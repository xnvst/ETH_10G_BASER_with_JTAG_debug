// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Jmo6Zb2IQFlDHbKi2c7GX3x0hpeytZL7BdErMgd1rV+6WGFdnrHCXW/1JSlpwy1ag/gxcg+q+zv0
GhAEZl2iIq9DbFvFe0WsY5fmFL+aZJlKDD8v2VZl+ADFUCtHE8qmD6Vz0qxjY79vLuk/SH6BCN2t
wyHw8KJF4vJ/JFt8x+Cxg7BkiFERTYNv4tymUc0dUYn1mJjSaaHyMrx1LlOlb5x6AZXBUJzC7JUC
Hu7JbtP3E46n6D1BBAXDyATkGZ07As7K4783hycC5blbzAuO1S81QfBBSqSf8fsjXmwTbBqNLMT6
2hn+14A1jN9qqt3YMZxlmpDgQgjuMMPlUqX14Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
bHq05aBpIXTGYVbuMXZ+8HuYpf7Z7HE/QI2zehSJlArRoJB0ajuaMA1PoFjLKPFzx0eXvTLzNbHj
jqZ5KIZXWe9wWy2toNyfpX2+gWnGfwe5MzivdlNuZkqdMET11kVY6g3zPmNg+32GmAWyMalgiIFj
Uy3Fqsvcs/fnZFb/2Eg/JCdC1+hSZgd9hgNwH1q5XM1ZA6L3ENz/mbH+iFYOXE+2dFrZnJdA/to1
GJ0TXYjN7Y/22dhS3Mn/+BLaWAJ5n6eNGArZCdB4Wy1AkkUJuQp4x6YSztyVRLpjBquvs3CVq1+D
9+L2o14rAosFwVbyMSvUNz54Ndo6r6/XGGmY31GnVdzeneNcMOoYXOoo5TrQ6CQLqSIZ/HrYONjn
aSpIc0OKGkyooikzR5FgQ6Uqwe25UZt4etUCg7Bo3kB6ZppBRruzVFJA+gj8+BzJ+SNns727nRS7
ixgKPYpDQTtaHll0w0NhetGFXOGmRPDgYp+AsxTQsQDGIgkwtKUxR1XOvWB0YsGxXxJH/zM7OcH+
IrlSZ5+fvpb0PKY+ZD2M+Rz9cBsRksw5nrNedF2QQfy5GC0Udx/GL1DzDe+BU/0OarQZUTJVzZBd
UT5bHj/sOyuWXK85c4LqtAE3oAoXDig6slHffU6Wi3+8Pi1MhoaSKtLyOgqYGCJn9uK+AS8Zp80w
OWvay09CjAxc3bj1sEdsHGpSJoCupRsZDW+bH/Ho9CrTqfTe2Gh0N3UQ3rohHVM7ypjUXUFyYYu9
/3t3swBkgtJqU19dBZFMRwQJ2+AGLRm1EgRKYXtLRg/AwB5SpQI3Onbxn17FcwSOOiE7+CzwSolL
UO8I9ORGuXTIExlRMOPo2JthPxHlDDDSmWT64WvInwCOaoZtrHIptWUI8JCUKuES3Q0uXDzsQkUo
efdF5G3kU5HwBOjFw61A7TyJiqZmpqaeQ3OO/jV3D1rDBzxTdA6z6pc7iObXZK1PiEPUYkvysJ6T
BqCpVenFAFEXFikQBwOMSt4Y9iZeDC54kHC2iGJjA6XHieXgvNeEQhJPXMR7BLa/tge83J7nm7Sn
hGWShgZZbzOUr4G+zOE+UtnXQKvY2GxUDOYll5iw5nph6SL5NMJKo6guG+bYdRcqp5gpVPgG/XtE
XOHjtuP9xlJ0hmAxJbkM7eCmbbBZVo2CBVw7LQD9LglKAg665sZi8vSNa04g9xLVLNBF2sMfOiCD
w1WuDB3XV5KuGxciKX0vqTTzvw0Lz/qazzG4PzO0bhcY7drhNm4udNMrh1bbQ/lnU4gWBGkPwR+r
TY9lCf0aaDZ3TJsfJeep4bHLiauEY9YcY++jjenEHwZ2bXChDBSxMsrTFy3TeDr5NZxg84s6WAgg
rYulm/H6FwXzRWM3LvHXaWRvVOu2IgzfCfjdYaoC9E8xI0Ft9l/m7mwxtDX7yX3+9DO3sIbmfI/f
FPnm09GZN7OzVP5dFoarb49bErRvbyC5ntQVW7FQzXY8UMHnK1HKHgoC7eT3gWZ+V6/GoxNuxb8A
VWUL3KG35xC5KLYcLQ2LIif+PZ5Ll20A7+Plte952oU9GZ1Cm7HF6FSfu5D2q+P/iaW76BROy/u9
wzbcZFjeOFbH1qFbPaVwv7DwoNKf5bQf+d0jQs3HQymoJqG/iS1fSQNJQJjgXjMiKOHSVPkQnk5M
Bx1Zf38gTSaIVnjd61gOERT048bgAcR/zT39OX/0dm5irAuaHGnsF0rHp28e027MFdScxR1xFyDd
DQFv2IfT2JjaJufmtWjCH+aItW7EBhpOTVx2Nzq1rnY2mVaiwbiW7zwFfMXY0SB7w7MDcYzDeOHB
UNeDjU+izAP+kCGgoEEWGWoi5JNMoLpP2mt63m6+RdIlZsNnbE2cNT2qdwS7V7fYCBpA+bWCV6xy
QFFvOk4gaagbIijyVB02yUhLe+quZkgzdPiwPW0XXTO19T/N9rnTwWsjAwD5xJGkJonF9g9Qw6fp
GqmItrkVRl3ktu0+uqa4q1rN3EBV0xZngb3XgZ4rTlNF59HvyBcNjU66FYrH3ritRkLU5uE+gUSC
4Qv++0lQF/4GwAgRVXlzsq2JjT5GUaF3yHHyJFgIh6VNtN1jXYNtvgkyFab2YvGbU1XcN9aIRj3U
+pzz2DqzLWZ1H3ZsX/Dux7EUqwODn2Qd8ZIDdZZe/eRdpk897GAkU2esZi/egF4jurnKMBvr0adm
MQhj/OorClXnRgxfNPik/UKEfyRC56NIDpM3xD1hNiHur5bfkVnxX64r6uGLadTtzGhUp02I1Vzo
oturaMX9hf6mqn17681BW1zSdFoHEnPUFZ+55iACO+oSqpgb0/IWrcJorGjd4c7VnTmOZJ6GvdLD
mnLLyZE3ufNKIAugKbPssVxIa5GELRunBdTbaRea3FfTubzDxe/VwkOwYEMwUewPYDuQjXcyZSSu
Zw3TauDNIbArRYVE8I5aCVMkVHabwT2HwZ9IKNM+NjGhIREgOmbEZ2ASHAVy6NsVXDwNUF+IPd5k
oJI5hBT0wcwlXv1Oasymc1GKxQmbMo1/mWX7WgMsB/n+laKDGW+mdX5E3pnfIdBLGIOg90xrtrQd
Gb27zkkejY47Ke1nyYUyI/R70rvgy2aCEmVgp+Xd3tQ686DP5LoUzQTurBZ3jSex3UXZ+2tZNr2X
8KLZjEyTm9kyy/MthOKoTLjS4zBhWpHtq58E+H5GSMzBfJE/WdAHOcIOeC1e5iAW21ng4DTcKUdQ
pn2ecsImkdsZB/PY2yLyMicgXROhptf3AViNGx5xoY6epUUzrfag4QErFmsVmlkVoY7RfPQ11UvU
soVPhswM1iY22OHiqqE1DYPuF2nKMSPJXsVnQySh9wMUsdJcGEXMXgy0zhucmQrBdhoXJAdBD7q6
z+zna2H3gmxbO7jiAYk65O3E0ksL4toexjK/NAUPikvE/iBG2OXG8Y3XjKJZu9vqZit4jfbmrDSW
dy9C3vMWrVH/sDPbGgsdkcpn19U6RwKydBWVeWMTKe3BjqSz7b7AaoTqHQ4RZyNYlDWgHoM8Mbrk
ODkSofdhzW3CqNp1T+9LFNB1hOP+Bndbt1Shxv+XPMtUQvRwB2O/IfABK35T3mk/tK/WasSeutSy
FhjUBFa0fTncuBWLIb9xK0H1TJfGXasAWacTzmBmk4ChLgWU46I/MgASNKwlucF8Wnd7v058kMed
XoNlPD3eV+uDbvOpjvJVY+rv6eaBh0+Vg5msFuCp8XQwzJBXWIZ8EU9a5H65ioHYVIlmdWmPmaF7
Ou89Q3CPYN0WHBQo35kHDhBNNtiJh8gD2STUyJHsngavmiWBD2Kv5GYo9c9tGHs2jeX5wjn53bUc
8UF5Gutk+2xIycowp30RFfp8GTBc17/zfhKpKJAqgb5ZJ1kQQ6zseplNDg5MWMtctajmNsRRe4aJ
2M3khAlvBMwVc09VvoKzxv1sdXch7Rpntaws2PHuy/xuwYVvUbjg138gobsB4Ayh4eKsyvD2L3Kb
IQk/NtvpT5juYBQMusdhsZJoxM3WTRLNbWKCw0SaSlbybsm5R0MfdTmNxvkktLGFMj6j7+3Ir3gm
9S61sNq5vJ+yncKVC5CewVEqMVpa3ph89wHP5+sTwXB+7/K/yIVxMexN5tK9WRcW/GPcbaZ26rvh
xuzIXfhvum3AM8/zQ2bvr3KfMWNixpzJXAPqQCCaISfIXxedZTX6qhZmQZKTGIKaem2yVY4n2vUq
8oabHeTRLBtfUmxzzqnomlOkyvjNafgR8l4xo2s0s/yRlPfchUlZBUznCaoBP2uJ5kojQif9+XGr
AoxNSpauRF1rWE9JLGZJyf7YaibE5NAenTVflgQAiH5A7AD/SUsHmG3NJROPc0Lq0J3sGcfiMbsK
xf6xT20hrIzM3emvf9oGq9EmRcAPKxR/xff5Qj4Ea5DEPZjO6JTGZNa9Ghw5gFf49nUazyeYQzfk
QxFCSFRNnXa1SaIgT2LvSREmg+3CpT9fYe4QRPSGndbZ0eATvc+CUVNWvqSAFLx0CG7XhLYdi5z0
M9GrkPp9+FwxyM0PpJjNIbS0ZdCo8hj0NOwwCYI6WWN2STkum2i0vXqOQH/R7UzFiiyGu38CMLxH
yUxo0MzuGNHLrKwt8ssfVQqzSsffGOWtwXHAuycFrd+uN4XUPmCRl6aH6+ItbkaTeYIXKKPbeQ0r
s+jVtpMfMEFwtx7vK0TNjC+iiRdHo/zEt0pEKE5ELTrer4KT9cMfH1ji70Zj9uCisEoLrlFMll7v
gF+KSl1XG75zb1sjeWtQyjrm8fw80COjKvtq/ZlsHmU0PDez9wnCQPCNBP7pi/oX0qirKqhLVfwg
1RjsGt5lg0RbYHvdMCZ2NNvuA7g6lPeLgqplOJIV84hR4+o/dg4ML69AqgQEwxBG5gy5KxEBz9bh
L+rHlJ1sgM/ju0IpKgk1v0Ab8hErMpeYnp6QlXkiQ/qujEN8fDCfZT2B3Rp9czcNANXTI7ynDLOD
PRd4BnlRbdyCQ6NIToKcmReYorgPKHZOEMp7cCn3wsUIIAi+AdgRiWAnsm+T/0WeyrW3jjEB3XvA
jxWh4f4WiUr/dKgy64NdeDEfuS72NGNQdSLK3Lg+hECtN1iAAStDjZGBNr/GKD5xQdNBOSXfUuER
tzjNk1dSokBEmD8rjwJJY5EAjd8sNsbJftz9HDr7GY50jn8ji0OUCTkRgGP6PRGzREI2hYDuqU7x
fbYUWvya4xiR9/ydw5B6NvhbUUm11FGfmjI+Qvmk6yppsf+95YDH7BlW8lmBLh5Cj71G2N5/7ypX
TSA5oGOaG6xHkiH8q6J2P8rFxbkd56k5IPjlOtJVxo93++RJTnt6c9cve+0bNBBAkSfCotijS/bb
7tYrf28viTvjp+orqK7U36VCwMXteVPml38DqEbpRBtbJuNlvZTSdWFTNYGW4EnI5MAShsqWrZOq
J5vqp1MCGBHhhNCuWUx67waSwbx2qrVaaL4hnRxqgc8hsRveM5425cJnyZUrFFdxG+VYRx8SbSOm
VbybRKId/Eb1N+A3AvZhal+Fssy6bkRKv9GS4ecY7BZbY/ZCUuBaFypIZiZg9NgnhidOzcq6cOz+
Bj+CoMSNYQEkC0ilhXLSMYkAF3+0SIIL8SpEo3QnwznIPNmCuIp3wj3oW7XnR3xe3w88mgILWkaP
Pi0QLnE5ni4Gyz0YJfxRaw5vNTZVejlEyRBdhYu/ssy90Ao+2aNSRs2nZ7lTAbPchBNsfgmBK2RF
yktnotQeC4PZAqkc24BKUg92Eh/tDvVFWkAiushrbQHPaRkWqV+8SQUPl2YyZ1DAv3C/+tOg9Mxg
EZlA9h/Ppyzx3yRyAtfdsPMMGymeoVZw7+Iaak1UgINLJjGyZacWQ/12VsOwWdA/n47ngnTRjvko
1aaYW4Lr9nEco8FWRI3Gd1Njh0rSiGioeRNmcn2VQFB/4q4NaBLQUQg+6/CujmCeLiPVrL6hCFI9
Zp3XCUyLnrie7Kzjrkpb0w8+Ux38yNUWzDhqwFAVtaBqpL4gm1BF3fO6aiB1BeYSAKi6QvwE4Xm9
cPhRe2V1KmIMpBspOyQRB1YanMymA6mLY+ancqPBwTvd2vKZK6fzoU+sMFm29NJsop8FENsenn3f
U4s2qv/2yZpeyzNlWbowC+OaSpfMLKhDJHrqSLoZvF+O5R4XKCaKr9jyCfI6z1uJMCPSXAWeOTTK
UXe3zjPtCs+vVZ8IgpFNNxQrHssOgktjGt/O/pNMMf556e9HzLMU08IIPudXc8UDsGd46smdZB2N
9yPXEIkErHxTZblXOYGizB40vwDb80BFxbT0zYSV1hUlALSJr1wbMpKb2SjH1nQk3+gp8vIwxTlF
Rc0OSdXDDndlY1uqDzLG4zNIDMX5eee9XlG77ngZ90tzh/AQzOBeaZnGHdHdwyXIMN5HpuNYJFFP
xB/C00Rf7XoOPjBrxh07+izzy3jA6i9ppRJk9t05lUzpY26pbDYOAsStcOrnP9ZC101t4jfDK1E8
4cUTre8P5WiMSXX93PSruNqqlOP2cVUgO+2CM4r8Mg3GgrclAOiz+ZXqa7vo1E+7YIBA5wg4WEXv
F1H/xZlBblTkbAZEqBbWcx1sWKVdoHyXqEOXZJCvwjIXCpK/cPKvIdhlLQXBe3B7aiE9mVjWHozM
RKmZmyLmHhaU4k0NnpHopzYaHT0Eedxij4cNel8LeULwDSkCGzR/gt513p5079Fp7u+O7QJnsy+a
ruStxNQj2nylIr8SFwL7PKfEM3bPaoaq2RLoA1pErfFmMnfd8ZYlnOqZB2havQd8lswmI31zuCfT
D85HrbluAWuj9tXsz+XzeH57HUnzvp102NbUyEWkTNQadffw4XpnHPDg6MmC914yX1qrE7G9EGOz
/9xeZIdUYYbq7afFMG+Gr3b+JwA8fKRwwxVMzUjxc5x90aXWTORbNjycKFLQ2Yo/6hQlB4uhbJ1X
GHC5Amq2cSA0Ef9tzTEa2ku9Qclxg8qy5cofU52dRDaYJ9ITR6di/ETyGfD2pOa341AQEH1yXL4j
ZT/YUceNEFHa+BQ7Svnb5+FdrAFAJJGiljjFl7EDBjvRaDvRm230w8kczuqCuBwHHs3TQa766x68
PVRn48kupPo70V54/IfQJXKxSV5o6fpeUfnAeWi2NitEHte6VjIlC2F326g3KnSC9aMhBuyPrh9y
dYokuY8D23M1a3N+L8St90XF7dN9HZmRNlFcNATyir5pdHH2u7aJrCiCDGd+8/Gg7vP3I1nwI8Sh
ozFjuV4UIwEAG/CR6IRuZuMm+LpqHVLrzgbyYMCca4LzauL4r6mlf0P/XivVv4CngxrW9v1gqkb5
fy9kEqzR667XIwI6l76mcFNIv8Dl5Occ3ij084Z0x/6XAR469zS/hZfTySgJvhmZoCrOmFSWRt/r
P5iaXqncTUPwZt0S8gsATGldAUawcyfujE5QSBPiGI8MycHbOdmBPtCzTaEl9Jx3rg8uV8NIvL32
JDcphn39HfjtVZZea0K5ArwQARStOWkZPEfK4T+dGuQ5W3RWH26fAgl6jO910OihJq0G+CDqucW0
G/BuCyKktKUD0v5NMi1SlvtzDzEEB4QoZevDMvH/gADpwx9+JvpiCEdEuY4Le6BPk+A2G3sKSXUR
UoCEwjUKEqYzUnFBUf025JMe2Evya/MP6hVzlnDkKMZntB8ao5DTFTReRyacF6dkTqxqSAgx1TKS
hRucxSvUUktY4Uf4w+O45w8ueM74AW8f30ogF/Jr629o4U+ranwsgMDTtzGaSNfTbgaU1sKwnUTE
Q8BQaza+2dXoY2fCKs8DvWqd7gLVp1Ws9zxqXWCez5uZ6xiAaIyIVrgQolguggQOMWrbHHakOmji
PB1V/xstGIWwphdtItqCPOuQpu7uFnyISCMAcKM9AcuTuA3IhA8SwiSdZiUqhKzPaVvl4Y5LEfnk
lC409DXoNIuWuTpCTpeJkFKex7fXHBBKMEmGD80ljYdriIBkcPqZjHgS7yb44Ixo1ZuXA5xpeh6o
raF1QPIPDSD4xkBbYOaeIpEiqOum+QJqyOj8X3c6z2kJ5Jt94usglOis+seRRUKUyafiLHRmNUIO
whv9jc79W9SlEZCGDX/Ae3Nb/8M0WFIb1lraV55D32g5T7o3YeDZ9kgO8rJGJpNVA5khipDm3OQW
+datHDeFlCV+2TDEjSGV/GzAAyBFL5pd5jw387Yh65gUnA9L/M2D6MiYn4egMF33RsdepibjUIMx
qPAPypgK5TEA1I/db7/c24UjNNenIjS2FfufwiRRt/O06acbj7DJfjabHTEJny78zotZie/QT+va
ta21G2hU8KxcaqkWn6n3XNjfNwFuBqShMT7v/0bUTnvJ8KHV/HtOTgUYOIbITmwNky341BUI7YYU
lOmSB91+0l04Wm/0u2pZ2+LAvvx0T330OylSI2F35bwJD/6U+ziUo2mYxYEorVMtuX8H1VJVE0He
qa/UhJOR5Kgrcdio8p+8hEyaMazqFTFg70l62SKvsN/4Ikc5H15LcdjKvNT3A1/0LLy7EkBIUQWf
x76ak6yACsO/QgORJNRubbhfBTmxT1eL2Pg7jvgkbvo9pkaAAOxZ/f+ZEto/Sal9kqkjpuc+6D/M
MIG4RX4x7M8lCyapsOPSHDCGXRjrIKSL0aklGey4LN/7pkBu/5VPEv5E18CcKLbnLAAg06Q0hVWH
LHjv6UX150NRM0GJPldqaZ3E5U9O3hguhplmugJf+z4v6I3567TlIVF/eWFaBlV8zkYfu18aUGHE
zCNJWvXVMXZ5eU9oswTNo1e54PzOqcdevKfbpjpn8tYDxBxczo6VDsXBa5M4bvKr/zKefettSL8c
I3PjqL1y+/kpqIuLxG74UyYBhXSildV2/1X1Ntg3+OHJq4tWD2KRndysZqZtit5nzN2Je3cUGz0M
nh2tKKxS21fQX6hLglE34Ghms7IBJlD/TnEYqC0Pq6k6ytKbA6VfYLivJgAMj6v6UyUvODS7i0dx
IcsTeEdyPrlc386xjX/6K3UYx7R8yo2yWrjklC7M8o9/lcW0XOhqgJ1Z5cBlSBHgVNZay9eFgG2a
MueRYbb4vvmftfEdE4F0dNgHgiizGw3um3dTmjGd7ILQjWcFKjpLvpkc2BtSib8UZhTsqN0mmP+8
TZoEzgdh7SNxiW0gxII2JpUFsvwYCoZ56ALkcACoW9wybDvdIvIX0D6hL3T1qDjftGpNKacKPM6Q
mdPY177aoxjCQ6k2OWYAZU7sU8vsd8gBQCeb4HA3eMOXFgA58TtXsEWU6YVTawaN0lqi4a/RE1Px
EX0etxfp90TtG9d2cOxjrS+V23XUHjdOFUwFpFJpdt4p/njypsXqp8U6V1I/IQ5RcJmrLUHs+17o
0ajjSBlA4ppsvzfB9RfUfWSPwl/KkcRBMYu8HIOzheDvXAxkiR6/wJb2VPUznCzjaqgfzd7TMzUx
jLAyPCUMpXHd5AkWaeWHugVUabqSgss0c2pgC9Tf/pSNkDCizy9WjKgvURPWmEl402U3YWDSTjFV
RQFYJXtY66nUdbuWtje9mC1p7Ku7TZs4axBi5dHzL4W4YZgdg583xWNA7IlLeJskiO0ZCtM9rioY
G2m+ybE7tnG1qmtZhhr2TRV4S2mUgWvm5CYF7pkH8rgJKYKSeR6+0Hlgw5rIjf8P26MOtsnPKw6s
D9jDh8EggTfjALPEMtZrBy0QgM4C0PH4OyTZcaYZUrIYiQAxxUjAsE+R0FrO3i0k/lR90413bgUP
xExipArlBjHGN2DCfjSWns9WuqlDCTBvTHIuoXyd4M2Dv85B9VgpSGwDdffZMgQery+3GnNnlt1t
tWUvLg0luuzxDgqcTTOA7f5Bqlso1OaFhd0KilQo5NJax/UkkjORx0vnRrEB//lmxUIIve0U5TlZ
AFz891oXmiuuRb7taf1/8WDq1wZWDYRAmjmK+9ZD50AG4MaQLIqPMQp6wE16ABdEz6GF4O91LuGv
yBwI5lKjrHZ0r+QJzdSJ4pvBxWYRqw6uEVI22iQQCMIz5yHcPZGRETk4ye0+B3Q3dVTHJEBNcwf+
KGC0yJEnjY9+Lbf6siGAxNq7HKWc0Nf0jlGpge+FuKp2qaYmWK2IJm+MpkfiLp1z4ds+qLU35T6W
+Lb0af5cBD/5JpLasKtzkKMtBzKahv/ptwSEZUWEZTVCJc+jZ+wRuCNSa8H966faM+QbwVMQFtfi
4mqvcMYaFQL1wtaARSjYhQ0UxnhgTPkSNoe1Dr6Lwyh5CDAKkG1Le1tem+WP8cYztGki5EVHVzG1
IBg5eRz6WZa9lptWsCFGrMzbt+YQSztFGbHNLlWEyds9XVv3EeGHxnHlOS7pQJaeTjU8VvW1cI90
oR2VIALPRRe2gWHb1t/rzUp/HGBXeBj2sXFGqOVsXpKsJbO+Wuy8tfj0/xlT88TukbnWqFajXygz
7XKObR3Fyh9kTiKE/W7w4dfvk6f4wFFFsuIAQBwFUXivCZVzTrVr45ZTVWIPVLnYI3+iCZkfxNlC
rIlEoZ7U3IpeLIWdS4wePl3NlUZrUgr3hemm8whhevuRXNTQEcyq4vr8FUxz0r5KoEKy0jNsTpPE
IXjwckSr+0kjgGC743tg72Ob8yaTA/XeDAFsPrKogArI7d0SKKtwesWvAO1/UkkUKkAAg+2f1Qt5
KP8+XT53SMqZqfJBsC7UMD3PNIHMDo0MtDVCQ20ijFIJNEyacJXmwcztELA4U/k7LZlzaA/cwceV
PSyFbbUzl860P6qyP3ykloFQpZVtfFZQEjbLGI13hEACWwz4wZMbfvV8KsGPJENty3FSv8zi+T6+
aFH7dkkIXnMVoUezpSBsptTCuXhdP1OY6Bqybg/+E92IRiSjqK0ZlVCh3BZJE+ibjsLXvsy9I4GD
20rzqQU/xxHT0XFTIjWCKdWQytYwi2xpvZMR24bqwLKY2qx5BUPsbIFPTT7jSKd6WI9voBy2eet0
lmM4TZqFrw1Fcg5J61kIKwgxGTZyE96V3f3w/U0t2m4ZUgSgPuiC5AdNPgvWwmLoO1SM09TO8Ih7
eJSRkz1VPVG9uhTa8g==
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:31 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZTbyz1beH0GM3MSFe/XE7fHWYIMcx0FfxfzO3LnEhN36QgbvCIOcD54iYyDKRe80
M5/s/XPS1UVlHtWNVxelEJ/Zdcv3N/L4xT8K6d6lH/vXBohSssFeqaJEsc/Bs6p4
+k9lKHsc+siMz7HJoJCualyMVIb5b0wZQzGnMWKUTPs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11776)
IX+XRSDJc4eDZ+WKqaScq9QYDo0v+F7080Hz8Bb9WgiF0/DivHFycA/I5Jf5iBHS
dNt4P1eGshOTsTymmshboTspdwaeJ+0wORa9OuEzqLYVH+QOrEDq3jh3xRkeJ0nl
ucJWUQC1DKEO3bCIrP47k3/4WnkTeg73jiGkkhVHkC6UxHnBYOX2Y4ep5hA3s5Fr
iaWvDvW2l1DOwvVlmaPStmQwjw6nM4LuHM+ODXpqazSZQjzY3L9GBTOIHtaLz6zr
1JlT8a4pP9VN8kFPtpF+/riM3TjCurYzG1WVaffYJSMGshSTh0hZ7mGBzNXMhghI
pzbGKxHYaFO88y+FXl79cINGctG8RltXdgczNVRnFiVfYuvjulk0nKlpfJNZsiAZ
Lj098s9CIBYpBytmvYBrpiRCqKdby4hYWC6wph7CYNKBlvBnCZlgAXC8KXzIbC5X
tXSniXYwCga2gOqcxAdGIWtsdQ5cqJ7u7YFrq2p2fdP2Y7hIEfwYLOSAQl1LWD4H
FQwJJqq2h/ybgMCrWky420OaG/2Ppmzaj+aRwmbw/LmCDYahD8ehECm6kqB4Di1O
XTwb99EU0+NWLxzRIzgXjSQiLG+Rx/nsJbIPfvUtUQiigaubwDntmYZpo9jKFbmF
VR/hZoJSkoDtbjpwg196TkSp4IGAeV200HZIoPQ5HlK/RZlCveQZNPWxmSg07teG
/rVpWFMbAgX4e6JnoqG7I22z9I/53bQfiJZmz7adNyXjDGqWm8eJfCQBA4as/XjT
Jd2fMmcUiZhCTGZ5THxW8vXK1Nvji7iq8Kb3dtDQnAap26wkbcyewrf7dvaHCALn
R/BQqJqFDQMLfs/Yo7RIhcSE6dz7+5E5l3yg+kPpDQ1TMDn8xC8ytgTBFvk10Owl
gPO/cx+Q4pvBsO3+oUB+8lCjt1BZB50v7uFQHe3roU4iFUvuJG7HBdndZSzzPfOt
cW6TUh6+8YHto4WiA7J0sXYgPPbbzUmBHR0Y87l5L1F/c/0dY/DryvNswcByVkDX
psYDjXHL61GfHCeVf8QvLaBzuJnuT3N1s46+lPT2iWzecALqPl8NGxEQNPdVGK9+
PHxC4gO7ImNz0PxDZLRlKrm8EgmqqqbSS61gZWpA2RY+zB10U5w3EjEEk9X9Szjm
Rsy3V9TqA8ZSOquBpb9IYNGjTzL3mRYhv+uYWEs/+OiRP/Ywwbdg1V+fUwuth82l
VNtdhkxLlumsOwlHTfPSOjM4aCNAOwZ0Vr9co3KEpqR6skIAeaJndL5IElmYUc/A
M8WxkxTRicKEqecQ0RczP4wVC/UmzPuOA8vJcAy8VSM/fz6CoXDTsvNAELxUT9wo
omj4Jditrs0QUNCTvpQNbMcCZXuEjSU5bEIh7cXQw++I2BTF+bP8Sf9KLP9He4CK
gx7WDJx94Q/Cxu9W28UIvs8ommwp2o085EaOkHMLU274BT0/OntQTdJayYAX+kxc
eTSZM+32/06on3o6DwrBcq9XZ8RC8j7Wqc++4W1lKtQSuqJ7rEOqGx2Bkud7TiyQ
FZgRzx+44xihTTkS2fAAuYZ2K0fNyNastS30OTdKS6OnBBxI0a4p65uJy/BLwl+U
GfECNPJ6iRAgKncn/AX5mBzxfV4Tj1BF+MRW71Ixdgbpxtq3x625JkFH+n4ionTn
6wduVBbSpBczbbWf375k5aS8BDBUF/pw54cUOpCLlMIeb5HFmTamhS6A9ZmyJ9Pj
z0RGeCROiC3gAz71DIP8RekkU0d8MmNaMAV+Uncm33HLoi3lHL1rp8OINkHzio4+
YQWsF7P33s2IDLb/mv6ghodu4745wDXktKPaCFs2bXvJx7ZGViGQUFVJGC0K6P73
ekgMgXb6F/XBFiZzh/0vGHMDSGBQU868H+lvUDUo4O61u+JNIjqxspE4FQZSUv4I
wv4YR7HkEsyWsfueT7SU+x0rSIc4PK7IyY1mGIYhoizeBhcp1mE7J8sKCefbur7S
5m2DmNn5CdNN7BWRRMLzzdic56jb2fNdjkWtI0EHC64NQ4pLiEtvLT7KhzJAwLk9
i3GM9cMRY7EngnuQ5IzLPjC83BTu/JWdxlhjG8ACG8viaKejm0E1fcO5ZKrbexLF
BjgsjHTnM1r6+iIrw+fRyvxkZU/BTVGY/sswomUjVTe6Dq/UT3TDmnSdQ0gwjgd9
yWltMtB0KC3pzewps4iL2Wbm+/ZtB2mtrQvb5GWKsvecBEhT2plNSrTdAWOiXLQW
b3P7lKkVRLarlrFMs7lrrO+ztJkgBYh9a9CITygEvn5CkQ567hVVI8nz41pW5p91
R2UHJC6yz7oOfgIc6fzwDarwEAIRcdHBcAZ8zuE7mIpEsD9qSlveN5u5IkU+F8Eg
DKaDq0mh6WM80Vi2zDL3phoz/QPCNg+xvDwWYS9NToVoThGAAip0+AS2E23BcGIe
4lEDWA7kANCx+4tNeoBo6Qrph0ksrKfl0OTCGXcP70EvokjDgu3rBIVPArOioA34
C3sPmb5rOzeuEWY8YuT/gkm6SwjuUYJwcO88izk58bTWQR5sP4cKfjvxV0swmD+9
lmPxnzTUqQOGbL+L7DuDNijdkKZDtDjRsYLMyJ/kXK2QhjSXqdajaRkEonGkdLGv
r99cuShblzgl4+FxWr9ayIKGG0yMerQJCHdeMJlP8iolnTHbKdgVwGBM/PxzmwSN
R594PkIPVv/HzoZwUjy3kBlw2rSsCy6+linzncl1mGzLAHTAoWRHcpSLwVzSiuAv
9oJP/kaOONFp8H+o0UvvtWwe0+dNXpGohNlgctNftkyhjVCKKr16lZO5d7ytz9uk
FuRz1CduZdma6ARmhiQuAqIW3YMPLLVq1/ly4f2gBXjr2pRxWjtdigNmlmSrRsvM
kCvTeJ4vK1MyB16XcUs5raYDLh7es6S05kgL0pdNfbH3fUnMbvzEZ+hByTlG+8vO
vfEu2+ZrqnaeEbiQOy/V3mQc6pxAQj49/cAs7ypXGLYsWyOA1pCXSGCaq7i7/Byw
UjanHGs0ICJDIa1Z5y0f+Dw6UTBC04T0gyS+1LqI/dcZF8YP23JCqgkEYkUozfre
XJq/zGqDJ4+6UjG3GzzidNQH50sBXa/7wOdyD2bcNkB9z67WNtz5dW37l/4qSLD3
n9AFVl7eRo/gHW7AQ//idVFBrV+wd/0DUF8quZRLDEnsqxRSTqUNgPowY1sErrXy
C/+Znx94WLyM/pi4ZIgHiQ4P+jnNN+WDCxZH5+13o0Hf44nw4UhFnXHEjcbhHtYs
THM/QdmqHdZM3ksJ6QRYlIHMwMkxsstI+geptDf++KUpB6fixgd5QN53jiiqbbE3
45RNSPT6fbKI2EE4i1yL+S9yIcOo0kSbqyTvwz5Ae4qGbyVAjoRitzIC0yuNkjki
kevenQrIvsin96h/qOGmC1t+UWCyPnybkT4ElX0x0Uj+N9bfpPEn1dHJ3ed1Fybm
mIWiIKEiwqCsiQ/LbtAxnpGmPIvF6oCgqcpts6LHU0N4CVtoOE5/mZoNjzrVKwzP
X1xnRs0ULki4TNlCer6rY+UG6PfvLPljHrfebWG0TDubblOAlW46sPhltuyQYdIo
/YaZzEv3ei1k6aYftmikKo1vcChVPLhIPMqsEnrpxc4/FlAjJFv6M0BE0pXsRF9Y
y6DOSAKzdblxC7g3EpbZGSg7pR3n7LDM6fCtadIRZFSbqd3R/bTGpfJfY0zg31nV
UY87GNW2Hz0DWepxa2jD4rrp8ownMWvQ1PJW6630oBO7O08SicHUU3vf1WYGuZFJ
O5yQ2uwSsC+NaGDotYWxSZgXlXuDzW0yPfczR4OGHdy52xn96k4pSHqYr19otKmP
1CcYdGgn0NhBPXlZBsrIESYxBIGpWSHHmqxUQ0OL/oOOgaEhaznGtMbfnwtW6TP5
OblY6l9BJSFkiFQEj6OcZb7nh6sAaj8356cw64fI1eW3iSjCpvim2Pc5upM2yW4T
tjLo5nh/lSDLUyNxw3PtS20AqMuw1fEvaw78eq70d6KN2/h7m1IicvgMKes3azb5
/UliYIcdAar1tlocTLEGwJlEo/ANnVcvEiV6t9DhCYUKygsEKmvNe+ynW/jQFNMT
i+vyXkvlzziNQMJH4Mepcsjo+c7zF6WK8zh9EscahSBlf8MPnl7qqwXGN4Ix4cvU
czyv3RDko8C4HfEBiaOWd6Hjf08h/tSOmSRv1KJehFGHlx26fpTlUdDkLXmn/mQl
7U7AZXRprE6IEV+6+yNrw23FxDoqnk8QoyFOB/pMfBE+0rVjwU0kEeq1L6W+XEur
PxVrEUjNWTyd1WhTM0e+XNdXduklVDzAS8AeQ+2lF9GG8aSECr6lojxfBaXVd2f9
NeOCHxLY2VMlUh4UWsd6waddCMseQMKWHwHSUb5O/ke8wkbgfWOckZ+WR9Ijvh5W
FlmtZnFB5SbG7GJyyxTJWIpa7GKl09/ZzhM49/X+aZ8pGCoJFZBUSQydSIy03QMX
2jm5MIokNh9AVS5i/m+C4VWg0rS7/7TWZQUswK58Ul48BHCpt46yhjatD9ZWdZ8A
KqeKUYbdyruDPHW7zp24yYbICrPgi6xSYWG+8GODt3Vw5I//Tqe5/vy2qBXB86N3
jPmH8uzi2qJ2dLNZx4AvF0gjR1vJE07qRgRViYX00A/Is3ehLahbNLJjqZLN5bUU
b4bCWcujlo1bg+jzlqGpVFCZ+BdTzIpwBdiqgJyTHbGNWqmEyW8bZfLmjBzRJ/Zy
upV+MmQasacffehx1zMcqjuA9ZqTWkxJO/4ZXeCGkhHjUi/i09k2zHFalrwApk/2
vwtNexOJ22QOKDEk5tnnfoqfYcZzXZPgqVNVvsskCr9kKvlT2TFtitCl/qFZ3Oiz
yjGE2nDNKnD/eanGo3Vz4Kobvj45EhLJ9NTst+A8jKcDIMnvAydqDi/MRNHfEXIh
uFHxxt7SvHaq969/lT22NheZmESKlTt4Qly0QIeeF042V898lY0C+HkJrwKJdR15
ftdBIF3ZOyURZs/phVS/eikdgoFw4j7Nd8hZf9p4iAUD7aE42sUxyPrlxhM/nFJI
h53bA/zcYkV6qcHRJr0eOfEtAo/RFnTMMymRZEMHrXgrtW7mWPgFi/EHV9GD+BZ1
NY+AnOAxjmYECg4PrXkN0tMGhsOppp6LQYrsYB53qKMkRJ6fQlzYfe73jJ+GdgTg
oDTTjAlcMMLrEpCK1QOhmWeRPtsit9bmjhcntkX+GHGAcMmOyDDWMBgiZNPNBRKh
gitSVB2BOFZPF28B9z6F78uy4w8iqjzGk3oD6XshwwZZSdDSdHQIMinElzSiqyIG
FQwAEMPLDfA9gu4m52bkWkNa67f4KSz7g5VC2/kRmqKHbY7YSSQYbt+nvnKe7zXc
KwcNFt94iugU2KyDWGu1V0HBuEbqQVmNF5KK8NtuuWDE9Mx6sJ5Vc0/c+fleyAt1
ZBjwffyH0+6V3pNaQmun12CS4bFdVuN+7QBnhfAotUnoQAGoWeMsqIILQHPy8O9Z
aYyerMHesq1sDwXkKYKf9SmWpml4Lwru83DyAZFsKsZSIM2IQucgXDN+pCjZeQXg
LuI0NpOUJ2RlAwl9fCyQ9/cnycyS+tlO5UJ/COJWZSNt473lcYCdTBHdmbKPSYYh
J+Qgs/0OAkghExAyv2JZJGXPvAs9jjS0GRjzLyXnGrNyK4OD18fewREstjkt5xrt
ZbUlhWC7RKsfHMdr0q18D3yy67bL4zX3lXs31+GrcR66yQK6VOMxAn5qOm0btny/
wf9TPCWG3YQUM+EPwJdPHOjhPTR7XjE9c0W4mIEXWO21BtEfr8k92zCmaMBpa9qM
E/koJin4TAV131INIiSbjTzCEu4AkWn5Vtuk/b2JBs3nN+Cem0OM9VIsemuEALUW
z7Pl2LTtLEuitXA1TFojh1MCYJp9U2zIi4piYHb6NR9Q0k/z3DLW3pv8ZKYlhbOw
uvwrs1FLp4agviZfMx3U3t+teOfftJfrVwkadFLDf+j1HdjA+XqZ+a9VCaE/5UZD
op/YTlYRCdCcP6xQUUfEPYhGUkcj/FIyBztAF8BLND+42n/KJ6ZZWqc2vlTpFMMA
70NkC904lQ9ATaFHJLObMo+R1e1iM/1yQovgtkHDdDpx/pFSYzdesIS6yxGyOZ4A
LSqxNspQDYVqAYxxj7siUjsykJqYE8qyxII8lPcpWM9w500GGWnDj1Oy/N9Ewzak
GgeBEaznWAUAc9+rp5bDFzPi+g3Mr7p3UI926kdeIL0Bz43GGhK3TtL+4KRuWS1g
x67kg6fseyFPzddXTTJ2z3eHZG+nSp0iG3DOO0a4f85H2Gqyh+rW4RMHf175/Yn3
RHvdecs57mv3o1mVAKldY4cuDyTH/OHTWx0Yjk8VXJ8DT3u2vdYSdicNFhozJZ0H
81q7di2fUeSgnE8nUFWlzyb2Izyoo2YqCTVRt1gTyw/8Cs5pUoDZe3zA80flbhcu
nq69BGnvigivkiP79DYmWjk1fd+ZEIallcX4qylRnPM8sBj6O0S/1RMlMpSAIvlK
MkPjxGU8voQmQP7G5IAgF0OIELb224zqNYH593jdssgh/iSCVJzIKxHEMQL+//nc
W9YATgmrSSvQrCJyIATPyoApEUVy1BAeR2CbxrHhQHVUyXfQ7GJVkAxArHc9jV5g
lxkl2eBpzSnJB81dCFlhm9JVltQP9Yqg/laXq05JeV6wHN1I8nBg1S9c8MO5/nEb
YjPefzltvDkVsAnitJxNnvSNcFAPO9+H75YvjhWnOcOulDzWLpswEdOvh1WXJ3aS
oUUvkLtid7WF+J+TW5h2DrRLHKg0sQ4SIER5udjexU74LPQkb0FG84xx6XMfNO1E
TwuoViTR0YhfHQ3W1GdazJ8qbfLX2cXUg+UdyH3qIwgZE+p2LJM2gVupvhrRddfG
mDAT2KmicpvImlhHBeumlBiU5g2k9Ni/8v4BCM9GldfcT6Z5NyDWMTdk/TrqSuVv
1H/d8XgUXstpFfMPisLClIcmNH+uD376Re1iI6+1JMiNXa1f4w7j/3r7dIegaAvT
1ywx5AJbCn1icA11/v342O7/LzpPQAcapKQQWCj/ltyd+dn96kArbBfpTwxXN3U2
OOqjFkdUFuc6heOykz520thrnT9WXAJKfDm0wHCEgYI2oRrFMTmDp9UqTa5j/8Bk
mOgrXpLPuREg3240R1oBrRo8SdHZs1chqsIvo+xRjCyNT2uajaYXfWfJdAVFP8o3
FtcTzwdlJRrjI7eD0cG+tYL8dszm74GzeS70XvqVYwmP+u7NcdQhq6zFzn6+keyk
cnR8ZromHyhzTHi0Ej1anHlmSGrWpgnN9t7zRcscV1f/lJSWzsrNcVYQxv/kmfem
d2KBzzCkQKPbNVDJx/R92Wxgs8F+xpIZAc9UE7aGHkvbcyfnRZny/vBK5Bcal5VR
Y8KnPnuMu0yw+lRrgi9W3+eTsvW99wvuoDwvInssss5wYVoriTDhS09qW+1L1yXq
BHPqiuhZlegaGocAbsyz/R/1/RG+lzwvaHBABW2Zig6fOLQb0UbNV+utGRwKdC+z
H52NgwP5zwg7filPy0RI/JhPiO2jP/9sCDhnSTFvfzD26zEDBYP06izJoOvkKG7H
39xCjQBxHVaMVu+2zZuJ2000CDX+3Z0XJ+7oPEKwXwZY5a+OmnivJe/ci3CKYRaL
nGXyVe7ykVNTOZHFYkkevAiDiEolXlL6MWHxVl301mHMg2aOPTkFzETfeT7Y2kgL
Vg9VQFjirknVdmSofgrFDYj389OfZRt5ytZojWz5X2jJQJpTJCYEVK70phWMlHVB
4LQ5/PA7Ltj0hsENa4xoB1Cf/fCp0xLUWw3Pv2cjHecTGnSOJQZuADm/PwrSSJYb
Z2SI+P8QjuRd6cRCNvqJ9mAgW+srhfnO2i5sGqR0cKSmiWUkQB1fS1iVBGeRQ1zO
BlUg5940qEfUJt8FWCXV5eKrFxjXciRdU9BlcASZBq2dVu4abl2UfD934rjY1nYq
XwEUSStfyuOgd4cx7HXpWE4qYWlv5PFEgXfJaNbo92h343cX6n0P6pwRsFL/uva7
4wFwZT2NFX/gpADbpRq5SMroZLTWfH/uqLqBlytBdj/pg/y6AZKtFx26sej0O2lo
lrZx0Kv9PNc3yw1+c06mzONDUFCIZJp1CTHUACz3cnLLxZN8vyw6ScUtXSEDmYjP
PPf28Nmp8lxH6AZ5XMYMFmUweZ0qEucagp81aS17LmKKrFSk5yk+0vXCBRmEJOKC
dZIaeooKkKNmln6dtXHE5Wcb4ziQiKrYMFuZG56j3CUiMSqdahxnOKjNMSoRe2va
8MsPXbHSDl5LT2XwnWzVGPBJTFi1FRYd2iPPXr9/E/p3lRSKhEkQjUGYCff+Xrmm
TbzdlEYGmtzErfdJrldwRuyPM3hAudw5V7+bT/ZV7gA0MvKcxhvVDKTlp6nIh571
xU78SeeB/z1Y/Sa1vKpT3zoFwHTvcMCqNWW9SgYkhsDXG1i6Q4892Dxm3qH1RR6q
Ehp+WYXAWLEtBg3nqzHjCwrbvQOgNViK9AFEkOk1BDi/gWh22TpyKpgDBwbca4FZ
E7Cux9Tjsp6gAREoRKk/q737YwOgxVrKbe8MAQhf4qreAEjteGhi+E3q4/AZH1ZW
NeQ0btK7SY018P64hC4Fovzw4tuj3vh/+iWqdRT+0JkBO1rr11d40tKaYV/iyLB+
XLWe/uP8kN0vJXtHnEMX4nIDFGsHMvBuBOcdKuyDnk+yrf1enObzaDGKPS9/LiJT
uFTEgK0KPOLJRFPbCzH1FvxLfIUoSuQ70VA9tYGv2wE7UlZjtjrc+m73erqtvkUA
UIkC4yAX3o7g0b3SuYWW+TIg65d+FKx/Bbgj4dETkCdlSOShYMD3++UXdSr/6dHS
wixP9kwTB/SytEnqnZ+BluLNdqOH4Kz1tfavpo2R6q9VpOSiUYovOsRFFK2bKytt
ezHXlzx3ObgYrYovvLX5lw5GkDoJfLwOt21Xj2Z+vpCeIpFT4PlNYUMYUBmG6zsd
1Cd+UINTyQJEdDdVtlEM0VfksQD/P3kPbl0+OW3P13spQJtqQnFYzTt/xICCDQcK
/TXXisI+mAcE+L9wiHSz51pQSudFI4DAgoiyp8BHlTickVNiNrCzdbA/cgvP8fPw
rcRtXVjjbiYfK8J8ajRMU28yaqCUd/S1S2bcGi6MerUXsldZJ+a2KDPD1S1xnSqQ
G8me5JtFlSh4t5pyFpgkSWycv4Tq8cjS8yZt8DwKWFvTPuwJPLwbF7Tiz20eLh+8
pGFNnBtcF7IlJP36UmSxDdqqc4ImX3vH/jUK4Q2U4E064A6JAslVMPqLLraC6Sqr
p7FLlmJxH2MnCmbkfjXHGuJlpfsnOM6Vec6zZJIC1oxmfo8V+rJHYHGdo2G3gXpm
yHHmVt3pk18+xcDtNzFoF7BuNte/fA1v/afJh9BS8gODxQVfYhWjhTlRwClUGYQW
hhVjnjcx7HThrb0ni7Rupp0g9+vR0Ed/AY2bcy1+YWprW0b0DzhCi9sjR3ZSZdLQ
KRKVFXjr1alFerXjomSBDSt3cE2agTSpyawFMHi0Avfg/LlMO87okVfFMfbOOLtU
s28rqYi2/TvVh2RRfx9BqaLdVCneYSFXQ31kDICKgzZWJfRRTbEDOyg9okGjb+7l
lVO809Yg36sYhiJylYOFQJUmtc56YSeLE0kDRycQpGYtKQvmsXeNtd7FprZWtPLN
mqU/nDbLHF+OI8Yb2D5pJB9Is0QNtAmDb0iIKDL9lPIDfJKczTnf+TcXHWGOhnQ+
cKXBETehNHVJ++DZqYlcsmFr5hEerXo0YU0zTJ4wNwApgrhFZ80PxjPgamYhV4kr
5mM/Ink343I5l2bVeofmWdZzDoRWX4InE2ZQsFSZmlcCmUs3jvlHCOrYqHT/+3pv
W/MxQ8/OpdFurVzwqetffgErw3QAiaPLYIJGshS4iORkk9bklInYZ5DYPbqauUU5
iB4/l78be8dYe349OLYzarADpfbXUeK4+FQxwK9fUBWaN/vUSsW2TkAQ5cjq3yh+
gxeXsz1/lahVvzY7h8aqHEJzgpMsvWgp/B10Z/L28hhYC7WJ3pb0DLdEYsyrbKsD
kSqyTwu/rrcVCP2YnbbcpXVqIcl2Bf/PTB4eFNOQwvxk/Af7VVAT8Y3VOhVTyKIa
nV5+6XE7Jpne5r7u+K4spnmFi9fuKkEtXoDyxa3wZdWWVPgxCDhCq9IgKh1bAVXS
FbqD4ZlFoDkUB9sM4TE0AKwEoh2sd54uyCzN4UXiGF6jud8wRS7A3N7mc8maGZ0b
D1j2BSNkRlNfW4ZYZANNbeewdX9z0rTqYk1znm7KYZzE/v5JTQa5HajT45kFzp+h
AE5Esag3cKcucrMnCtstmKC3QHiG7OxGveJ4SR9iHEdNbxPJ04bHbC9XCCtAt3rn
CqBOFLooTPCahLuhdH7AU4smB/NxPxn0ez07IpjB6Ko69RZm4JKTtjoIKAXq5aZn
sh//PXy6OCOV7cd8Dgo0dDc/+Oid77j9U75t6tZJQBCJ75x6oCpfpVFtYbr5ibiV
P+vt48UvlXAYQZnbnDy5JJHKAshq7n2Zd/uc//EkzWJUcJ1MgAqYjePUACWG5TFx
aek9HoORyPvoZqGvzQZ/NPl+/k+5dJ34hcjw7Z31fQFov04CJiqXeRl73YcSy0FW
af2RkKkA1PbzX1WDnl8qRxLk1Y0tuPp2THy8AvlZOlPfHQc222nnZgchBzh2/aVI
1CS811wWj8XA3bx4CLBDQVSwog8OdgGFxX9F4NrFdJF28q0qfMpIt39m8022rxRh
MO8AiE4ScnvpHvCjnWYAsgieAh+CCM89PEm1vdBLPoORjxBp1rXOGF3eKPWILkqM
PDMn5KnZ4ERSG9hhuZYEWyUZgRp1byK1uTekbNUerpnruVh25MO+jOY2tHs2WdMz
myTzP3xXyd++jYs9ZoImQFesBES5mEE7p2tlrEhnK3nNSFW9sZznD73hVeQKzndC
78U9ob2DXqUr/wsMC61tDgQ3JiTrokfb1xObxULuo6cmi0j3AroCHr2rIFjEPxGJ
Uu0VtZOMJrop38mRFGfLCUYmlhXeB9HVNompKO+mdw3JcUEp5C/VPQUhd5t4E3K3
p5c7P38xddJDT9bi3CRGC1b4nRp+cCfgkScZ0QXn7C39Cg6UrOhEP2DHpAwJAEnS
KgxtJf/CDdNjmniVDCrZEo7LTJkvFYVVDxgQ/FDqh91AngbCUr9NuiSZDRlVkLEP
9G+Dc5Qfd5jkmjJ9GZ9LgcX8iHQT4EwWh422dWHrZAtbfRSur9QATJ0irSaKanK3
h92mECMiryy5S6NKZ31rp4xgQ47xVxvUc/TUlIpv+DtARhSzbVFkqHw/kP5R2l1i
27/nPLRayw023yMrSAZTM3uZ3k2tQ6b4zgRnJnM6Jdd8NB9sZLLVbSCd/SQLNTsK
4xny5/t+3+vyuL6euEbZuQiv2xU4LzY8/JGLaGRPh7F77NlGaZ3kzsNXI3LYKXC7
oVf2fjYrf+8IXU7iRZ7YA1D3/8ujp4yINUdVKS+TBH9UNB8l8EbruzoyyydADltB
eIUd31koOpUhprmUeTJ3M8E1Mb/HonJ9DP3aYWR1pIBAyA+blOSd2XMWmV8V9dKS
6Fvkgx4luulsnvjXhPRNuHlhWepqaDFqc7ZYf1+Cdd56tYytgTdvoTcjMIvWZx0X
a6CzNq5EvdwNkEWM4QPh9GcJqIDYypZ8TAwu3lKLhgdhPqFseIVXUael31Clibm+
yatVgng83bXL7OEAOYJBguTv6OdoegSesX2sk2uQuULG3+El4SiXJXzBSKZEGPl1
AEaqPetgh1T1OGY11X/PUYerF8jgP9jyhBOhS0HC7M+MKatp1VhoNe5sAe/sAkdQ
gMGidwvYB+OZ0ptDac1avX3xG7389LOe8Nu5abs1mexQ9Z65BDwkf2JvuqJp62W3
wpqa3f5Ndsjsa+8V4FSt9zgZTqZzlmGT0BdF5e2ue9F9uiztZPdP6+ilSOf8idq2
0BWEPm/SE8M5L9BJOS506y4+LTBttoDkj/Q/DQQIlQZ5T1whXXojNXvuvmnyP+6M
p7GzRFB/P8rMWG1daHtLxvab0swTp7xYwRR7cHSAel4buK8ne6sMMOycazP1VOb9
OkjFtI/LGXMHtEjffOBS7UgRXWt8ZmTJmdXiG2ljBegBDDHCaiEctfZao+xzlBTV
klYUsSSSnPXbBXQHQusjR2x2lwe+O2b4HQ8FWvVMomYsfPl2yIGXlCTtcnNMT8jr
Xiyn1lKSKRBzSjTs1EO4bX33qjrhJdpQ14k9Ti95y1dGNxX97BnixAbnuXioU/Sb
hd0mYzrgW6TrjHmzmcbUq6YXv8dEkvRXj80/+QEZuLLrVovBajh07Gf8uwQXnzTz
8GqmG3izhTOHflaWqzkrDrfzbmI/zP0f+29L+z9O49St626A/vnijQ97hIvo2D5a
xTaBbn/2yFLzyZCOyaKEZqxwWljrHza0wWXZWnM4O4R+cXg41Zu071jwGl+RMVb8
CSiDNW0ExT89pqZCcqFohJfaLgc0QH/dur1DTWLf0qtWfyEZS3bUNzg/My9VK1d1
XwgrxCbnbNURy8PYC7bqJfexqm1Q6ir6C0pbvenV49XZH76vazGNtEdTXx21thry
W0VUEnz+x8/XWEIyfAs/eL5eYCMnhTqGNBufvlvJCij4GGF2N2/bHDJgSYkk6b3m
+upp6cfaZ1W4r2H6PDJxfgrMN6/cteh4+pmgzXxuSKOyruoiq4LjIJpTUW2WOcfC
WtVpBtpFHrfAwG9pWSQZD43olLBS/Ccbx5csa3XAMiwHtPvIjKkNlCdjnBrdqCcP
araybwy2VySDGOplmB2IJyYJH4kbq36n8N1rhP5XIb8ZIj2eOsQCQyDG2bZhOcT1
pFXH7axcOk88GhLhkgY79xx3KmCX7HXovTjoogES+of88lMp5myIpAzIuLExVN4i
miUVSUap8J4JvbRiPUgOZm6e6bMAXGqlAnBUlZbqoxa3+f3wXwzfKbReQUUhefBS
VsEsPq4sxrIZFxJ/89nipNLwtv/z5V30mEx7/K042Vvw8mUk5rWAXXrUz73TxuoL
6E/HQL7w83xqo9ON+F/4LPsY6WtJ+fLS2s3bp2MD1SitxdJ36/Jak6fuaUEVat9X
VRC6yeKjW6mkXLnpkLZBpjDHkqWslq7ekhcV+Nyxgp830x4LxyipAc63I9Aa7rUp
T5l6PfhRGxapI+/yhNub+Rpk66+L9ciWnRzUWCz6Mludtd/P+6oO7nWzczL4eU4Q
awuhVPR77T2007eby/imxdGc9/vG4MePS5qQatgUMF1fqZV+PpqtITWVvfZCUMXq
hQgBwq+GzEVA19EMGz4WWzFVUBMRGfiKxDdQk9zE127HviWXVrrCCxEiGyyZO1lI
17RJa5BdzMqqDNN8lMyDv16gG0y+aPFxXRY8fDoTWcLWsfQw6xMfCwXY+GIje0ES
Raqgk5Hq1G6rNJXFNSZfz+zOTbCRxei9Bo024WhJmxVF5UxzLKt72O+1PYpooMFO
wiTXU++3rsbHAt3SuGI6gEuWiLbiDFKCHYzFho7hprFT7BetvxA6pGhHL6UNs8mG
a9eachq1qJ+GHB1VCK+217Sr3/vCWOrj2xu8o2xV6wIhWvZCHiMDRUQiaFrNGVnA
M0MzYSEPeJVyya0EwCYVQZShlw5i1bXYXDeIbYauk+9NwptVej0V21bcESVb7W5P
7YTNfRMhKGQJ5Tb9vosFiTftQPbJ9c7fhq4G60MAxHLe8bWbpbhREMbn5AQF3Yji
erXRgAoUu/0YoQ/Ey0x/qVZf0HeIxCc207fqAfdgo8yLuSG7HEUfxzhaiQ0w31Yi
CCPtDch7Trb2O2E/y0v77WsyXCf0gkLqljL3Qfv5WNetf0FntJXYmOQmnaBv5c1H
6+VZKa2D2XYjoywmFF9IT+91AWj0xCWnxEvhwafda1KbwHjoxr4dfB6WHES2xyoa
quFJlgJ8JDQUUiGTG0wNDZk+QfUAEW4GFFDdgLUwPXG7GcR2kez/6XsEXbKDwozg
lJW69+73EHnFUkyWGvCx/bGJWjY3pHfdRJjS9dDoyZmOE5BziAbMTaqRIBJqORWe
EnwG7g8sexHcByHzYUwHGpfNbs/i/WF02qWNLRDnYwH9UPfkyciq+GVgZ/5aUlwn
1zfe3cln9ckrUR/xqsaQJ7+v2Ud42uX98rzpVY5zfDT58A8ZL8sahienxeljbuqO
QuJL3h7xJqXFVtuPdoWYW4gvAHxOvX4qtpyA9rw5PRhm2uGsNPIbVngfo82sj3fJ
gLa9u5CE5sFfujdGmw9ek3RGLTAuKYeGa57acTK2dLy0HgQbio0FxO6CZFaDflNk
0GPBOYtRxSV21c81RJR5zOPKkusbhMoDEnRF4BqM0lWmv8QESyNgq0cGcCr+WTgX
Fa7OAfWVwWqoF2xG8DrAQS8X4SN0QxkKCAILsBILhsMRr1jD4XVHMiPv98s3rjPK
cEJj9bM7ldpRj4JZIfPyFd+zQoR5ln1RGpyIL+qzKF0aXo3WYW/1qlqDr9e5wL8x
bIkxL6Gl7OkbdjXcEL/P+KGMpHoSX2dQ2tbtZkDKO56TrUsdHpKCaO7eh7qLWJuu
Ko80viXCdfq7xkZXA476CWBGPFGdXztvjE7eSAEcuyJaKIyQqchG6I5rtX8qD6We
3GlLMfQ2SbwCiptukGwv5S2/twSD1t1zCDf2GWmq5L89S9Xzi3ZVMh2Qa/8hO2xl
wB9gv6u2U5Uy1Tc8eSYm/NWEI5UbO8cZRdS42t5XdionjPS/8XgcU4AGqD4BZL/a
VsUhR3VPYcHSe+ftUCQ0l7A72Igyh+2UatR6RCfTsMxKKWFOE9jO9fbxYjD4PaIS
zzwChgwSxeHMcemKRAL9AFcJIi2aPihsIqVYr6wzhNHaV1SQ/S0WNK75AJmr1IiW
c3rvPRtVXWS2vmhaMkuwQn30kvnJD49Wpj1uQloDnBMgTXyNL0t6VZZ2I3DaXPnh
/MbAnEUN0K3/KSwAorO+vi0Bo1i9iUyRf0Icui0KKBrai4ttSqUV1sOSfxZf9o9J
UhJ05BOurzbBjNuGHShbA4nSCFbwzu6dukD/4j3S4om7lG03IwTI/L1n2SXvGaS8
TuY0RotaXxnw40zn/AJjaakJMgy01UK4BuU37BixTJKXRYFEj4OkLYjb2QL0UO6y
V+gAMdGZw8x6vhyyHtqqCcBFdQT4fdWU4QoW9M1Rj27PruYStuZId3Y0AAinQkMi
sLq7lAD+xjoWu84pPk/2c/LZg6XvizRK0Ii2F7gWiiZkZVdvxE8/4KgOT1Mz+5a+
0vSf+gHCX/upo4SytPsgckPMsuhdE1JinOxLJ58J8TDSK8ibngl0tRkF2Ogxiv8h
lH/LmvHaPzjW9u/5yDAfmBR7t+zLyHbmUfMRc0lMnfr53m9MX+emsG0c9DMQojub
UsFgLSNJVDdD4q1FxotpsbYLG6p9nvzs3U6Ug6gpZDiKdnM3zDbkhOleEnqjSEsj
3pmBUlptOVhKV90nZNoLi2fZDQr6O2qqdbvVeAV+nC04S0Iv+5qcbcjW3vHDcJ05
KsNQFtey98MI2SXEXI8U9PAJM/s/fXY+KXY7H2/VpDOoZqHU1AMxW0PmsDvfGBqJ
MBp3OE8kUx9x4MnF91ZIGQ==
`pragma protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡j��-��l� �3Wʴ ��ȟs�/�\�Kڰ��n��T%���#f�� �J�R~�\�s�ז+�k��p��e�����q6w�c�WB#�=�����,�����x����u�K1��b�#����q�6j�;�l�|���1���ˬv\y U�Ԓ���e�u�O4�U��_�wL��O�12+������/p3f���{q�mj��I��F	��|�416(d��]�T?ϥ�c��7�%�m�SF�]\b�R�����ȴ^5uݕ����U�G=?�{�(;&��gF���E�eW��%?�ө�_���y�&�I zZԹ��0F<r)�r'&s@�O��"6�U��3���_˂R�W^F��[J�6��,[���`�����L�ؘ�Z.���l���x[X[H�Zr�p3�"��m�|�lid|��a7�y�@�֒H
�%���B;��d㏏N��OH!�v[����󮊳يZ���T�Ƌf	��\ڮyW���`Ӝ��wk��**v��k%����\"������vA:7R��%u��}rI�_����^,ܐ^�A�[����=+zI��6R�lP��RY�'���gݱ���pzV�C�mV1��k��z��Y��0A��W�x�l* kވ�7��Sx#��+4������^;�7J�g�3�"J�3��'��Yb�W3o�'y	�x�B�Mx�5��Wr�P.��\Q��v��˱/��ב���G������KR-���5�V9cOd�hu>��&R��[L�0��'g{9G�W������[Er
n^�V S,
uY�	(@�X�f ��F.]9�)���U`�|�J��PsT����P{] ���i�2���]�I*S��t!ZFbΤ�ogؗ�w?Q�ԇ$`���~g�,/n���]����b������wr@�ՠ/�i�餍^�#v�����0(,���%Ρ������:;o������Q鍦��B�^R5s�)�կ�����Wˊ���� ;ܮ����)d_X�"�܎qJ�-�1�1�_�s�9�#~��EB�J�km�F���of�����܌�B��}~�i�cڙ�#�]�ikL֟�p�wRߜ���������VC���^?<�/�*������,��D�B�om9�̎4,g��[_�R���>�+˅}��A%��_��Ļuw�gn����@��������\��=�Q�gQ�� �9�T�d�~f�9ʞ�o;�������g녮�܉�-��-�sf�JD��c�x�h�|x��\·�M9K�ϑ� �o��tN��c�vE���{�&�i�� 7)H':�9fz�FZ*�%є�N��*�dm��pJ=E(Jdu�N�z�	.�H�T�Tk�e2��Yz��e��V�Zd4-lhl���j���R^���d����Eao�Hq�Ƅ���8Ō�vU�FW�����e���۬3#Z�Υ��k#|iV0��h��)Q?��D�g�����Q�3�����Z-�索5��{]>��,rK��H��H�;P��j+�f��'ȴ!-�$Ї��?�U�Jm,;������X�ɻs ]��/�fV���g���q%��*��|��'���!�+>�i蜖)XN���QB������"��h�����$-��[/��*H�\vd��6@�:I�[:��MM�W����KWʑԚ�L�ua��"��DR��˹���u�Z�4�)A�kf����0��
zԌ�߮�-�\���[�*�(�sOC(�
�L�߿��knw��[1.0�/s"��`��a�4��TbO��w@|^N��v\������ˡF��##���q��H���.%l���Q}�|�kB�DUV�B��)�+�=�ApKCW��שr��L�Q�����ʶ��i�]{%�
��[r&0��Q��w/71{Z_$�$��"�H?���wޯ�q���/L��A�'r�e�4I%��L�*���Ιߖ�p	��Z]����_���5y���ۈK��Q)�c�C9� 0�+!����U��(.���.ｏ����UPǣU�O�
�p��SZ̯��.�%��~pP;�ԙ�����ِ�R�=��>�H�q(q��u�~�"y�~�k�㨔��h�D����>F��}�-�Ce���q�jp�2 �}�D�`�c`��2�|�'��J��.�Q�fk��x�8E�EN-���D�H[��;%���qE{o�3��5���j�&�_�"������	*M���S�/����N@0�!�8����|�*Y���=�:���q�Y�:�K{~������͊)�Ky�Lh{�N�=����Hf/�ȻBW����o�$ϾY���RU�d)z�𢫧7G{ªV����R"᷐r��r0*�L��*����"?�%�/����w�8�Y�kW�jaTi��+�o������� �����pz
�W�f�v,�I���6�b$��!l�RO ��u��C~Gq�	��:��(><F<�?e�G�Y��$2/�����|�&��FP�s\I�w1�6g�u!D��v�N|��bKxaCy�M�^_�s���m�I���nSWIKK~9�(�,�v���4p.���uy��p�lV!����6|�G�$K �W���C��b�	c��	�٪:#�O:��'>��p���D���p	�υ|6m�yKRX�D��I��߼�Ip�8���@��i���<vEʒN�>l<�B ��k$�e���6��Ϩ�fb>�;H]ɔ3y�6��ӷ�ou�Yu�֫�u�BMvO����(����O�H/��$�wZ���ύzq7����̗�+Yu�yg;�8�Qn��'V�k�1����}�+�.�G꫗��F� R-�Q��@�9۲���͋��С(����UB�Z�e�|����qN(� �F�qq!N���	ʕI�� �W�P��|�f,b}��	`^ѽ�dbPcQ�~\���Ǐ�?UN�������?v��f��u��3�IF-��A�Nɶ$�����1�Z?1���1��A�5I'��>ceĨ&&��k�y��;RS�)#"�7��g��%L9?)��(�2&#ϙ��/�6h�kq�n�o������)�����N �/�>Lׄrx��������V>w4���T��^6fy4�b���z���b~�~#xhΟ*%����D�)m��
��E��2D����١h���Ye��(=�	E@����RZ�(i�B	�q%���<�h��!��b�S���T����8�����
��%���6�~#�6m����I�,|�~�:�(���ڮ�D�:�@H7�0�r6�c�;�M
��
l@��n��U~�k����v��� ��uW��Q�D=>�zw|ۣ����'n���=�{yּ��Y}	�B|oT��P�g峐�����[g�Q^������P�:>3>`6�� ,?;C�@�gο�9�kT�Kl	�gU�,�3Z�QrԔ�� V���t�_�I27HAR=�����̽�'��I.>�	��d��D�2���D۩�P�����[�i>G���}Cn�X��K�[ 0�V��O�cBi����8�g͔֞�C�~oG�+���G Ғ/}U�?���k��rC��jC�2�D+�t���*7l��)�QMd�\���v�u�f�=���n���y*+#a��b�:uD�$���eSP՗�V�B��7bz�E��l#E%����W��� �#O������	�c}�/��+&l*�^~Y�_n>J�/=U.!4��^����"��。�7|&��[dAWAD����t�2��"����d[4v>Ă�����n����]��?��5�P f��t��Y��<�U���d(ۣ���X{|��1x�	o�jt�rKCk��Ե����\]����S�P��J�</�P(��qab2a����L�R��?(�|�|F�Ri�r�omZ�L�"sY0s+�a�Զ��5��*\�����g[L�U�D֜�3��*U��{�q�'4�+`���j��IE�z�c�LŶ�E00uU��>�yʼ�p��.�V3�B�yݭ^<�u��Q�z��b��1a�/����8��G�X'ݨ+�4�+?�"��k�i���C��o%�>Is{H���]����;�ur	%��ӥ���e��ԓ4�?��3��I_��8�7#���T�P��6q���zĉ����t�+���d�0�����`����|I(�C�fT*� h9rh3|�@����+��{�!�k�49�S\�d�*^Ph�?����O�j��c!v���y(��d�L��Q��I�z7��v�=��%:��n�}�����˦���T��#�m�핺(�7���c*��O��a����j�T�+��W�a��r�V"ٹ�UY|�����n�9���&�+�:�t������EOU�]�Z�l��j�&R�F_W`T��@��&P̦�۹g^��z�wLk����c�b0����';Ñ�r���t�la{ܭ٘V��7W[��B�\�k���ى�'�صLC�i�+���/L��^]X��۬Y������{�}:�αĸ��_��fo$�$���mt���ް�)}�;$�T8r����e^1V��<�=l��J1�AlA����ȿ]�mC�"�	8\��ݚu_P�d�&z=?�m(�����ai�����\�h��Xo5!*'\ԓh����S�6��5��_)�Aw�}��u��j:먜��
�m`����v�G(�(�h�-�ȿT���wց'Hj3޸F��¹�u�*	T�H� B8��P��N�R�c�ۉ�1���	[����ʗoD�XY��^Ɍy�kߴ��d�&Xf�7(��Zr����36T�s��U�*������W&�K��P�m��u�œ���^�>�����PY�S���J�s+}�f�o�Bd�,�"�r��W���`:��ؓ{ɇH�h�k��5��̴�`p/��&�R6-2y<����(ul�@қW3V�qd���G��6�*�{ �'�����]�^��hi�N��`h�f#BMja�a����3&0[ѿ"��{P%학YI|��'b����9����(����J��ӎHڄ+��)��ױ���6.�����&;\�\>�'�{_JK��"q,(j�����!�,�@��4�F:�޼׌΄���� �������>�=Hb1��N���sI_��Qߛёi��e�OM@��n�?G��6O�ǐ�����5%��ߺ1�HS@�:�\�{�h���������Ϗ̞b�����U��F���k]7�!,k�ꉹ�8-��V��.�J�rP2\;����9%А�M6��jzS�#5������m+��Ĥ�t�X�p�
����MgW_��m��2n�!Mj������J��ś��i`{��>��WV�u���~��f<㱴Ć'��}���s�����蔑�ڻ�8É��_���O2ꋕR��Yg�LH�X���"���'Dt�{SE�ڂ	�$޵`P^���i�%2�mݳl<-���P�����>p~��X��O9���N�G
�+4 � �4f��I��~z��Vn Fۆ��~�U@�~�ǅS�՞��lq�W{Y��akl�'Xݣ�@���?DCM*��6�_�k��Н��1�%�Y�@��NO�2�>���k��VT�����5x��BKM���hl=�("VRې��9y@��d�Zv�$��3���8�Gp�1�|�r#��뺽"����rF��������A?���ܤm�B?��uzI���3�=R���4T8�����p�f�ߩ�>NIf�k&��`�S��2��{e�Ho�/m+7,�"��]@Ub�5���V��04��tV)vȴQ%;�+I�b��U ��}�u��#l�:��_��T��2���ou$�.X�>Ơ�[�5��2l8��:#�u��n9)h�q���+�?����x=O�J�����Q����d�P�����>"�rq!�ǵ�ٴC�q:r:_�̆��� ��*bOs�/i��Y&�II[�fp��xi�b�����.M3w����l0��J��͂!f� q��л����+������X]/MDъ�]��[mXOг� �@�6$�L�$���c��R(ν.Ŗ)���@}&�A�)̻��ew�f�
�F�H��k�b�~	�Q�@v���*�%��[=�d(�EǶ'��
��wW|Ј�$�l����:v0�U�Nhl��:�,bҖ�����/�ac����7�ܕ�&FaE%��)��p��ѡ8r������GvGgOG���G@�[m���fDvf}�ǘQ�d*ΜN��Xg�7��O���#X5�L�7JԱ�@#�QU����xߡ��\�?��I�!i�^�C�*]nY@��ݞ���l��%����ZD'p%�Ϯ����
�.�{v���m��I7�"��o�Pr���zh�%�[BaƲ�Ԅ�ϊ.tI��w�d	r��wÔj�d;�s�dĲ 6H�w�۷�Pxp�>kZ�1Ơ���t���wNA�V�.TAZm )W��(	��W��D�3�/U]��yF��7�c��%(ٷ%fI�S[g����eL�[�3$�/��h}&M�4�O���[��Y�����W(�mv�d��8�f3�zf�Ѥ��J��]wF߬FC�n�R'�����[Q��\�=���>A��y)��u�Š���n�����T��?E+���&���K��X��'N�警~
��~�45ի����C=�;"�
���o�!`�c�M�ڏky�:�mu�,Ғ�\p�J����r���=��QQ�@�tO������Y�8e�ݕEX���%�>�]��e}�t��Q#
o���֏([r�|*��IKߪ3�_���j�l����z@YD�o�6��_/dg'��ul��k����W0�x�z�G���0%�b�`$��x��OB����䑬�Z��O�K������97��=�ik���c؜�5l���d�׌�|�~��-�(���wD_o򦼾ϧ=�5����EjqJ��i��y��oلL�
R�O���w����9H�f���	.�~xG�!9�l[�huHPt�I(̺���}I�M�i��.�n�SѠ`�Dh<�Z��uF���|T��
�@=�]���tD�����dҎ��.P�����䪛��^�Î�����gEt�4��@���w����mp�q3�$�D�:^4�φcl.��6���F���l${V�2c�m�{���
�H��	�:��y�Y.ꂝUH�:G���������v+�Ȼ�BP�5���n��"�d^�/��i�0���gB���>$ӛ��H��4/�
X�(�E�gb~J0I�)���F\	����c'�֔�&F㶏xPe�0�a0��O����V[�(gՒ��oz9�>M�w�|���;��s���{�n�$q�A�@��]"���4�O,��A�6�w��+;���j�"�,�ք�x���?L��YP�715pI�Q��[:]G�:{)���u(�n�"�vj�թ�5�j��Z5	�3�n����	��>���6���q���_j����c8r\
(L�WI$��S|4�/)�P����m������	��cRɨ#鴢r�#�W�c3�x�gMP󍀮6~%�.��!��ܪ.+���P��,��È��|b��<�+�Z���9瞕G��q������ж��Ɗ&�"����[iK��'������&�.z[��S��*�,Ba@�l�~��UƩb�iN9�,�e�2
�D�Aߒ���[��!b���8�o���򘻄,�ٕ�������x~픣��ԉm�q$�p�*�7SY��������K̉[�#��N/�έ�9Y��<�������"��pE�F�R ������KF}#)��lݩs��yV8tWGNLS_���Q\����Ink�#˱�����W:��sN= �pi}Ȉb�ḅ�(���'�0uj����b9x��mR(V�'Kk*������~�ɶ�ǝ�RSBbEa�Ϲ	^��v'� F�+Q��Pm#Pt�E��mZjW�$����4]�J[j?��_Նu��	�&��+&�v>���2M�'4�&Q���U"����W���a�=��o\��oX�G�qy�V#(��o �&�\k�
�Kp`����0Q[��J/�{��b�T�@�&̤�ܒ��:sK��kj&�J_��#�~�N�"=��kX+�������|��9���N[�rM��;"�"^?9׺3�NZu��$����y��w�
�R%=k^���ꒃ����"��b�@���_������)H�� �	�`�.�E�A;԰�[�n#e�-���D����5;�N�-��������h���CȈC9��f�D�D���Q�����e����\sL8���,�?v�[e�hv\s��N�2*ê�2#�����@fv�5��1Z��o ������H�<�׾�A��G�f9HhZ�������ߐW��Ą�9��5b�I8��y�V> ���������-�DOOwXɄ��1>�z����{A�>l��Ļz����*�¥��h�kBxΙz���Y�l�y�p�MB멥�hZv��k�ϽI.�c�nd
]?>s�PO�Iz���mٱQ,��ˎ��k�׼`��}br���u��{��q����"�R?���4.�.c[K{�����;Տ%�������	_��o�c�� �Dʴ��� �qũ[���.Ou;��
�eO���X.@�G�*�B�(�9_k�%��Pw�ܚ�>�qH5@N�N&�_�Zuu�J�c.Lw�%T��7��\%�Mf�Dk7�ʹ1"h	&����4�҄:t�ⷎ�'v�H�4�ha5���ju��4�����~�y��5)�-�#Y�� *��`7�y�S�i�yƫc�F����
2�i��B�t�;IhظJ*?�i)���E��	�,7�`��87�$�ŗ��L�.��k%3�� 3��b&=.VO�����`d����c�b���ێu&��;���W��П�v������R�֬V�>8�?m����X[��r�"��5l�}Q��wY3��(��m��z*m�u�Ӳ
im%��"��,~lC^�z��"��<��<�|�w4��Y�6X��@����u�0*Ű=��>�%Q��I��e���>`�r��D��?z�q[H�nθ��h��0�Z��|�:+ �8��V����@9����d�S�x,C����M�%��=[ZB�k�=�?�C<C���� ���?P��uc�һ��^<�K��NdZ�8�^�JO�@D��Ҟ�X��X�0�i2�yc�1���-焮&.U�=�����M}/�-��Rθ�ʞչv"����67������;1-i�Ŕ��2MJlC ���>-zwi�ƈm|)���ķ�tR��p]4�.�y������D$�öGD�M���jS,�|̮ICB�Bj]^�U)K3Q!^X!�K�u����=fC��''+����L�V�f�o��:���8a�˩���4���D��)���ڦ�!	I]?V�n�p;�[��`�m����~�*W�F����"񪼦�4"C�B�2�K�o*��㛛�Xӳ�D�I�V��=�3��W{�N�����=/���F���>�,� 	G���:r7m��+�����z�k��JI��rn��� |�����pP4pO�dr��èN��ʼq�݉�G�P����2i?��}�eV�L��Z�N�M;s���-Bfoc+Θ��[��̌�X�:�5��8X%O���tqԳ�o��7�.�d����%�#Vf�LQ8x��"{B�;�_�����1�#�I_ ��lT��`}Ρe1w�(��,|p�?�/:"e&	x�/~�k,�����/���B`	�į@��I�CzV����3�.HL��YfE����_�Kw�V�f��&k<�W��ޞ���bP�G�U��ӯ��Rd&4W����6K��X�|0�a�*Ho(ё\����f`}oS?��4�Ts��`/��w-B�	������<���+<8��l1U��㟯q �Q���Cທ���"��"�ґ��X9��Oڡ>G}$=�c<���[b�#kLޫmfzd�$�{��)��V������m>I�7`�)\���`XB)��)�Z�t�7G�c�6m/ҸrwW�|O��{�aŧD��rF
p/+��hJ����t�ቭ[G����2+��*
�O����q gl�t��Hz/�@�2w3p>�V��6w)ˈ��`�; �8Sa��
�=i,y'�sugyt���iӪ��f6k����(��m�1���Y}X]�|b��I��?�=�+Yp,���>@���p`��;v��i`{��B��C\}O�z82-bx��oW�Rڵ@������������ӥ��F���'Ȍ�3�C�a���*C7y�����17-�'l8{��ktB�ſ���DgŏM�H]f^ta�͗V#�yv ��sfT��֢�E#;��]�5�v�Q����0��O��d|� �W'k!�&`�3q��s��º�8���.�[�%N�	
��:����/ɩ���ّ��L'.��u� N��DڹX�2�� (f�Į.Q��Y�f���ۗ�� C�9#{�
3���Tۆ��'��.N�.��
.�dDښ|f�k��ځA6����U1����x/�.ok(3�2��Ym�~oA.r�˴A�P�ūy�G9w+h �e]릉����#���M��<=��P�o���Ǐ+�+���k��8��L�г3��н����_F��SK�t��#(��V�Ry�ak�/L3{�����S�[��;�%.v��,T~�����q�` e|�g�w�Ҏ�mm&�Գs�%��%&ar ��)?q��CCc_tՔ�h8�z�$@�����&�1N�]��My���0n1��\�;�#�۩�a�м���\���kF�J��|~>�p9YUW;�XrXp���{�ծ_��E�X-�m��S� ����C[�4@�p?������1?��Zx��O ��l��J�wA�2HSk�F�F�G��9t&C���d���M .��C��e �Vy��9�8��
�z���S�����Ͼ���p�2��F��_�~oC=u�=0����F�1f��G�Rz�	�:}\�ܦ�q��������~H�Q�v�~��i-� �d�S:M	��(����E�|��("��<�CΏ�.h�J63�}W1~��-c��kc�@�0�^M�i�X���H�*6�㙽-��h[��;]�]��ȣ\��ڣ��Us�H:�m?"��Q�aϋXXR�pi��:B�.�h��dN�����)�� tś!�ue}w�g0�p�A�n���+���@����Uv���"x�pTً1Z�x���"}���S����QZ���@:|���"Wٞa=$�J6�8*'r��u��^l��
�,�
�Uڒޘ���-�pP��pΧ۱�����JɗZb�!�����h�ج'Ӡ��QX���x� {=Ϲk#&W|Փ��޲.
��zyæJ�r�}/��ywB������z����_1@a�$oV�C޵����C̹��Q�Cw�C�b��e��N�9}��ʷ��f������bj>F~��������eAY�D�NԐ����E@֋��OX#�G"{/3 ��(K�3�1V*F�iBrq��!��K�4���SD�@���� İo�j\]�n��|_ǰ��J9
c�~�ڲ��S3 _���:z'��L*��ө����u6��`2l���Uښ��N��ș*�'�e�L0�*���Z׀�<bH:_��ٷ�A�)�G���Pk�_�N�]���4ν�D!i�J�X5��xXRw�Cłw�t(�6���K�yr�Q� ���8������0�3̵�aK�%z�.�)���g�V,�lAk��� ��Nc��ױ�汄�9,O�Η�-2g)����E�q^���K�֘`m��[��	�����yA��p[�fz��������QTIh;�/���|��#{�M.h���[R<8x�t�_C���b��'�bn;?+={���:�@��t�%-�QEz�a�v��}�<�jP�d:��2�2N	��\<W�r٫$qj��Y�����
�@J��+�jl�!ϡ�\$?���J����g"͈!MD��c����o�t5&ϭE�k�=���N�n��k��!����a=���YI�|�[�Ym7���]�%��ZJ�����,o�g�l�au�VGm[I�����E��@¨H�`h�[Ⱥ�l��cS���F���b���m���Nm+��Ov �-^��=��$N�<d�B0[zx�KcIhI�q|Y��I+�v��ԥ�5/hhʧ��;��(�b��>[Ja.���N�����&+��{����G�B�kp}�9^��!_hcO���	�����`�5���=�@թL?����f-�N�����K�`�϶{�,�j�貤�pO
�V�juWf+�.�ٸ^�
,��Z�=@��i���9�a4��Ttl�P�h��"oHPy��B3;��@��cSr�s��P&BP�L�&��{�l��O�a�qN�"?I�d��x��q7e�k���鋙�zo��0c����B���.�P�W���i��Q6�Z�>��Z�w�C�~�+J'ǧS��EA�^��u�(l�=�gRѯ�Kֹ6���򖒁`�Mp7�c[��r�9�_؁�R�h�
�@b�7?H#s����׫*����:ņ���ݜ���^���YO�\���SX�� �N�Vx�Iv;��kyϵ���| �eJB�^�,�n14���Z3%y=L�QUo8Ҿ|re�� ����c�AD %�B�m6��G��]S5�.��o{��r1�KpB�t!�� �t6[���H�|� N�V�H0;Q����5�c7�UczLR�b;���+}Wg\q�L�f�߻r%��, w�{�辉�#/w��
<��a�O�uï��Tb��|U���{�dTl�����7P�����6f6���5uI��u�����վǡ
�(�>᩷_5�Д���x�y��N����|n{F"�$��/�o���>O��ٷ>�N}���:�dJ@ � �4�� ���[Ծy��]� �G���5�7Y����U�v&��^�֔�Ju�.����?+F���Y�a�Jb27�=t�*�R�ə!�(GH���Ce���H�+�����S�ea�]B8���Q��I���B�����I�#�Z
����;���ݺ��p{��?��f���ߐ�dH��ꤒb����Y�57�Oע��бp�AƃR�l�\w*� n�[��_j;O�l����&�V���-��[��O����
O�f�-���^�(����/��e��,�d� ���BfIFI��ż-���X]{b{$�g��VR�*^?�yRSX�f�"	�[��{�2�$T�q�%r�N2��mC����ˏ�������l����A���a|�+H^����]�6o�8��\ �I����^������0��nMX�!Ҫb*�Jqk�������/5���a�>�?����5ܗӮ���.��>AF��$co��V��[�f��(���+����b�<#��Y-g�n��[b�j��`֦����-�!��h[�!�Ax���,�:�[W���0����ȀÆ�̇~^`�JT2�,�c��h�(p����IC���<�6l��K��H���Q�B .��0Ǒ0��&����Ą�N��n�U&�94�=Y+�o��&uvI�IH����'@�!մ�b���o
4��g���4ɟN�e��`�}�\a\�ѿ]m&�#S���s�OC�NQ��+�v�l�K�V��R��?��#G���k��akv ev���x�8L��G�#���/ʖ�hB���v�3�U]u�K� �Ԣ{��(2��7k*�s!$e]�a�5�zl]�y7�]tɱ=�GSJ �7{ڌ���o̱�EvD �!]�fv��f� _��D;���_i��ʍ�
�	��򉒑��Bq>�6|QeZ-�����l�5��޳;1��>]��Xl�?<l�ӊ{N�N�a���P�|�' ���,��ަ�+�*4�6ʂ���H�d��(YB��\�B���(����z�%V�;�[8ޖ��.��͖��ڈ-���0���L���&�'��*�b��vhm�1,A�	W�?yܳ�=bCb�݅��k�����# ��Q��8�X��*S-1P�8L/	��[�5��J���ҷ&�:Q/,@�ؕ!�*S�ܫ�)E��|�>D��%�!�zw+�ߍλ����C�����+�?T��Ԁ�Ԓ5.���F`c��}Z�����}�ی�w6P��贤�	���$.��ӿ�/#���*�0�t7-�5;Ƨi.�t���c!��5���|��o���W�m���G��e,���BºJt�f\� �-ޯ;��˃���*���3�C�	�i�����F�4�C��
{cQeZ$��3J�'|6ʅ���P���N!�/$X��:�����m��5}5�-ʑ��בC�]�{��J=&�{왊0H���4U��`RSF��!�Sf'e��t�6��!��0��iu1�Ո��ȑ:�@቗�l�Fs�����Y\�5�9��sT�ۨ��'Fj�Q��i�/�}��W	d2w��C��'k��ܝ.�B�Sg� ����u��<�/F}����5Sw���`�	A���>�~��g�� !+�^]�ߥ:ڱ�����B\����I�6���� ���2S��W��C+H�i�E�u8ώ1�.W$�2�&��^$��8��x[�vr1�" M6^�]j�Bv�_a2Z�i��,e�W�]����Ƨ�r-�?����Bl��"Ͳ=/�r~DZ ��@�������W��'���l�qv3�˹����G�pE�d�"�$��Q����|F�6�wo��r��s�o���;C�Z���0���BC���0/#},�����+�^Y�v��M�-�6���Y���O��wEݢ��e}783�Ƨ�c
9�Z��i�l�u��v�%�!���J�(n�.�����1����H��S�$b��i�e��������s��Wa%�-eTY���t�R�[�ѽ���#8��{�)`��VZ:���Mvh�4q��A?�x�����x3e'p�?.sF��$2�)'kɯ�R6%�]E����{KFX?�L�8�M��r�*�*�/�E���9��C�_�Fŭ6M?�G�u/�D�Z�?ST=��c��U���1���6�H�JK��D(�L��,�:5ݠ�� 
C�,���)8�*C	����Q��*0ֹ���N��G����Òd��sO
��@�w���`_�j�(�d<�K�
���X�����}Fh���!��"����:���С��'}j��V�D�澠橦��X5��Vt�i�b6p�97�:o'��(K�_3�_6졧����)�`�0JX�n���Hp�nP�?#s��B��������4F�Yc�\}/;y8��[������#�<� 4�Sv�}��6�"��?��E��� }�
�^o��U���^��]�*P�{����j��%�Ɩp;�� ��&��PL;qƊ�{���I@��`��y�=�k��"�f�?���:����Y ���E-V#�vx���c�n u&������8�����38�h�'F/i��L�q�u��+Qcj(��1a�!�ƹ?&�KC1%��)�ڧ�wr��l7���8��/� �h�{��NNE��ľ��nBVN���\��+���V\���2{}��۷' ��Ky>��]�u��ź/{ߍ�sqTLG�.:!��[�nR���P�7J�i&p�L�Q�xH����pf﮾\�X�ߊ�ʚ�E	����lv�I9��B��Oc�1DU����\U 7��V62����E��B��ۅ2Mp�a�g��p�eb[�����gJ}T�t�Y�wCȶ�ӳC���9�� ���vF�ڠn4~ab�N尞W�d���K�6�c "v�x8ddδ+)�&�@Q7i�6*�M�)�u�����h�p��@�R�Db����Z� �OD7S8s���o�i5H��yuts2~�-���0��]��B~j̙A���X���d����cz�OU͘�
���"�p�.����������%��֡��C�='���i\mD~�v��_���"���;4ؖ>W�	�6N�燯���5t3(S�]t7�d#�z�pނ�b�:w)�i��ʲ|_���|���{l�[���i]qAS��ɣ�<>�&p9P��}����;���R0� �zN�f}�C
���JR���_����?WPUڑ��]11���Ĕŷ�KH�ny��ܷ�ڪ�$��+���HH�ڔIŶ@��ek�� +}�����v�;���-�I2�*�T����h�!�Ŋ�(�ű�Ɖ�V�'z0C�U�� $��T���W�
nr']��f&}G�H��:nlsIDJ���">����萫s�.�Sͤ1����k�;8G��*��67鏰[列?��F���O�a��쉘��&�O=%_�1�6���
�7Bkz�I��� c�_������Wo�˶�I��~��57��wb�_5+�Ч/��-|P���%ݕ��ύ+S��]Z�M��>M�9Hf��a��		�����&��&�ŻSm��
�>MXq��r�xS0W+q?}V��=��_�>@�e���D��+y'Vś�ǖT�>g��)GS�b�[-)��ؚ�J�ff9��D���MQ������N��b�q��ǣLG]���vw:������X����7`�?�%	f�CІ�3I'C��y�����Ay7*I��x��gf�*PK0��C�[< s��c���Yqe�O��ɭ��\H�t_�)G	=(�!^j�e��GVP
挑߅����F��������5R��n�8�0�,��/a�S�T�䬔D�N�#<�C��d��Dv���\�Ǚ���t*~."�%Ʌ��&WFP#t$���$�,Ct�n�-a�E�����!��Q���$�u�<�v�ۏ��t�/���޿�sG����_��rH�W���g)�B�"�%Փ~u�d���+�DQ7�Z�!1��>�GW��|&o�f}���Я� ���w�TB�B����{�jaWz>�R�#��ɵ��P@�����̟��JQئ\�^�xЄ�\����DS�S+@.+��\W11>[I�ڥI��G��
B��&p!ɶ�M	�0����lU��K7�߰^uwJIb�Y�1�*`f0��I�ٲj;T�
^��dĚ�Q#�H������RU~XGZ��v��ێ򢬖�~O��&��Jk�-��<�;��.X�M�$p�{�'%���[��mRAfP�S�*͑�̼�O���%����W�[������^kB����%UӏU�~��>�Ra4�E�h�����EpSJ�))09�k�6k��^�ϨE[vuz7_ԇ����msá}`���}U�o]��t�lgb��1[th
� �n��5;sC�g �G���4���`�ލ����B:=.#R��8��$cRH�A9� ���0;�ۦ���� ]��ظ�<������v=�j�R��N��5=s�;oi=��{�0ˑ�@U� +��Ӱr*�g��2p��B������7�T흷N�)թ�5�ߟ5����adP�[��O="5��]�-�L]r�`���SZ��3�Ï��4�t�A���q7"��9�|�hٴ�%]��q׸����;�"�p, ?R��	k#>�غ���Mzkw��Ղ�S�T���슛k��G����+%�Eu
6�h�Ts����o$k�+ʳ�濸F+���h�=��Рw�6��o;Cf�˒uÕ#d&�%$�&J����gչ�Z�zj�dkK�����|f	�@~^ޜLZw����~����a�,\մ�<	Eİz���z{ʢ%B���=�x�8�gS5l�IR-�DQ..�!s�-J^�V8�Ye���+��� ��7�� ��$�������$
I��;����jAU� 7� R%���ы���	�W�P�(cq���뼆L[�����+C<@Y=
{g�0��s+Ί<dP�!�/��
)~�PZa���9���;�}���@�-=SoU��E_�k� ��S��ur0�#�i+p6D%!����?,$E7�������MKZuYy�T��
�c��Śe��P��k����\�&'|x�,\�Q�}�/LL�9��N��8w4T
�#�^���p|�k�k+��~}��(|������F	�Y5���7&PN
[�n�b��^����P�^N�F�����BN��C��Ǣ݂࣊X�;}-�/lZoݞ�:%�p�-h]��;��k�t���~�٪���x�1�u��إ�`CU�����n�w������n�Y��C$]�hz��oRu���n	L�JC��ƈ�sx�,xS����(qg��7�c�M>9����R�AE��GiܰP�S������ԁ~�\Ri-rKf�:c�dٺ�,�![1�Y���Z�07y�z��羪T@��h�,ڳ����`g��X&�5I��8u�)i��>��M��_�O�m�����m�J��Y�iJ0�4'�P��m��@/��S���hj�v�r�i�I�Of�� �"�Z��hMƘM�D��KJ5�	Wd�Ɲ�f.?�C��Kv}wgálw�,��Χ��{�xG�<SW���!]�s���b��m�y}>Y�UՋ����^v֗���U��0��6��z�v	fF����;Vc¥�Tڵ �S)����8�*�ztR���mW�諗#X�@+(���T�H�F�Z䫧�@�\֞���e��h�u��;����j���I���P�#<��\e\������K�.#��r� �.fB#' �#ג�(5���o'�j-x��j��b���9����q)��R���y��y��7�~y�ۦ��������]�H�ྙ@�d�Lɋ����1(��F<��Ah��r�2q�7�����1/�ՙ�SB��iňU��m(r�T�kϱ�����|e���vsTl]�,��!\Uj��x3D�j�Mf+Y�����}f����A�r���=�+�.���x�|���y��Dg�VvГ�z��2}�5��'�5sԉ�sm��m�A����/��t	O#�rS��+�rN�"��B�&�9p�c�w,�r����}��X�?Z�:b!�OQ&�KP�mq8����O(�4��_�������v��x����s��|�^��q��7���pNw���L\v0�`W-Ɉ)�;#�&Q K\��ClaTط�k>������[�փ���4��P�����6�����}���^Xr3XXS��g��a\P9:�WɻDd|#��7h�V̘���#����X���^���W�������G:_l�=�'/������jw�p�GVJ �x��~��
(*MD��*:2<���x��	������m��N(Q���V�b�:8x^C9��:�<5;TT��QrL�2h ��_�,��f��#
��	퇝�~�!
0�b����p�	Ϋ�����`�r���E��A��5�KPyhCkUU�"G��CT�;y|]�z�oKn��nep�D�5 (9abUޏPJ�ԇ_�L���e��`/�(k),�ٴI3��2��3]s��Cd��:�,5���y���ɸ���V=%2q%�懴�G�<� NG~��+��f�lRq`�������#v@L�)%�S��r�^�dvPU; �1�w�J�����؆�F�++�^�kA p�AԒ/4R��3�:�=��r��u�4�.�l+���$ 4����}�zRfN�7htp�j��ö����L�93�����[k���	�<�~E��/���K��s>�
T��yɠ���,.C���)�hD����j(�߹�֚���vk^)+~�(�I.'��c�O��%#�D��x�\KSD���-��ϐl�k��bڬ8��g,��'2Zn)�ۮ��e[#d��Ǝ������ ���b��#�N2
(�PkC+,
E)�SAl����.#L��(��{̷��Bn{�\�,`�'Q��M3�C�bظw���ih}b�h��7_�%�-� �����gx{,p,���_��˕��h�5%��Bg��҄T�Y�Ř��ή�Pd�8�Z4e��WM48��2U��Ê���^5��1�~�~S�kC{Χ�ȿ�`�a�6}�q��x����4�`o�gt�91*W�O"�<hxJ��'���䵬�=��� ��z��?>�5a0�������˪����H3��Zy�c>����l�vf P��<88�)�x|5��Jk49�4��0Ǌ3����J�E��BU�O�-�0u��Xpt�=���І�⼫2�4]&�M��=W����	�����~�0�s�Q?e0wj��h@�C�@gл��V3Y��F���r�-j��i���:(A�`�6�@���0(��@���S3+�t�PB���������� �̑u|cg���>\P� �X,��
;\o�/��;��`�A�S�QyU���bW�6�!"\�d��"r�=�"Մ�2�8���$9�Z��_���fDDh:t��B���efO$��m�lM��7��^�^����:Q��8�Li��|�_'�~��D)�,��)��������0�`�O������`{p�{�&m���=����2I@~���7�KDO�5a���#�����a�5�}��
m�P�4>�Q�D��4D/��7���(�N,}�J��\@�g���st�L*0��r�w���"7-����3�M�Q���T9��L*�G��rwF����5Z��Zn�ڭ�\�f�T�Rw��Q/ʦ{�����3�=RE�C1�|H#��I��Ux "��8��1^,��^$i��=~g*� ���Р^���&�ǂC~��ǧ�F�a��.`'g6tٶ2q�㶚J.-|̡74s�.݀չ��0q�ȋY���N8(�����ӷ w��T|�U��p��mϱ�L�<��_�^�ǹ��#��[��V�����4����O�n|�Fd��� Si��:�c���0}O߉����k����a3����;�<gNlf�1	�OS"�j�φ��p��!��{�|����8x�t�tX�g��f�'�ܥ���$����fz�jY;�F�=X�+O��ge$Sޯ|���I�5�Z]���͔��5��Q����eZU�v~�F�Jp�9��ω)�Fd�0������sv�/B�멚��<��Q53s�b3^:P�T'���E�ؠ03��"���ʘX(�w`�����yB��&��!��^��6�8'���#�qIIV]�w�on��B��Ё @lv�7(� XS�n�������ig��C���%KË�V��E\
�p�ԕQ��~mL[���{���r��'�u�S?��j�a�ܝ~ �o��¨�u��������m]H�����E�L��zi؈�H#�����{�z����쿃1s �h��9�1Kе.)9<����4|2w!Oŋ�x�Oh�Z <�	B��!e-�ՙsy�^c)�B>3������#���E_"v��İ\���ns���,0HF��4�U�����٪�\eɍ���]�HF'Җ�o�cXt��wg��y�a�u`y���X�����Ho���ىb1+���ń�b�������>2;���L�Vۯ��%4�̷�����*(��5W��Aκ/xGc3�=і���(Kț�9@-��Y�}<>�}�l`_C̋F��nuYD9m���#b*D�p�)P�`o~���-�Z4�\�b�����$0�Z�� J����\�"�-Ú�el��Ÿ�%,1yp�@F��p�f��V��e�#���4��j�u��g��h�AX�zOɺb��U�����+]���W��7X�	��<8��l��a���;������"�B�'�����:j��ֿ׊����h{[�P��y6Bh{3�.��$�g	gl4��M��О���p1�/^�9���v�LWDj����!��R$鹲���4T��=<���E�/����!K?�ѥɱ����%eQߌ+���0[�p���N�Wg�V9�{iP�w�B2�"�0A�$�j(�ЬԱA�#�zY<�UZM�.Q�������C�A?~39ڙ�3�e.�#lB�C�i�a�>O`�x{|X	��#(�_	.����1V�5'A<	���˷�倕x�!H���`������&��{Mi�[}�Bm- /�!tK̙�Z���p�����dxnjJ��B�@�%�EB�/���H�d-b7��,k��0^��%��&v�G����s<x�^s�D˧	�鈗���Ք�
wrZW�Y�]�l5��h�F%��[�Im���ˌ�dP�&G֡A�s! ��I�o�t�z�*���h�{A�:3�⼭�5��}a�%J<R��]6ơ��?G�L����R�R��/"A�=�cd����d�.�k��,u`�
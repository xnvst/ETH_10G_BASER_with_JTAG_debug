// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
SMGMHrK3h+1O2nuilQWwjiFrxwflZWvH7oQr9HuvmV8tUYUbpXXiVHiVHm2MfNDpM08ounNDsT58
1YuhdpO44au/m0+paTOLUktzV1NqnaPO7kkLlUlhkdFlamdU8aeF7YfPm8FeQRXXY48pJXgKUnGN
rHrkJYuGIMRljYwrCvmYNoPHwgcj1lFc/rkKA+wNw09mbjcP7Ruq8wwg2iX/YoHiDccXNj/FW0AN
tkUco+UPMuKrDEgBq1ulCwT9CLFz5qYPm53xC6mcJZnwIa5E3mtq7sQIAxaLoK33IB083qy72KEp
0GFHR6UGOkc5YJW6CJEzxeopEAxtjko2Phg7iQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
jkOSJZlGumOaQ3MswoA9ETAd3qNI/RbNBiQoLHco0y/YVR36lTe/c2drJIFwn0yQPSkmbvJLxcuK
AImHh7tD0ViKatTEvOrtnam/fN1UsKHafTX5cS0Wkvb9vzSMpPCwtXWEZRpTTXZNBn3KbrvOS2sz
hI+qflS2WX1k5BpRj5LhC3RkWCSwhWqnUD2SMOWA4sOt1EZOAawJ4U5PWDxef1+L+uCIevO3/ggD
bhBU264Vqo4WrRO1HYsHETpv3Mloq+ejJzTgqKMoqCo/BvKWP179kLnVkrKkwVJ1G4qP1EywIw8R
CClfc6bscmUqH2H4Pe3KWLHHhCOAD2VP258ztEhIQnnnP2k6cWwK8UohKcND+F8mjHkL7bpMUeFo
F+AtMcGSSowuKOjR2CjDOozrVd5GXU1lXaWd8w+2oIiSEJsZLh97/34w62bLbAE2oVXgpSEFqNO6
8NTFdJW9s4YTgUC/DM7/vXn39FPooaX50wK74IzksKFIg2BB7slB60mWSVL5UqLa2rvFkKYjArzG
CXgEjNN9y/BIqATsQnEK4tO+ef59vk/dM05mQQTEy0caYeqh3WCpBDuACm3mx3SAzOzXXOhPrkAX
uQ0Nl+o7it4PSI8IELaDdS4AzZWRyRk9Wi3VRzR4hNU+0zefRoCyp8+9Vw2WQmaFdXHaAx912nFX
0m55TeS0a6PpE6IKaWXV346762atUr8z2DG4fBW1XNSN51Oen5Ildte4r/A+8y5YSZN4ASN4Y+gn
qY6yH/kWBUtTHC50RN6H83hOg3zt8KCDRyMzw4lqf13AKt07UNuu7QVV3X0Wco8oXZTQWRws+raJ
F2vpHh5nmfuQ+ZXOzPiaMOCWLSmUDu1bgBolU/3jFH9D8NAAEUkFc4HwwmbB9U9Nl34PUL5aJRHb
Sc/NdYupGWkbmq54MsjK8MTyrVIQdiKZ+2lVMv1g41oA7GW3/2uOw7thugGnvg0CX7eUmu6cQqM9
tCVJsC3vRTiN8LfOg+DhSb6IJG1Nttvvdo66mpsT2Wai/FZpwewwOV5i0tsvcIzqUNxYdcwMx/M/
0pUaQOko44orAnZDyGDskTlXaH+Tc5r0NkOXF3Q+0sAZTjK8cyEKeGD6x/6HTR8zv6XtaByvp2qb
lznMpag2erVvkGmk6uKxPTLB7wfueBs2b2HffLuk9pfbBhIDvxyDD9eXyOdyTd6MDmb/avTLcEi2
rUuoKXrpUtXTU5DOUFLYkHwuQ92KkeMPZ6whlzmkYnyNxZvhtkAHQrKgln3RIT7gw21dn7q2LGej
6EbMdzMmhZGIFXEqRNbZ1tWHdEi+WjR6+ZP5P0aG90uxV5KoQVbZeVMtz3qyyDOuV6+sdNkGs+K+
af2JW7zJ+z854whRtx0rxIQyBdQBehV3jv8unZA1sziU5LGMv+4wEWcA62YwgwDzoDYmFQbdzitx
nLJl7fYJGSuWaiGMi3fZXaI8P8L6zEi3d0bFWYQhsk4yrTW38H6APnRq+cyMS6tJK/foNBChy+/L
XnkGt7otX1MOaltHEmHT0um+uLV8u1H12ZzVFAIcbOSPtEkwHsmRNxdXrGQNgaNVU6lwrR5ImqJP
ZkDmZr2mq85MDowbw1gBcOwjh780sqJdUitR9ouExa/vuFfumWQY6vlFNRP6VyYA68zeOZSEbjKJ
GBWQP9IvE2dUlHPQU83/W+dGe4MmLvmBHmxbIf+T2n5cpaAu2GGapYET7ajARVZ1q+6M9QLkTX0c
DhhkwuusWQBvT/LsXLFffwjVpwZhbeMLy/Y/UVcsmaypUr7NNzM1P208d+gwSDx5m/is4gKAgQND
mB0GtsDe5cvac8AR2vxc7ozd1EnGQTPD21HuheITmQSK1baFQ4+3h20+JCmuwmHr8p6CUEVw8N5Y
6I+p3RnnAycfsJCOjgKGqYAYEQXUZr7C8aPC2joqeTPvzxpq8qregvO2ifzwIFVCf0TDXMuuIhdj
9Ptpf8wQDjT894uf5SXqQY1Ac/wh6nC+TF3Lp1kBRGavWqc0b/PEaOXMF09rFVD5tzCunhbjnuw5
75Tp5ve987DDS/E8nv0/IJi5Zx6dHzCpfEhvsKACH+J2Kdv1U/0uNSgEZRCbSzRrytuxp/+pn2fs
LpYOeJQWyvxHalW0fSCgHWHUXuTy0uk6YDhTIZIkJmP570KrHfSZMj9g+xgsTdz5OFIdAkmG73JX
4kGb73N+uFQzBVdNeeG6xo/v6Sg5RS0cBvGYwW1o0ZZRFwDdClkRwATX1W26d3z9c0UTXvtr1rci
qBRIGccibnqd/9csMBNW5fBJ/ZcNAKgof6EPITEkIYXRjCWtqYl5pZvv0Adg12ScupFHGn6HUZiX
wCsxxCKgdvpXp7Fniv1174KfuT62od6LRq8WQ6Ifln5p3qHWJQTP7kKsQQ+gE1Mf0ape7eZyXWYT
YavWJ8JM8Q1rATks0zFV0kl4CbgEJGBmU92Y/0MbmInUUxyLYq5Kmv2Jc5TnwW7wiUxBFH+W105c
Oz8JYZVQubWT9jREa0Mcqgn9s9XgYQ4A9Zap1TefL21Kc2ckmmfXCv5tiBodrCmSnggS7XkLQy5z
huAVBocn4/YFGnC8tmaLN3L20yD6f3k/E8CXFi3hqVBETW/cHBgQYp3RxIPBDVSHh4TsBvEu+EQK
dLXUADbWr4wNCgdMEVyWuwktET0+YO10zBFcjVQkTdL2X1BdhdqYFmW6zNASDHcgdqWsYykEIoF8
ppdh9JHD8o1GmvABsfg7JlJ+odio53hyqyh6GTcx4KWHYCaiJJjTLkisXX68jwKbj5swsxPi4Top
Z2FkFVm6V07FCt8qLml3/qU8j1vkDL9BOeAhsud3Sj0f3QF2dk+4uAvnDWQT179Y9V9OTOFbOl73
wf+jwRfhHDM1zkqiBKvcK5mnwN+NnJ5PDd6oeiFUvdpcUE6wKXXm0ETz8aOdMd0fIK5ymAm88JTb
LtNovAih6FALQ+ECOhTNpzRrlEe7AD28fV+HqN0AF+2NCxVWrpNPwnpr7UF+SAUH6BrEZKq87gtJ
LaX9bc/k6v4oRJpHxowWKIJw3BcJJUNzmK8xmM725b3FwqTA0quXLXNpjvkqmxd1x70+Bt4F56p0
e93IFzl0aqFZ6DQZNvAifba3wvjibLMeU6bDHKwk9NB2R7m9ZwBUgCIIX+kUGYCID1RgK4Gsd6/+
fxHj4aolrJPzaZP5tCA/G6H5zzdM7T0Di/4KSb6kqBckCtqAwq23JJRCIcFS/w9vtVleuyvsvGYv
msNG9rVBkidB+8AmBa3pS4Q7cTb2+u1HKi+971ATxa4GZZ71QzB8QTEErAgsn9rXBv41T4PUSNyw
LhaiejxIz5LYfwFmmrJtXUU3vPbZSSYODXbdU+Zrw0EWOnlJlKsrDHx12Cc7b+aTOAkZ1HPBIw5g
dvZA3e0VUE5V99g/09GzuWAEGE/zfjTsfMZvzXsiUahgxJjxxCEOisd2Q4RdZYDK+0HqkuIL+g8J
XhWSDoqhYoumx6xV9WqkW54Ltcnpj9Q/F+OLBBeZplGABTQbZjDSRBcOdjSX7WR/9o+rZL/QOAgw
+i7G9n7t1gTE9HJtP9yKh/kCZsL1Ce5VzZZd1qL+Or9PIzj+XRhbnRAcGhBBoKDuPUyRcphgx8eu
ql2MchuRKaOmQo+Rf5u7DXNHhrpXJvRIWp4kmbYlMZuS+JWC15EPkWppOB9Zg2K917d/dPeYdlBB
g0xSB8qADoJpZnR0y5eljbynUuXZBiW14C7GkU7ygqGG25Bvs7X7Z2feAz9Fkv7ziKjqr4WnQnvl
NbcUd11ucaw2uyd7Em39OAkZAr+5D2YKIyYJyJkg1EKZ9scTmzafZWZvIdn1QksHxbwkeFHrTgYX
9Wh7DVtzrh0EAsmwD4k6LoQrpMX20tO2YviX3QhFzAmw8Zxv7ed3koryoArNqyDneBwVXAWKlf92
U5Fi8BERkotc0lcp1/UhsZ2LQqYmpeFHnOTUCyUJwWb9yXb5hV63hbR6N38H7BYjCG7vLWfHDekO
wqIQDAD1nMq+QtFsm1T0lC+Ohp5K4K0CXP2NGW73TEAgNKb742F4TEE5E3dYn90zxNaKwfm51hNv
i14IYpXKQbATlMDOkklrPY14dIWAovAZVeCY7dJysSE0qfUo7vEUAxdVcmHHZuTxSXxy8iWztBU1
RmIDUCSF05GW8ZtpnjJYxjKV8T3kWvSwOlC85FTXM8FAuWrWxm0XtCU5oTn8yjpaOyJrTdxK8mTi
69Of5da56VmGcWN44xsu/J8Xw/7PkMqNYT4xpgQkPfJSrHeHUcq4qZcUmOpZJ70DtrzQkM9xcjD8
r0APtWcWDFz1vg2kMbryslXbTeXXLdgXh8CIB+e0S7CNN9zBStORJMVRApRFuv23r17dY3UWImZn
JkI7dOPbmPWkWzvmwlEEBOAV4eD7J8XtxnzdLYUZNnXQVXIJwHxUWE55v8V3Zr2CoIGwZeHwwQtX
J4DsEcfGnjzcIC4yrFCg1aQu6IJgAw8BQLP8RejkoX2gi29Tuytn33IQB3U5Y9QWZo9jY3Kc4oAz
Wlo4k9BsdnBZ20sft5VhCirl7vS3zENg+ajj1DpcwXrPN85jzEWSVdAAqT6nG7WoFn2YIml8k5mg
QftuY1yuxdYud/E5+z/+l+ZgN1QUFmO24mNDu5yu4JvJ96tO4ePffUG7a356Qg8qdpbinUXB4eKZ
FJGEuv1dKlb6Jk4kU/vwQhAJdw8X6vg114Rs8ag5O8Xeuxs8nGqA9DR8VRxE6uHZLcAkoykLZqQG
gaL0S/CZPTwkuYmAkzw8I5GRqI71ZDKfeu8iLIQBQQ6XaCTEG/FfsxJsBTm0n+zYrwh80oQnKktg
8mH6Fzc3RB5wNIO5EA8BxTR8bNiSv/n2Zins8/egHfPvz0oSbijhtQgyzjcL7x8nSctuYMfPeql5
lNzqnXdg82KcI/VMRXDcDWv2M9nZ78fpsU31H6KWspvJDKWK0M7LupEvAniBAcCVzkBeCnjVemqW
KUrAc7Y1dkUTAlmOulB8BQbdILAN+X2+Si0GCmJRdwn6kG7AH+53yzozR7pu7bRgKbBvh7iBFBLW
KCq9cdOisSLVLhuR+yqVCK++s7ve41w4ovI8E9b4gJAtfj1HIAsyai/YSjBgpd+1NYXPISKa8eXe
8n5FxtzJcP+B8Pb1UwZegGCKD97UmpMehEDyiLUEdj/BIgNa+GL/wGETIDV/Ue8FBjgPzC9dhG3w
VyvNsE6FVLYV3FqOC38Y8hEI3Dojvh7mZJ+nZXohCRxuUM0dFYUDL4GWs/US+ztiT8tfnk6uSmhF
G8UsJ9mrz6jf9VdFPuLX/oTfwKrDhVu06IaHU2LFiY9bKu0KW+WcpJXCE6eUSciZuoFJpHHMqHvm
f71lNXDzzCzMGF1nOKLH/Jv09BK2Np+INn0QXqCbiFo61FxSgONPjDQ9QvWfAPWRAs8BANVIKe+b
ZzHWoe77+5tyypBv0nPYDbwI9iMqjKf8/30u5hBg+YcNrue771+TOJ4M1jNQ49sSPA5dK3g2RUfG
BVt/BylV3lKjXPd3sJS8KHlMuM9jSPi5ysFndHhpY9/QZuVj9M4egWrQ1l/2Ay4VNQKnZgHfnjqp
TyAiND7pLCHOIWdliM/hTyK2ReM6O0Ouu1h2EtnV8q8XAVXG4UxByKr+lu2fQiObKGmtXd+RHmJK
BvJz8AJ9ezUbA+0zXEeq/vikhSGw8nTs2Ty6o+51WQiBf7JXfxKy7tPB8pfmLEzjpLOpHguZWHGe
brOPW0zvBM5ZsdsqLjdqUNsahbuFWPxOVDKEYXaLwTvQCQIA5rFXHn50hPv1Mv1q64WoBq6XOXzK
ByvACYW/Pfr7TdcL0Wi0gp1yMUAF91W31PNacWvf39JQUpniRt4ltJ+w9sppl1ecNmoQIv0s4LNA
QJ6rgSbe5nm5ALtefQm1LzFmw3+T5lkyQdNLkmoT7lSxrg==
`pragma protect end_protected

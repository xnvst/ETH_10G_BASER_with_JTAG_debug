// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:30 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IqB3tS3rSeGJrPyGHQsyEBDWSwRyeNfLJ3h5xyRgj6/pki4tFDauy/tM+fsvsUp2
4lZWvsRxTdeBAsa7NLxYpNj3ZSzeyzOAzAhAb34yos2b7qkR23lzE689JbD14WVR
KxUhmr/xxnnQp6XaIY6W33WNxYhQXEMMWgiXnzkGlBE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28352)
A2tLCKaX4Q+CIIqORZn0gXYv4yLVmq6fZlglBw2CxB7TO1xOjCr0TBERWruOapfy
Bqyh6cXg3qK8Osdqq+B0SBP0+BylTncEQc/kDhd1fa74TkBbygOPfvn3FgRskeDM
4xEHpqftiWjrSX1iGkmQEndd9b3Cqk7muHSYVLwX2fjXaCKgE9rfnmhJcJJ/j0s1
bZDEShqvjAm1XnzG4HaXAgUEl1lROAs1Byis61rdm5WJHllFT3FqiUn+KcB+B2uO
3psfUbknKRmdqUMwXk5GwxFCpf6DnBzn01ZM+hYKTU1Pfauc57oIhewIdY8b7jzl
IZcF7yvFrN6vOf+xLbl8E5h6Yn2hLhOxkm8NZ8BLBHooOZKq0x0lZkTDgZr06YYu
3yj1jCPtOaUpCSm1ODbUH5fUEobiiIvWoktjtSrr3Y7YR7Usa2+w5BM88KLtvZdJ
xR4PTzNATPUjMD3VY+AYKjNxTj2/08Mwvr6XszBt30DmJ0HoQbiH6PvBdOvsxKKF
QJn0bm85LF/rZAZQnOWs4atYFbwyAMd2NPLkTUPuTUunHl1OJezaPwq0dRvPRdrH
RHvSkqyvXEd3RMVQpWLriTI2TvU4KzrOAGImwCOyS3SdW8q1iR/m6/9EtXGGghs+
h97fEl0hu0Jb3ovIIa5B3/eBBC66iqQ5+TyBYAyTr2SE9fhb96hmN36ygTUvK8jC
j38uXV1PSl4nlJgg36PwbnhT+dkvcN0BW7lVqlWsN1cdQPPkR3dugxx68NQQUN17
JrXULeex2+MlQBfYvMeBJLQfilTb1biLRagbSU1SWOuxDBSBpdn+VnZTBxS4OOkc
CuXmHUJE98JMEiEIfJBDhJIhlXXyRH+sxKV8uZcIDN7QIjkVYitN6dvW0eFMLCbS
BPZoG2J3W58IAdZK94Yeq9I7V8szynplZJV8wmHhnVm8eFRM8L/SZJDg04HVMPgc
BQUYAXyEef9BWm/d/upNyK/MEiUus9hWgcNAI+srav23Gc2TpTo/FhRHtmxDjkUk
pGaIU5cqtTJ0O2UXuowjgS0ViqypWZqKpZAOUKRNq7KrAKYmtdEXpgj0Lj8hcsmC
kqqaUyUaInIVU0/QoXXuato6AXy1z9x842o5GAg/MCS8Prmo1CcjXR56lRMm5I9Z
Ye40kXitCWt0tyJGLTafGyR6YltM2KXsHOy7j6LbUA5bsjWx42k4PbEeaWBkgic9
/ldrpm9Jr/3bGhmYVzlGHk9Tb4ny2plxBRxSS3HEn6knkOwDaIbZQLOZ2TYxP7sK
BRhWYnYAyh5qJDtbrgJROaDJq9ezeUrXSYxGcltVYtfxEAmyUL7wo7VlcNAfHV1q
vnsnBIKhM/VHKusDrSuduE3FhjDPr6bJgiW8aTreeS0tlenRmXfdcoYjkW4EB+/a
1nxXwoso94yAmGoQ8FrwKNE1IK7ZwgbfXVrt/D2jNPSFawUM93QtDmTM37r8dTfr
201T4ty3fzj/l8gZA7F5NnmvCkbKf+G26kwNhaICS18Rap57I9HGAHuMyQeNd8q/
f3/tW+BP7y6Vj9EX22kwvsx1qw3cadwVdUbtcQzUCcY7hLk0mHxIphw8t3jDE45c
cnu72EvTx1JOjM3kKWK1dh9LRIhbJqQwDiuqYVMBOgeLyRKVmirQpMWNUBvfz0bB
dLmSO/GjZpSepyWbQJMRRxNln4trfhebLuwQtPHTe6lxGGaOgQHdGfTOm0uh+YGr
/sjUdp/8Xf82XKdtaSKx4VoytR3Rh3/WMFvKI+0UV3olBbaKFeKRNAdbiv914Th2
v9YXKlXodmqIUOsPAq6kSRvdvV9uqapGEuRvOfaLHQ6Pj4NQ665CPdFqIKnYjAd/
nflviP4r1efSvo2PjJMkGICd4iMZes+ms5WscxNL7gQBZYgjL7OTW0b2vAXziPlY
g/hSWeVmg+PjW/X1ihBpKxCJAhRWx953R0NlxUBNkTMQqKy/p+2RA0fJtK9u0vG1
6PctZf2UG8osPohTdE8LBfmuibCBlEpZpRujXx+3DLs883qFutx1+72fHHTTCj0d
UbaF+nW09QT58+uRlvsu/H2H2wf+ZYegvHDUGrTt2Po2NdLh+KlrP/J5MqMCTKRE
X3Io59pJJqe75Pqwm/iWURvH5jNqtiD/b3m/6TScnBabKNMABxPLr3U+31SPdnj3
0YQPuArWMyRY9rxVJugdcXpvf2odsoWer1DR/6yhpK7T7VNuYN6EFff545yMbwig
izuFGuKpWp4DVaqGFKCUZ2EegoFRKqeYCWCNx4e+eL2N061oZnOXVVMC5DdOCGMT
jNCkZVMo6LjUBftWMWX3+IDw37STT2nJiZxNjUWR6OAcuASi1pd9576mWosGAFlk
YdH4jnNxkO5WoE9q4qzEatC+2NJNRin3foUl6AvhNpMspAGTJefdajtJaDXR0PFE
uCZ4R6Li/kpHYkaSxbxUEG2La40VO47DKFvvC2+F923Og5fYS3m0/gBsiAONnJiS
j2PWEvbJ9lRnpt4/8Vy/2RIrKI60gsaBacRoDQMFEIhphThm2nW3yK63jj+OvKz0
ZYA4jbV9Sgk8kXI6hOVMMy52wXp23UgSJgF6ansjNjCzkBCatmFn0sg2fU0VEi5e
UGMW6QNvzU94DjOM9p3Q6PifsDI0yzwn4aNlWts1EVzesg3zl+Murh40L1p7vozm
y6GE+fA4q/bsauErmoz08HBp6yQIL2fhVz4kd5T9OLWS0Qv5r11rfwkyMc3/P5js
AAyAX7p/fSXUgGOOKegKXdCVFir7SZhcyINpPMAJJSzUW3NKNIZK3CzWqHW+X75k
xuJh4dQOpBO37VVahZRS99EO0gdZgKWORphCNWkQIZAuIyf5kNJHYHB3up1SrTPE
MFZo7+uZGlV5GS2tMbaPQcSx828fg1Qan3YQOjlkBtple0YhWsLxbBT6cSofdF7/
KfcCdWhcwjz+Dk5t8NP0mKoetdM99WQVz4ARanSXTkG1gbSYzSkUjvaHkvl0pY7I
hBHNj4ZU0xQjjeA4vNkbffKt0A/kzT6uH7jFGZK9V951x9RpES9SssfALbUzkaJz
DRq4H6PDRavaD7B8kcRNsivsS8ias9IrG5OgvRI0gheVJXpaf/1j9+Zqndu7xd2W
ZLMDR5q/DtPVJaJF7+j7x9EuVfUKcO2p++3UvnlbqD7F/Q9RXb+TNpnOD/qT9oSv
r4GpJoEDwFjrl7VOi0ZwP6VZzprHqgRC0BovnOPmAi3LzCY+HrC4KrBeE2osCNeD
I/x4rFXDL0a3cdfPbnMxHq+M3/Tfo3oiRIwHAvAfCByU66P3WiGhKyKAmtfPmXtp
Sov8J76DTU1eAp4rqJDTRGWq3YOcbZ+VpiziLcMgG5HJDbNUhcrhv7sbWZedTxnL
m0bFEbgm+xx/v+rsvOg/EyDmFpyOxDJCF9Hc6EPnnIGwsiMgtyJVfcx2QSA/18Df
sM8DIrQkx214sgwDrTreBhstv2MGzDo43C5059NndCyUIfXiLCUiaV0XWsJpVHci
kliunR9OyxDloPNYo7ckzuErcb8n6Kyllwnn1vdhlUoii/u3MsMAHnvWwXoQsTor
TiCUVmp8JtQAEU0/WYYdkVgE6P0DIVQoJK0y6Z314V6zVO60ePfV+SjwwrOBQvl3
x3joGhl4n6COdRKp2t3iIJioBlc0KHFCY3vow+pARQtsB1lEtytRTaNTn/WzHxLR
Rsh5Jz5hSlc3ypAwTb6Y79CQLasewl/kVEjb51WdE2lb4qtiUSPbIGxZParCfo71
EvbSaq3CzZH1OhnfHWlonp0EgbQZvnDhb0nD6Wh6EyooIhd571+D388wCbfP5Sfq
xPt1hkaBMRNZrbWtNCU313xTFxt19xyuvOx0wPho4KatdPt7+rnEsEHmPcSqAyDw
sZ4Ik4jYIZf6hEV6XaOWgzD1LVGPoy7ilhQU46yisgetlYNp2wjVVsTgmE5WX8qo
YyeG+rZyCDD3pPz1SW3vOJcfTGxIhjx3QPz2VtJxLn7GlUlDPBCUv1eoHOfOXub+
GbmJHZd1RDuzO87W+P8Y0b3UzgE0JoWvFbRG6fQiOigwDwYFA03GyBJbJXRQYRXF
m+icTBDHEmgaVMIt6bcfmIL64ANu3Br2+ZfYujr4Ytz71HSjpvpEFzJRSkxUoTcL
lnLHOQ3yRdfJfInZdWn1Oydt6ZCKRKDwdGer2hof0e6LE+Noe2QJLtmKF74lbdlK
xO84xaesUsJrQEapE37j90DeFJTRYphYPyKdVXpli6++2w+CG+7bdvx5uLKaYqoD
LnTkS4uUjzp2n9OJU9e4Gw1rVjId9MZ8MXWpGsHxKc9ylpKqKVfSiIa9qc0CuKga
uLWHRz/81wOqJMYYB23EdTxpIG53XTDw9avnvJ0RlnVEKwJFbkVi3wjIaOtBXyil
hdi4DCATA0F/oGAfv20fhnwTC2HyVn0qDtO9Ug9bghhGE7vQF+/Ur31ren16dYiy
/rkkuc6BKYDUl5PCGLVI0uzc3Je4YXg1NMM1adqEp2gsGOz7D3G1527F61z4Q5Yn
Fpg/rqE1FhdjJkt7kFS/oXqJIbCV4/1bDmwfDEF0k88mPEIgBbz9pMfZOfc56zsN
HtZlyv4pjJYORQs8mJ+C05qEwt8lGKY4mNA84ZSJMZQe/MbfWVSyvNDKRZwZ8S41
a6CJgGrq5GDsNVxyPmlJds/iO5gVYej6U91oEtyjs7nomLXHDx1BmM4DxUUO1s/n
CJss7d0Uknv/fT0PCAX8WEofqenxq4NhgvhoD8SQsTbsZFKmKLMmsSpb1xRy8gZC
9GzC2p/DJAJ6vWa5z16jFlc+/oZw6lGygqLp54peiSViOnH8uujiUUPiLnPNc/Je
9VC2vs2IcKNMRHXpCpNHq/m8x5BQfcIcH7AIveOmK9gnYDHQ9geIoo4CHuTzHkTX
sJdJgLCYO/SHlEWa4PpNOJ9LkgIY9dxhYI3/eef1y/TpPGQazRbDrBmSkFjdWSS+
c7OmpdG7sjTofrtMuAPVSOoixAcXE7meGv5rSzThOlrH7lXynzbIhoIL0cLn+ffd
SZKPsfWbL5Jjr6dsThY5H05NrRZAhpvte45ghlQlC5GLc4eWTHTd7PWEDzItegCW
F4y1NLC6ek7sSpB/lis6VtoTiZuQQpuKJTn3rJ1g9473d6xVT5qQwYyqKp+z1bEq
KHCeNDcRi197qBJlBbY89Npd4P4ePCUo2LrP1k5bonMFa5FLczHLDKvbcnTNhbI5
L8bPg22aEMP7gjLyQ90RHlWvwoAsAip1nXkoRD/bmZw2n/CdCxPbsH5GIHvgIodk
CAJgFNDwY4GiwaNNiT/varY2Cb34f2vBPqlqWMBwABVL9L2uB1Y7YeiNhozd1Gtv
7uLn9w0iJ7tIQwRbHbNMZdgrIzOEx09C83f7QBGMd5d1fqbvXCBsK5DNhQ89NRnw
7uiHlllSjV93B9niBqVPYBRuVPnY7qduaprcya+ExwjYL7BciuCiV1EAuItlVi8C
vmJzoDZRd6/Svis4C4P5NOUJ/JQtfdmUhLzCLiUj1uEPnB2HUbfm5KqzpDeVODLJ
GJb+JPFCgYu9cVUxVn8VJ7JYvAbwkQfZGeRMBZkColTUzxDUbFOoHDxC5sSRCScX
CgtSromQl9qoGX6NfFNcV0oqp7WvzwxyqvvKZ5aTM44S2p55+SooX3ZlRJTqNg0v
2UnZUqpLSuLDrA+yQgyARwsrDEwAt7LJr8lZRduXowRZgBeV04JiK3xbt0MTsZLI
HaYl1kWXWGo5zPtLFtVJkjQ2fUiqQ5ka4P1I8Fd4DyFOUMBJC2J636IbkIMPxJRa
j3D5OYWpCvrYtRde2Vhh7bJ/q8yiqg4dnql4Px0eAVir5ipXDDfTgVTkhmmdgixe
yHlQNg9i5PcQSlhI95E1vv8+VlYmoAG7EDDsGrHfp3u3uwx0qJUsBcRF0CI7GcFi
G4L9kt2EyD0NVoZTJQq4EIrECF3klnf+a/ZlC4ZHJEoIz30wLzarlFJIuZgN8k7K
+UWVGOQyLVNxhKB6ZMCBFtqgs53mK4mR0GbQ17wD/UmqEPD0WuoWLlPk3zlVbP/l
EOqYMYf4Y4bZMDxJNHfTbQ9vtnd+AuEsd/NwqGcXkxAbj/U7ZsukvhfK9lZPm6Dk
BlwRxUUuiGQh4lbDd4Vmaxpmemh9Y1+E730tUi+TL/U+qZxm0OsD5fAZHn/YRqBL
nCxX4034mLf0SmGUOl1TVRmWs9jAssK3iBO7jPYZQyS1vOkkSzxnuGMmkBBy2aih
Kosdt4ijT6QzhyFhPajpJdsbrTlOCxMHGhZs/b/9rhR513bdlA/RCMRutbOYsr+k
qID1WLEhbwCNw7oxrd9k7rGG1orLdEhG7xhO54eBw7GepGc6UwXtqc970fd1bNO3
4FjI9BhDKCW+fGCEy/5RUvhD9/S7zxI464xvBxot40p231ToyOsjGmdHkeyE1n72
JUqznFiATT5FKQTMdtCsK7nKmj6yJlu5+B8WFD/spxwPuv73lz/csq7eGAg2lQ49
3asI/tzxygPlgxqJCIFOAEelMixOHpkFP9187ZOeF1GqVeOBAIfDc5QixgzW+d2U
czxK7v9Zg1E2/wjcsXWqABWvCy5nvRNQRchcUmd29WG7aUE46yDHb/oZjzo4OLxt
G2IKJ2HsEIuCalsEan/UqWV/sdd+w8xrylJL16HmNYIiWe72UbRYkg97SHZZABUi
eG4yxnRbzaz4uo3BKmIwiWZac1S2hHINwePERJVw2DTRxzJ2V7fZd9kxTWZpdM85
hoAv7mYM51a89x6f9koXTBuIkIUNseYCgUlEgZ61sfnXUrFZTRqkptaczWpV1Urk
QS8+qAMDSmVz2+7eGmZMyMJqNRPWuYI/cnsuVUpSu943/a2JRFLs++wyYuuDq22/
z88LxsGRhMCjU4fHNT5f2HK6kwWfIY3cZ3sBoPtZfx+aEEE+/vvHWYi8p5AltzrW
cPc/rVJr9AVsPc44Xc3VO3kmIHff2FOHgVFvFKZ9NL2+AJCBfurQLfAwhVZgrg3b
kFODqZh9+S7ILP4Mds0uEj3isLnmViHtTtLNDYrx4cF08Lx7VdfOQEElFwvcAEcD
38SAwLUtAn356ZJZnR/pBDzdgjXg3SxCaS5cuEl3RvBbHdiOBA2QJo+19Ryr3rG6
TO0AlqYigvNu/7U5zG3dMcNlA/VXfSHv26QSEnbenGGBCpOELVV6LnGDI3PeXZjV
VqruEXxg5kGIMkgBum5qYHNgT0shqjduO9UL6GY7gvkYmM2r8kmM7LP9yx7BYz5C
WJ8E7aF5WpeoPfmpaZE1o/YfNphCXY3ttBYz+R3p3n4NUbrCUv/pYiQT8jH99vH7
ZDz/vQRA302B81EMLEY3lmO2/97Jxh2teBb+jyezJEImJIp5jxI+pZyxE8vFXYYW
hvpx8j2aHwsjwjBW/mRyNn3sBP4a6EwnQbFINJmGqoUI8myio0ohBOW7iAj8q5Xp
9N5Le9yo0xbFVP6qpbkXL0RueZki7+dpm5fkZJBxqyZv7k1I/290xa0KMzaUW/ct
G6ISAcDBdNfXL4j17Gf4JkEJcaY0nOelkw/yLSTKbpC1rkdthjHxJ4PStqOR2Byl
DZe8R9cmusHiVWW9C80w9A8rJoTwO6QVdgon/3eBqr/p0k8IuspCBcBDTxOzINqe
gI8yTuofCu7Tl4PfLV9dK7L4vQPpuF47d4X4S26g7AgwY/48O94xKbkLgZrCVMVr
OKh70L9HHt288CQeEc7IDufuvuJErHqKoMrWOWXXihoe07vsz44HCHN1LVuBrNZT
AfSOxKCBW+5YXg5ITpeuZwkFODkcqK99SYsL5cpVLfJIKEczfa0cJWsnnG/io+7T
R5hhwap7H1hyteyrPFo0NR9ynLLPQvVXnIZx/lCMaJWm/gvzm9dw88NMJjK4qb1v
jlvxGR87evn0DvDMY7PqXtv8K3HX/3Zz1JQ+coe1jlI+MWtinBmtHt1LCud3T+1a
9JWYcUQkCHlNQ8dZbq1DmPzPqMx7vZePDjGa+TJ8s7WTf9d6EPHdspNRPqezuE8u
D0ddEJhAXR/I7FhPuqBEACc6tYD73eAzCAlFf+m3/u/03TfgqkOJjakM2KybGrJz
RM1cq3+Qbuor730b7QoHYZI+l6iOetftt5z4dK82GlKTUp4FhT2W+R+cAqin795s
DJBBwU/NrR04UgZGwz7nfMAxv3jLGxBY+YxQu89WGU34QkhosSxHsOVywwiBUfcy
RNRQUjjA3UvbKnS5VXFm4FgmkYYv+wyCV3AwaoiSuSiAu7khbvrGwbmnBcAt9X+t
1YShaUghnCB5/LyqX7V2moQuxJTZSyQTCoFT2GWBuZeGwS8RoFhgBdqASvvJ2CLU
hfVJddXOjn2NYp2rF/u26uLTZiQ8i0av9Lcys5aJtwQJTr5sFLVDhCMsNRAga57P
dL55APITzTIfiE1wEL1QZR53YUuQoHTaHc13A/tAGB93W2/490CLifyDq4KUBi88
c+feVzAcrP7h6ml1OZ/wR+I7pRe6glcqOlW8ZINVbqMnD6I6oseRJKUAgu0j10jU
A1oP9jPi/IdCsVVJgQ6vJtqQ1Q8rmMQAQ5gVB9SCBnxxy3tzn7E7xXe4bGpA+xZ8
KM/MoXZocuA3NBjfRawyFaGJUYTdUCv580ujArKjGz/Pl843FJbWg992kuI+YE+d
BELAYWlGS1GpRVBbEl2baAVVobyRs1tC/akkZcwh8O5Pwd39LsgO4aprxu1A9oIj
FjkhnVciwzkmFefXcFy2o06jI+9PbbPyvg896zBQ5O2zDHMambACSZi4gBCGx2Q2
M9O5x3wEmvg2yf7WWuhxDR8zDN5IYKYuUPYKtvbYlhcaP0n84eIBe0/jKlUTBRSg
xGz3G2zLhb7092VLHoaG6RLRdloUqNwgfC26gtHrL3Lv0/p0EWKv9ZIZV9an6iTK
2w6wfzzYrLbeP4GDMxNJStBkYyiZPhwNjq8aC3eHMXQDsIoDyF9rZKf8AXPFGHIu
7nBhdNADwk3EUj4tbpDKHJ6GRM3sRQFBt8MQBvRtaIKmnKRn61B9vWWu64dif6AU
Y0HG3zcrf06hW9NzDSrveVgv9xxcTP52gEXqIPibBSIWUxaX5+izobxEWMKRj2Bs
8YlVlZl9bvF72MHx4RFyDJLdpTvqgED7jWXr40HNsQesMO0+d8+7Mzn2qDsa07ez
/vH05wDLr1LK3xsLhRPNjFYkWTopWmBKLxmv+u899D8JiucEU/ul3swGdELJcscE
7ZZExAIvnddvwyfD56sQ52YVMNijocSrO917i6jHeGfgSAOH1SXCMsxF1J5N78//
hyTPykpEiGywmUYqScnBrNpMb0YnepnXslsJOzACojQ2DzfC40ko5T4K/2PHkkf4
puz4iLuZXHKM/eZ7sbqzAq5mRmXR5PHpAHQ5yo7lj8ZpbMo63a1gI8OAVQ2bvm3F
8CfkA1oIKLF4uotdS53bmDMW+PJQWuBF4lZHVJWjTMKTmwJA3/3oh4fiOQLS3m4V
xzKWLlQgiqL6+TvI+88SYaiduFf9UBpi75flNI5G1/54ZmMOog6ugeM99P2gWY3T
8UFfXi69BDwY3R4bfb8RJoZJSOaFMbeduEEdbkRUZLkpA+f69GjWw/htqdvV6F0x
MHK1vq9BVOO+8kWcTZkTHebpXobDmp8JFJtmTJy7IVym+3JJBERjgCT0ykymg8mx
3q7y5HsQn400L/Zu1ucWvazovxtbkQ5oi2YDLS8xOL69rA5OvhDWWFmw7wtzf4wr
aTXqmDK/fARSFOcv/7IhTh75rkmyY6N4+S1a0iJa9wptBMFvq/IKg/RvE9jH+AFn
t6NnMhw+Zr67MMyXlQp7x7XVEmKTWbF5T2p7fNBtjBARZy9OnWtxOH9zLL5Mcgv5
co1EuyQ9QTm9WSJoGP5m/7goz9S1S4/y7KEBLoeN6YlcEFn1ls8NNBeC90GO3YLj
uXgBcR4bxMUSkAds/sgT9YYAfDRII90xmNsW2hYaejWFBoPPL+XiKa0pR7dILZ8q
bfEsFKvmKhrwof/Z1027OIHM5AQ8cto9BMQf1mp0KZrJ0HmcMkjzlkuD0QeciEaO
onXq1+RKvF7p7Rc3tOeuqZ9bcla3DkTZQ3S76+W6/XKsfeDV8nMXHIsP6IJz6IEv
0QTUXEVEyeum/9zzsdT+h7DMspV2gv23gZXv4T/uJWGefIHGeeSVicNueBuv+kzn
aFnxdWogU/ueDhG9C66zgL1p6IhrPF8sEtWC8JQQJASjhcpYtYOENqlJH521ltAo
aOtx9fMSdrCTgdeVwR9yhX05rGj4SK3ebHUUTPep6+GHU1QHttyCm2vRMmLRRYJv
8qqmrLIEseBHMtGphqG32zw/UQAiI0MMTndQ7RS6f7ERxN6DcTFtC3G+I2qttgH5
TUXnnYS9GqnxOpb5vcKYKVUWapDrtXdxUt76F0B66C4cwPpRaEt1CvKtJyF6XDnd
juuKU4C9Q7zeuL0wDt3Vbb4mJrJ7apoIn9neB2ZHkGDzrWypOvmdhVsk5zDIbTWd
MIiev7Waim+vsuMkYdo7zkYoZGfNH6LhpoNN7DjNblehJOF62qncAJfUXV0dVcFt
yDFFW7MjWWISkliOU291tfQ3H9Wf3bYLsKThPCevB1/j9vguzSuLyldCxMs19pd+
aAY7/Vu7rHopE8xnum/l8DUFNsyUgu2etDzV9/oFYhLd72qgVfzik8Aaszm18xhp
5WaBHjc2PHQ35OgXNeZyGKczGdOdu+U4oOFtPt7hFt/EFBTOR5XNbsCYpuudsAzp
ZtcDq9zaks/9o4XNTVUVDwO9CqErrybQ27PcqKiuBoSdOwB56CGVrjbH+PnOT35t
Zn3JYQS2BezERhbccdoT89gzty2FfQeYMcxoNYNkw4jvEC4oWawxV7EI9JTFaSEm
Of9gPVWi55/zVz10WljE6QQXXsnW2y97IvOc+l3GCGZMzAH2kCvttZT+VPQo732C
mHGi7P1vI8/4dDOLR2EtskW9MN0hifcjX8/Th2/1Bxoa09zCagQNTMVD7Ri1LBAo
LtL9A0q6HzshdOK0VgDjpdodmKa4uQdMtKcf9Zn2OHu5kSRx0ORQSqhiE9FKpbHu
FHkkeRQ0D8+iVESu1TYeySSy/X0pO9hlunvenYXVmePhi7Are6Dxj/ux4/spFKpN
ju/kDY7jjXkB0pja5Wt6tKGxHWwLvb5KaXFpF5VvUfCVQoV6IMEe+22SvJB+n1//
cfXPHkmoWU08Qtg3Xp1vcQgZaUBnn8us+eh/9RFD6rBQXD+d/wZ7QS2OT0oya3lS
WpXwtZDvkC508A7fIJUvrcbRb5T3Hk5Lbj0folX0QBDm8QQXtM5InSjHiRRHz7rn
32GLQ3G34F8PUJNMlIJeSzjC6nt8erv7CzoduMonXjg9EyuDb4kQg13M5BR+mVtd
68/6DIospbHEZVNEC1e059oz/vpeUvgFPkM/09X36jLLSu5TiJy7Pnz+s+ioAfWl
DmKtu7VCG8BIKMk7GI0QLgFqCgXALaLcUuTSX2L8tuvZPMutbajWUx1d+QbXlY/m
x/P3zigLsHlpLMx+/uNFvjBDpR8/Wlh7evEQ+A3CZpbGtIRM9JACbFb9UPTEP7lJ
vzbi2HRupZZn4ObsxDdu9gBzBLDSinwiI6nJnR0zuoCvIj4LwmljxqcT6IBV+xiZ
OS4Y/HFRfChu+5r40ly+D3QDY3KBTEEkF0JvHc36NwphjoxnT2ExfPYxS3OmWxwf
IZtVbvfbdkrDU+ZmtmlL+FBf23XIFD+MR4qh3Sm6ltxioCNMTZ6S1E3J+odBLlxu
rRRKIqj87+I2MLDpNO3w4PG1G6XQUn6ALuh1COytmbCdX6lqnYnAXCMvkvtViDVa
wGOta7+HoLld283yrhQd3KIH1U30PQWZpg7rXDaHEvuoFFzseFggFFl6xhaZcUlM
ybTgv7rl8Ql8WwbMPpqYThUGP+Fi+U9+9Wgj3BTFf6i7rOCHjtEmP65b2pam2Grs
/GwHjtZnj+ByO6ies3VQB+lO473f3TIjpMscZvS4bQSMXTLvSfcq73ErQ8QPTOlZ
KXztj7SbLriLuh5oCWdviylzJcwb/yxT7t6PusuZBP8Cv1VLl4qaIQY1zApR0WQq
jb7UMWnBJZ5xfEOnUPzZC7nx2mj6Ul3t3MxbGZICvVyEEtHrXfUVje9NajYPxLq1
MrY4fXjNB2eXIQOxRHloM1WkddwG0Emd2nBX5w/x7Bin+gOfNXfeWWa208ALSf8X
KabE+J7HfQAIxQe/IlQ4PrLuyzd1ouQ3uwpM+n2Bo14wJkFHzEYqGF++HaHKsRNL
myTxPdOEN4VGkTTf5yCu9yXPgFEgXueQrgbobvu/V/43WQk6jcYO9AS527Q4AerU
69SZTDh9SgJrtgmKRR73sChYqVgwuz9WPKbusQSHeBXAwbnBx9sdNDlDCa98Iuxk
efks3tL7sDhNYvs3owE3Tyl5CcGT8KewLdBdpbsn63KaOYxGfiRN+XulPbfu/156
367JltempG6XVOIL4dAsdU4vE2kO0kd9nX5FXbfNS7arn+d65Kw/bZ/N5RRAKbd0
KdoFpjFCPQIgXI3iKaVXB18DTnwkXxZuQd4YEmbUmjXW9vUz+08ZmOgZ0K2/ohYt
sCGKDsZrUVEwP4mj3CyS64wbhqem/xiYc7hzLXMKJKcGG6jy41/B9DJgGEey9wBn
oD+KUMBPKfTl8Y60ar+vUDCcNxy5tH7KAmzT2mbmuVWUxHvwGV6f6FhN9NZz7ZEf
hy0GhQtFWj/q4AvQyMFPeBZmqo9rdbEMFHZrhiOZ8oTp6vpn9o/obGfA4DIWAEh2
ZWBq9//z8+17u5xZMnHA6sW1hThkTPk0BkbGA8ApS78hTMkD9iBT5wNLp5HQO0tp
Hq6sr3A8rSqQHE/iI31LxiNtvY1TBhCvkCzJ79WP4lQnF/Bk1WwiJbWBTISwVPg7
HkPKZ8XKmW+nZyuaSTcOeHoRM04RgZQf2izzTL7yMhMx7JWFjiWI+QjplV1F+G5V
LvWAjs/GvL4Y8F6k8Rwl9MxlRqiGdH40LUWX/zZRqPofoonkGoixOPmWsmMdm0Uh
F67asQIJzDQ2SUSarVbSvbxk7YP04VBig4qd13ZcWH6BfN5X4IssK+in1VGZKPNK
augZEQyfzdTc7qonR6waqu0PC15ahTEQCeJN3WhKS0Ewju2fNCVxma5WwuqxDwVU
s9qj1ESMSt7TiZXTRZqOBXSOG1RRIex/j9tqqWOSqadIbQNXpQy27//vbeOWHfjx
s8LKFT5UO4bHOXZJF3sbyEMLlCJTIVvMFQZjgLNomcvCHO1TBN/mqSvjrO3uoDsY
51uRubpz+voZMeCn4ygvxgDiBs6CBVsEdtxnwslsBPPy7gw5aTxYUY9wyBfsT1oH
jLatYDCzZB5QGV7WM/6byB7cN+7Pj/hZ4UFnkNgP82SHuUwDtxnOCP+bs3wRdouP
NJaMgprBmaOxWNG0x4A/5BIptUq2Wjlc7MtOcewW+M9r2SnDiUj1lSqV3KHRHuqm
d7sBMTjM+y+/tNcTiomyB0iylCuTuri04Dnbb2jag5gIsslTOnZRBxTsJVlsunXv
OrP+9/0YqidPa+PGHvAytxFL2ckoeliMMUHtZVGanbymcnaQffvsLmGILs9Hs/ka
epYC0BXHbf0wrWvxUXROtN+hQ/hyZzQKK0lwD5/EsWfYhGJnYGzfjEAUVKVwsevj
Id4AGdYltkJ/odty3yCOgiWvyw5wz22H86uwzjju7b8medtzJmIsdK7Gr1CF7TBh
Ce7TNCFlkPocvF+MeyaEi1ivxrwH8biiU8iMTyNZLz+/tm2KIyS5EckqbFueM3Ps
/ugIgSkgz+xLJ/kTlZv2mccbvwNGV+M/i0pOg+wLEKVHzmt3KpJ2V2v/el9z3H2e
pvjD+Fc4e5/bLfCC4Mv2exe//eJIja8GHJeoiSJdgvhhdKSOmCZQa2uosgBkUPfC
AVUkzOj3+LiwfjSfXOtCi2mycvYPSiNt5RoUyMy2oOWzJHsXylatQSY6uSRRQ1gX
1yuKCkCDB8zX7YhWQLNOtuUzo2dseGWSw/mw4vRe116ZkE+tjUOQG4FL4LTSSQT0
hVlSTnmFifI0gd7+j3FEkrKvk1Q9BNaWqZzj1dNGhLgQNcUyNyWWZ21ztl9rbTVs
Jmh+yrzoGQ+ipvQ0vOJwfSZiylNfw0GF7Fq1WOonaT2bgka65CxIpBmDEL9osgvr
Q8GGd34dQD9PC2zVB5L+lhXSitU5ICPj4XwS8h2t6TVg9KSnwb8ykBuHCOJ9paRZ
Nc6wGfi9EDnfVbvppI+2185HlnZaJx88YmxAORXFPufAVfD3awANvDTzGxAFUbz9
XXr3fQVjolJnNdJsyeDBZKkywko81ElVAGbOKTdUux48F/5tdQvNKmbYMObSy9c3
W76Adk5uPP2H8sE26xBkw8X+CWjtOfGIHvLvgIyZ57V628Ulnz0QrBg0YKlFs6dh
Pt0B2P4/cO3tOk90QSeQZ76CEL9rzmFpUI8Xi6McoMKHtQRwB+OnWpz5C90wwnL0
KoCGithWjNnpPxG4mLOGNI0HhEjVRofuqzTKh14tixVoOjCLgWNuecljocWM7XuN
QNVeMLmdy7UHIiivfI/9pjLIhxJ/6nwuY2bS5vjT40YuufsPt/lPWNUKafq4W62m
BE7BqeyHBa6SqH4skGFIJb1va718veguRkJDHl7Gbm+cRaZrH2Tx6IoUvrBlhcTg
8byTfquYF+lJqBtNq9fxJM84yYOKK7orLR9Ah4nuoUdhKRS/ckWplrh9GUAwF4ss
j7OeV/WcqHh2rcS2zYksHlCdvJcDG8pplgdbAJhtKIyXRNsQFPwCJXlezgO/DLVR
1+xhU3Yv/uiLT/LHikACcW/oZ7IRKffRGabHaiUSyWu74loYkCCk+icMajzqOktI
rvtpTenSORtiTbZGbZ4doRHEWSMBfDzayPT1r2Md+aDruxcSMcYjGFMnpCtIXiTn
EhWGSyAdPrjMEv8XgybP+NjVCTisz71B4gF6N5G1XPuPGnajA0r5S9EdneU3fdNa
zBQcX5s0eiiLyZ4j9hoWZmY7mbmdr4+PoEhRBMcETS1OeylfVmGNr0c/yqDL59Sh
/NgnBAGXjxHCzxWs0wsFh036FTVTNihSNwlE1seGXToSI468TDC+LSC85kpJiaDA
tMK322CgHDQw/BQ7lY1GW9JGH+BXz73dUyKNf7flp38GWx6nzId4lPsB8hSaLXGI
fxQS+q5WleQbjhKUZzPwMAtioYB8UEu2XD8/cYgDophMa9I1UL78SUg9e9zCaiW4
Mprsiwu16hmxmU/RvXxYJXJ7qx69//EkC94TUtL8jUwabopjF++k2xbOxePyeUeb
y+6Y93fZoe03krAZwwqw3W4TrHA+ynLDjNBlESuBGnDujJtC4mJpW/LRHG+C+6F7
q615sUzVtMppfqbnCZc/F6olPMJAccVgJFjULVI8Ew/kH5GlRpKXaSH9qMID9dtV
oOwfrf9Jv+08yJB2X+Jt08ntpPNQxAnHawM/DvShnRMg6ej4l/d5y76uWYWpZndy
JMV9b1s1LuTmvudhPmLmg8+n+ZzBm072Zmg45LPe8/YIpgwnPLSs0lyTo4xeZUQ0
3Xp7VZArRWnTvvXkfgWXikY014ij2LTd3Qs+Myib5r3rFvni2z57+oMNcZd8PowQ
Q/wAUAg52Ug4FZK6idSF9y2yO9oUGo0Xf8X7XsMIgZlkm0YHIWXzXz3j/+/8qDFI
NfyXqwm9JOIBQGjXZcxiyIq38hSZGlkw72A1Mui7FtbjjuxCuarM+i08oM8lwXRE
rIo+N/sadpwcnWtgt89YxLmfVSrZuKzCF1UAyBykbdZeh32K77mbo9vVKniUq0l3
kdb1BxTs5/0OvZ2Ul7yyyChl5Ze6xnEUl3vp0zHr/vLRtFeWD33Pvg3u/GSpXjAR
m9SvvLf+N1D/iI7MwN9jnTYN931qPfzLUIQeo+f6CUMY0YiYpce4NVbG0tP+djQz
VJLC58M8Wa+lEJjT5wVZX+DUpQTYwQwagniukuIECOvIOJjQ7Y6oRqcooPM1MtLX
8h6eKWRttqXsIptouZ9ASuvzel6Oz5Kd41pP5RS9O/zTEhx5K8vRu6CLARURLyV5
q1yPUrsHwbJ5l6y0a7UiSpu43oO8VM7sudL6Z7wpoDnu3twbOcYktWAB5ULgIJcL
+Gp5NMcTAQpdMFPoBa3K7EshXCgiY5h7V9B2/U321lhuoYwXnfdpC7w7tzmk/P8S
9XcdoJbVnM4FkrKHaaa/75/FH1VYhnju9IznI7PQWv7H1QSt9zzquDWOgJ87GZLi
EZ/UYpsxr+LdsXZcE+RwuAlbzfE7FURoYTfC1KKZ8Hn0LjSXjDlsWeyfEfmEOUNH
xWz3GtvVxDkPSetpGw9qXktfp1vAiOtHn15Uciddja4NRfRB2DVxuxCSIsEo0Hol
YZjWp1m60n0GvYAvNdbB5HqyK5Bqs+PJix16n7+jTjvlu2i5uWWkTAwr6h0h2yYm
psp2Yil9esr2giwvSVqKORVFuc4VXSJtnUTilDAceSl7uod85BSCOVy2kF9RUwkg
8eCqz7b+yzoL5O6K0dMUR/feTrxUVkNXjYEySGZxN6kmQIcTYRtU5ZOzBkE14vX7
mtUUseHTSD5gWK5gIcwPNIzWbHjRkN07dp+bOK3n0I8LQDU0Up6O29ldm1YHeHhd
s4G76A7RlYafKGQV/Wgzsnl7ibSfs3RxTocQFJnwc1r+u0Yi4vwpW5vxhTWwQR8A
haXnv4QdF5UyANSvvLTjH5h0rxPIsVTkv6ba00wyWnKpXZ7jXvYkwsVR8UwJLMJ/
pFHeV3hNCOMJPauGNNUvTDDo/EgCe334qNp/rKT+aMVju7VOQ1MltW1ScYuQAV57
X31nW6j3kzXJr/+kcDXqCmaWcVdNnQXU9RcF6TcGCzVWqyL9jHFCI59bUuLTgq3K
vtJerhdBw6uaHGnn4w/sxCIWPZWpmBn5fUw+GCH7yjYmwb7zMR4VtrCdEMS3uqh9
YtSIyyK0aDxjmu1naxVIwJB/bgx9FD+X22qHhgfKEzUQpScmWdZTza9U/QmRwi1z
Sq27W/aFlr+kNzCLtJUYhcAviV+B+gjQGVoZZlSz41tb6MjC9w3D4E4VCZVlUzKw
B0GH0yeRujJuJyGXN+emoGcAbPVLEhQFUCR+2orizYIM+ChWPoc55axXYHSPyni1
JTZj1HD2SOrPbKPosV8tMFNDVdkIppBziLh+fhsVWmKoKdYxQRWdoPaTMznBuiVe
/KOdLKy9hlrpmchPvngthbACuIV+uT1IVwYKnxsd2Fh1/Ge7SIQOl2WEpXL5BYOA
eTBU32IRgAjerpvQf0V/H7/SB0ABypWLqakB0mgO8n4Lo3Mevh9zgQDUcXZNy+Mv
tkL+LBlmNdrZ/7f7mAB/GaOj8khMfELFtmCHzkjRHijCnRBf3+2IuYdcJsv2vaUy
GGQ6g8SMONEMLoM1yyRjlL4eXWeiEqA8FbMiWKXq/AwAmI/L0Po80fOyNLlsEkiP
tjVjr+32I2JhrQm6Iy1c+BKTxhPcLxVYLDkuEjCDYoRzzNoNfvZ1CW7roZNuud9u
Lb+WAXTAMadUKUq/4BfPzmHAmnHei1N7Ie5NZPp3mnXYuflREIsWWd4wenqD/jQ9
p+n4X038k8qWdepSzTRNdNNmlFec8MEsp/KAUY7IqI4xFej9M7r1saYR9sceN5Oa
9JX23+w773bxE2Wtya+KuLRyafBcOmuflioAB+cg/v93dK2LfDXY7BR1ChDR7VXH
fzeSfRHUfpaOjsCAdaeNxdpDxkluPnn2KOXDy+CmI+x3/vlnT1Ci0Utb/TkWM1X2
Xg5zVUl3Fsd+VwOG0sobjevm0thGSTWe/GVCW+zxz/yPITECwU6bpBp14Jz1CtOt
8Rb5jErdVIYkaIccAZ7fsXUxufC+oAK4+pvLNlhrE2e0INPuRiohugfpD84WbC0i
WFqT8L8DG2unVe91EltR3bcilf6YICuetuK7lMjXeE65CiD8n+NSo1DrXS6bPo19
3Q10wFS8NlzuNkp3iewlS3ByEgogn2mi1Lfqf/UpRZFyALKRKheWHCPnCPWsXvDP
CN6vZ/sTdZ0CjlM73oNka2w4JRKnMrxDzFwM6k1kUPU227voBvhbdyNbpceh1afc
WJ4gNwxznSBAMz+y6wfAh1M1SKUyvmAXpzhvETmF4ZdbamWPMUG3sDzAb9eCjLKh
h2AUtyjxxBNaUba48QwRXjWCDsAlakxXY5WIlO1X1xdp6/1TcgmVLjXkVl9vBu2K
S5QkWZXs8QMSVgn6PuzuIma5L8dLOooIrly2Wwqw0Ox+TIK0kKSvNln1edtveZ2/
17NZ0ZSnYUsQf1vrS7FOlpatAgsVMFoyW2fBefzaV9ZJgHEr37p+Cbx4JGT52GqF
KExfzz4m3sU4Yfq7PGuTduVBJSDfR9YDTZHLiSgJ50Zg/L3PhlMYijNs3humyeoh
VPwIrMsrhBu8/tBf/u+r/I9Heyqemrur0OgVAtP5KpM0f2w9QgGOdRM+YlYQChKP
nhrejNgLupx+Xxxxh9ZbDhiF6WWiqaxDrgJl23OKKt+UPSWMyvdKMToq74lFQ2Zw
qC1uGvFoeh0Q+hBovoI9iV4VhoUdXWMOWXcI2Xf75UhecrK1CIJxC3dvjiN05Y5M
quVy12KrYTiPbMr2/e82pSIXX7PN7B8+L/MVPwT8LxgOih6fwq3+F9oqOKBCrDhS
DEcO7FOnDTO//t8ltPrTTCiW/GpUTJa2YaKGVScgb2whG7k6kqPWVL4Qkmy5zaf6
p94TjXT5HazbM8d0royQ5X/+FIQjyrdfsgPgyw+57E8RbSzNprB4CApMtn65VXYi
teUb/VmfYPEo75mvl7198dKh7k0SzD2Dfi1IpB6Z0ngyqzwrTT/cNS/EClipm+Xr
8bku8G5BZqRk2PvD/mtEJ/Q/FSFs3IXVWm5vNO2l8te8WpKSQCXznmXTmJLr2xo7
+SnOU49D5rLAeBKL2V5hCOJBoW3dO1OLvbFAK2tvYHzxcRZiAb9VtPUPm3g+cqwF
ZrXBuZ2cY/CPNUCGhQM5Rjw8Dt3EkK+I6PTk0IvU0StER83NsOB0bq0lVUraRR1Q
zstax6rjUa27J3Cr4nK1RhsbUVsgJ/8SVm3gD9YybDYiRFYGqRAIOtS2lZM5BH7H
uq//Dy4eBhf+Y1I79bswbKF96OjKVO/Bo4Tdm1pJ1KubdEifWg/0Ejj4gr1r8o4i
Zv52VqDoLttM8KiN7nEdc3QBdrGq50G42GMtYMGIUPOMeR0+JvL6klXvS+HXmC/p
2GNPUlRrOcN//m3V4uXxTmGId7p0+Ax61QAcdS8EyD+UQdHbIALmFQqOy1heqZXI
2N0kvwjONdd813GTXJ+x2u26khlR/QLbX6xDlPak+8xYE9mZdxKYHo6KixQTEXEt
P2UXZxWWzpPV53f9e7ZA4ecQok22pMP8c8PWGR8QvyWRqhdN9yoMzCTdv3kTQXG4
r2BYp5ZJ2eswiclm3coj0+zKDRvjP0NwT18iO12wnnE5gGhPOiwMMAJfUdD7GEx3
FYvufY/Kp/DYVkcS1ANrdBGdQtL1vSHMCEKNlgj1IewkcPn2GVMgpvGXwVm8nisu
ZxFxotncu61+hI+4T7cNGOC7jnVMirahDBTtTCksoM/36b2lYGzwnwGBdU6piKBh
Uus/i6kmfJk+s/glXstoj5DqPdhHukDP7aPvPUuyrG3pO0gOmqHNBMXm4L/USPbR
OrQIvwPNlfbzMxwhc8tXlF7DkJP8OF5g13s0jYDncfsCSen6pL8aGP0E9OHFKKhf
LCjjA/7LrcQbbeKoifCQNIRASshGSF39K6fPLEEwSbieliuNs6sFs4zqM7Dtpii5
xOpDkM4tP7lBN6dCOUmW12r7BS+wuFFt1G4e+pN6ttew0BOJJ82p7qEL7rYoHhQ/
B6ljsmmhLfqSm/dsVe6PsbT19bUqAeXiccM7L10ElSKK4n2fEJQnLj2q9UM1d+nq
9vyejv8wTWCSv1Oa6rVuhdVoJoLgyx9fybwu6D5LxdECvPfK/HZIuyKraSNCL2D5
wXDFWllrc+scSFcVQHONRbFqJsAX53vu1ZdduRMllGAL+napPCogTseOlgmeLnfN
L11iSh7qNenaA2eLLFZ04+SYkfNOKrqMUsr132v3Q2EYgJ7/YoGiJl4oz/RM8oOV
oD3fcc25J9T/kbHCWAxVSAuUXKuemAVv2MhcBGXaS8fnZQY2toT9IBP88RhIVRFX
B/C27O5TdbadYbH2dng69TeG7Rup7FQlOhJOfHH0+TtiE91bzQOU347BcusUJfq1
EPRQ3Gt94iDjXm5V0IVfTJ3u36aHI73DlIxpDvrkXPKP/GjbqXWDLR9o1JyJLLOs
pHuBV1NmFWiDD19ahT6gHKQIegrI+xOYHi1weU+rIat5A0v/qZnIu1W7/jvf01IK
Rw5kY/W4tbx6PwWl8O1wkvyWzRzjLsbwUsqA+YrRXHaf5uMO8UMFlCWDxKU7h0Uj
gJ9WkUzmHRykchmiBo7jHvy77No5Hl1inmpXX1nM/UouJmZs9xib9VbfYVfSpVvc
anMY/Nxq+o8xvrJTjql1w9skxMUmevh5RAmxnA82j+BFbXKCqc2Enp/JFraaMDLA
fKWeYYI0XcaVL6E+P7iEmHIvAsQqQN1TK0QOPszGYaS3KibkMllAlv64ueSsm3/e
9sYyD5eLLM1NBWqVQyUEX+E+Yaue0N+NiUbvOVqMMtXqdAJw6Y1h9I3bl9Eq1Y8v
+4FsCI7OdpG67RE24mJ0MytP48ltCo5qDaS0PzkpVfLzA23rlVxxesWOBfamo3Qr
WdB8oqiMZnl44u/wKRo2MV/eNYZ0ITF2lVWswdckv2Nwn9qkGI4JifNtRSxxkDGS
/xnx7afyTuxlrpD/9CvjdP28cy771UHLujiHr89+Z5kRk3uj5zjqj117ymJu8FwX
YXZvBEgxqZdVV6SNMS6KLHamtenIgzfp8DkLAhCigQFNdKqulmUts7RmuwmNDK2Y
xEZ8QTdsxtmW+aw1qtnpmXVG+Ndxvmv7XTatkYDdsfNOXUKk9CxxrjfGB3qhzgTz
jQQZ6VR9uUbVqsQ23ofqjhteCqnZJlXO6bmNo91jpITGSKcJxCZxI5i6i3s8+TRV
cmuRb0jh/mbds+BUzvOOY6PXXvmDlGWuX+5R0aGTtymBhgj397NbLPrZ3Iqq0OKK
VlMPUbPMBnEYtbGj22E6cAYJl6Uvg46LFSmgHupYy57jEUCPr2g+dmrnjqt9nH5u
InsS71WcMVqI0jfKRL4J3LOxO/Ml4zyppan/Sp94B7jPP+H6AuWxboGZa42DQ+mU
i9CWkGdlXpLepOD8hrlAcS379nJPMzUokA7meOdYPPWjWWbvCOV0m7kWmGSu17rS
DA/rvqYAdjzrBEXSveV7tuGVruaZwowLCSOOTd3XhECizv1lDpdPFjD3Kjk5G10/
Bm0JQd3yD3RU+tXIYwHPOeMDl9/ZZApM+TqSEnAnqiTwQ69thahMjwuaW4nU1ome
VrqesZcB+weZzxS2E/2Zkle8Op8FhJ5elBtoKugepjw3s67g1DXa4ZdIURtu/KSl
FRvSgLbqiQ8v29l8i36N6lhVXAMJdUVoqa/BcWOqm85gdjqZlKjyYWFi4CSIHTAn
BFqVg9Sqmr7V5ctCLmsPQswAzWszqSzU/htwUIiU7EzssfVku8RyMS0tn4FPDDI/
p78OE3kRTwHjLrezL0xxGuQUt6uwHCQ5+ffWc/nZfU+HyHGBPFETudwSO381jV1o
0sTQjz7o4H2hW76t5+1wQDuDMMTdRrENLxOr0OEvkrB9ikhgNElz++LGEFdiVGx2
tTpLhPIA7Bczv42ngfd78CtF1VHrZrbSSCzsBsmJzN62aUTXYsb9FYIfmukXed5x
T77PFKbQ2REhpclOsE9apSPmvPD0B+ZZqOy0OpGNJ3jVyVyUMmHBoqnGhIbN3FSl
fvjK13OEAW5tbbkyKxM/nRlWhMtmnk0M+nVPy0NoPL4e1rahY6AeoXY7kf0ryxV2
Ph9dZ/xgrKp7i1wSaCq6qqctu3qeAl05qVMeT9BLRDX2J534X+5TXnmEHgmJcI6N
DX7UL36/EDv71EsgPlSo1oG6H3Uoed6IxmY1Ri2/3b9BNwpTJ4I5BZqP91+tH5rC
bPcknzp5wEuMINm3EqaKCt2WWpgjCiyOotez4q7t4Z8CzmCPzaNaGlhPr7ChBYwu
RMM0UgLqjNfsnzTOhsclOI7l8mCFEtVUl48mV+WtUwc4d9bM4m5G2jbUVB2RhXyD
dhdTNq4u8Gf5P4+gvRVxIt9QWVxDT4kJTrdmSqyYI1D46jedmPcUamP3pkTMz/5/
D3KKEWGu17xYKI9qglHXZH/j8ES6SkYmq32xvxaeJ7O0IFit6ICfy2c1XxKos3Ka
A04Y6HL/Vio2wpE6k63R2Kc5Z+LzXo5HiqoLrEGtnUMJYU6kcWFTsBjNwFdRx7ig
x4olhWvajpCELVLkd8J2uS96Wj+ChRGkCOOnv+ZshpxWD22cPOSvjkdtLvczLJbT
BNuVcEv+7kFAh4jLOjIzkhY3djNRa2hgkdzuAUsn6kjjWqRC+r0u2cflCa8DSKb+
iusIPnMTvh2fVvb0YK0TV3u61qmAetYCS7vHJmvxedZBWCH4NVtxu6MhKM7fjxoH
xzpO+vrZc4X8a2MNZMZGBqzAU+ifACrc4Cx3LvEiYO0S7HthZckfFfLc+9lYmq2o
ChFSh3rNWcUbJZsOBFzwRhdXQm4RtNbtSIJNVa0uU9VjyH6OH7T6BajJqkyVi517
aLnTihTWo2SiiFK98gbtjot7Y8KsHqygsajXNullKDAAnwGyEf7kutYLJkQGYiw+
QBnRBys7isT8aynv3F5ItnFWmSog/nbdBkOcHkibucL0P58QhEHjgBlHNUUVSZ6z
ybicbzPht2r5hRBNbAJZalEE1mq9/GGj9tl+UveGdncGVCnYnujhGt6e2/u/k4pG
lGjRab6R42RgQQ0WojYTTtybtDJE5Yj0dvYVRKMkOahfXLogh3ks3wBvfdtGV/4e
YrcpccrsApQC+cuAih3h8Fvbs+bVbmkDjY2CvuNXEpkxxnHh1Snl/YEJjN4H62ut
3wMbzxGvg9CbTN7NHovmUMQ50RF57eOgE/5f2Pe5hd0F18ztW+AY0LIN/T76rX14
uasMHgDRdle7xOq5YTiNP7toUTRXsmkLlZvrL4cK2tQHNMMgU2JZ4LLy690EE2tI
pf3CRL/gg3QTgSC21b805sKj95XdMZkqABNG2jGipi3BCbcGPkcjAuf6kTjC+dhP
5QiCw2pnB2E88cY/t0GbwhZEQwp+Z5Aqt+iJGg4Cwzf5+49UjsSAWlt67ElT/5Ub
wU2T+Y0G+MgGxbqM1rsmiSd5uU6deD8ZgSLpwcuTT9sjbl/90AULdbliC+PUMT/7
zW6CBY/1X3svD78v7uVP6se/6ZLho0XJz6ji6gVDiowd7buPMoV5KGfttGyOFzmw
FbsbEevjqBg+lmdQTk5GZdgC80rXx+W5/XH1z40+ytfrZMYm81u+POKDd/m1ScC+
N9bRyz8dZJFlpohdoWYFtVlci3DkD8vrdGeBFa5hoZSzPa9Ys1FNm4jjhvGSL8i7
xuPcaL8iFtoM46IbXB/S1SmNpWU0dyfLCzIJnjV9ie2+owyU+OOOIgHc/zLgSpfr
QimX/6VeB0buqPakAvfYjV/G3qUsUNm3eYza/bZDU+H1S9KuxthuR8vzeFxdWN36
ov1ohUWZsGfHwxYGLnXOUPuGAaFO0bOeDIcwhHL7/XbejLuuZLkowK03jZONvY98
gIWR94gyCDU7+1LDAWg7WTw20X1CxEJpb4VM3yXeI3Vta7HDdee/4cOHRi847MW6
uypGeMSDVz43lU8+JJ6Tg4y4KSASiwPKcfVSyJaWoXxfR3KB00axQtEQHGHq2G5K
KnKsp0sw3CePwCnG/Uov2OzUP8BKNUTth/Q4AyGXzZrOHW5b0gufIiWraeFd4AwA
PYqbL709EWNgBAadQAqcY31YXa67xk7KS9fqQzmB4v6wI8P8USaBC3zVjx5SC10O
X2zXjAbu2aYZBl0aYmlSLyop434jmJ3uPAaNZBRenwZz9iWc879fU34AxlK1wZ/s
Fg5brmFxu1E/6D8UF3yMMVsS5VlwclaJwHGbfT0KfnCaI3y2TEVS44g5SgDIweVb
SX7l/vyjPVkc6yefILeaSaVHSfan4GEWHRIWk4suKlD2eBC4MKg16pPsWzzPLL7T
+j4fAc+cQt4uN2jNXsvPc0I4AjKmqBIRzT13EFj6ZyjfHM1CUrFWfIeswrT4SnUt
UQGy3QoaAc7ibE4UWuwYSySIZWOlErT7Ge3ViCyIB3cnaQ7H8yre3EkFGKAGx+6V
ZcvOsZispcnwrfa8fAyac9Yft2SyX0GtNnnEwq/oy0Dm77mMfTkiEVcZUvlj+nFL
JNrms5nssHZF0PZq5Epk1WMJIvgTXmOf5K68am/YwJfyHezCLoKWWalT9EUClhpg
0xNPts8h4f/1cAsbo9eohh4U7WxlAA/eHjyXhaMW0/70ONtlBfetPcq+uagda7qm
1S9syW3c1RcAyufGvz6F2XmrWBlzURzzxp0gA1CvLAEOKT20/+zuDH+sYz7Fbdf8
/bYy4xfcgQGujLFiNiLruT5CTEU6qwRVt9jIZJFXYaAMi5u4jxF9omz5EETvocVC
P0EfYHV5zluENHvbz53jA/mEf2ltDqEUqhWUWNWctEZDD1d5nyIl2JTr9Deqykn1
eOaO/i5eINcRIQDkYmpqQhDfZhJSDaNIRvmiifWKKg/KJfV1AKjtdRXYceVyJuTb
n8Fts7cXu1dg+lieqy83/sVUQbUTtbZCRsJH2jM1NSH3YeQwxqSdpSNnH35fkREa
L3QbR3ADWep7jFkJBzhMRUdL6sw0VcAmjnRFqTk8Mgt88WbDh9rEyzaSliIrwPUE
RlBINeKUvYd8yOSSooOe9qOZZiXWRN7k78a0bVqzJHCzDeBnkGC5C8ZDO+hWSfHg
Im+MbEe2wGEtXU9UwuGnPh+opMOw29AFcZognAIQ4SRT/vQLCrnMqbZCmKRjn4Mw
ttGS0qN44vkKQQlmXSy+7j5ooKRsVyYpuf/vpp+S6pLMIqrpPUq4n7+3NsuSsJJS
ahOro+trkhda3A450vkLwLxIQVwwaiL9mqSap5I4nN5Z1Krha7GYKgYwG9+TCGXG
3NSAi+NWRFK4Elg8neZYI/6AWbfRF2z0jU9alF7NHuhWLV8Pl4n/nk8GvjEpozpQ
ul4FXEWhhDh1n63BTUGuM7N1yyaj3l1he65byZoNiQil3gNlpaIfuIJ2LbiJLro3
gLKZYtA5JNT557NqkAR8WWvAR6Lf5obyG00PKkHPqsMitbfzIs5nBgodFFtmTCrf
W79QbXCNjIjE6PJ2/GG/8rJmSz/UlJ3lEUU4DR4w8NLwu06HfjUDccMzwHz12431
BxFfCvSoCteeonjqitNm3hdDpXL+10vFElvqw1AStOq+YEaMHEdB4jcf+BMQVDH9
gswPq31oF+e7ZhRqatQ8YTqkS0PgkSjUAb/0OzFj84jJntLZ9YPVu9VaEgA1sRI5
z7Uz99o3cpbW7WV3OyTJhP0rcuAzTxzDMmkNC+pqpT6h54HFG5Pau35oFtWr33J5
Hf/pEOAEmomKPDCFmLiyGu3538bBQfXg0UkXe7k44qqjKDbOy6q4J8/qeuE7BGS9
FaHNMhNPhvM+XSij/1ZZeNBhK2Dfo20xhU1jApOQ2VJW9kO15e3wPJl1Gfun/FU+
1BP1IPBfU/HIT2eL0kkleuN7+geP+rGkMcnwlAAxg4sAbQYnKEr9SJyb+d2l8xo/
TBXnC+a5Nop9LnKKlQUx0IhTW4yM6wKVpc9ooo7+gVkzY5wP75Xb+SeLC/gP4SC9
2XuylSAvB+X4AKLM54HdXpDxBUCR2L7ZQ26ykoKNQW0hA2nqDAfJ0SXNI3wFJMmm
VkAjTlCzYRBVy3twBozKrrH8eRyRHFmzinjtv9dlPR84IGi4JEAaLM2YJHkGJ+uD
OMQxR1zj364vYRuofFUzkkeUlSR5fVDpZs6yAK3043rfuDmNWW9pUqQVlXFbcfYU
5FbzEk8NB7jeIoYmkBypwIOiwAFlByW08z4sBi6wHUH8nxsZlLMt1zkZIXB4h5uW
09MvmKqVccwpk0TIwci/1w0gsnLJTpcc5e4m8o5ZicAQTJklexpit/S8Qy7z7SVA
aN/sOWZ8NJnxqnU4zRND/WXaHnentW1C5eR7ngIFv0Rqx0A6re6Ma6nxgS5keX6J
N7VSM4IvSW3EUtjvAlTptSLYL3WWm3soFmvLBIDHwp72GQXovKBl11+PPeoB9vVv
eAUIThHL//ao86stGLclo/fkhCGpFspzFW5sRV/eW6bJQwkl70Qrjlk6Ephe63cV
vKwClY9cUIxrGSB+wwbSpgABtKRV4y+RIOYBKSnZvSbL2KG7RnG+uF3dQsWdmEJb
tQD05EAlWvytxdd1neu384sC+q+aZ4xJ01Y0XdGmFSSbPUz9s1Mei9Cfh5o/cMkL
zfljOAe6drON34p0KRG3yOJiT5iQGhsqv/NFigl28vAqtBWBmEMplc75nIwzSOlT
pjtF5ST6XQZfmdDsSIkaDszuAiWdjBuTknoCp1ispOQmwEvY590pkGipOsXnvzeV
Xw3RMB3/qz1rM+eAIXOMH+TFSqcw3YKr2BjIux5RG6kKd9U9Q0PwSm7ws/rMtnGd
tzQosAL9O/o3ElX6HqTYCREAowOsSluwRezrO/+TV7djdrUDBMRJFPKjFngJs98m
lQAGqjnZXvcx8/ev1Hsyr9NVVqj1ZvqkDgIj+e8Bte0hceGgB7DNL40Aj5Et9j8v
syUI+zCy2BFSwiPDMcjWCMpOKOtUEN+HY7TXmrsYqNOaAXc4xfRROy78j0L5P+nQ
Bbrhns/YAWUMcVBZqVsgs6bNJJd3lHNKa01Mjl+Gr25u18dlks+nnsisxxHbhHTd
5KKkYeiSW4MlXqb33VsQmb5Z838XWwWGjN/fiDLRLMjjOqjl6pqkMxg7YrJFe5Qs
zuFgC2SIx6NhOv3FXBzZjCkzYuGAHKwJmLF3CyeOfbghSP4neyPPDnz1YBvHSQTF
8mol8h6lKgVqhWA24aKy1G7wPOEznbjlznp6jU1Gy7Wwp6CDMVYQsqywRZrWcxz3
6qOYi4lRzc80V0d/eOR0QJOg5BHWxlB1Z+x5Oq1e431Njzi1RHNkEkW81L7+q3si
reFRzLApz7zFRLHC3wkbg6FtioYqkc80cjy89ITZJ5z2R0Dw4pHt21NUM5W9inM1
0bseaUcWXMkM2uen6ICT4QbVVnSZ1lGWUW+oTVk6Bp/KrZyx2L54EXqwy1MrX4Kb
84/ICklG0DdYgBSS765CAKfO7gOsYR5RE4AxYydbKg/jrdddblnFqHzCK39P2y8H
Dj6x2tMvPiuqj7EFOkmA4NxhacEdOMKa9lq9yBs5DHLY8K+zTsYgEjMksw4m3/H9
62RFV+LeK85m+x0FLnuFbqBhN8lY+TdOBsOHGioPVm84jZQ6vlFfFqMIa07GAdYS
v2Kd2F5Z/93enr7TvQqLCGXj8AVeYhkhVIvEfi/SMoOT+IULA6A73GbzwPAfuixO
TECQNn12gdjimJ/3+ckbNKPUnuIMAFQiSVwGFwMob9D3wpjZ7V2VTascbbaMNX5t
ruOQpjk2SrY4jZCSgzWhmoiEquDwS+1bPTwn5KLYpoYVIr2UfWWg7UMF647KkFpe
/Ervo/ShiYLaCyhgvee5tHfJlkotsSF+bYpDquSJ4JjxnhyHmxum9OvfDpaec+le
XvytjhEANwx9fbjbLxXnT3ogtpm8QLdP98s+uP3pgEHyA3FuZtMEl1p8kAAKsNVP
SaDMn7zL8utSEryyw/5FKZ7P5mA9VpWa2gXnvEiMCSzEOe9SjWE7WtWwW0JtfTjr
HhLuSQK4qhUsUBM6B5IBxMic4nxQ6WHotzklow02oicGtz7rJtqZabQq3sWmedFL
QEhU98NFtgAlrpvQ+Omtu1B3OCQBq6qBN2xyuV6eiapAVBBoC/mjlviFUBxLMV0m
mW1BU7IuhJ/AiZws9Vi0MopU/9x7sMpjG+S/x6rRJjWyaoeqevAVU/ClgxujbnEP
c/LvDKt1s7/yMcQQgNWHlHmol6hX1/vJLyU1sG9UDPSgMHb8mDMHjafCTXeQZmAa
3WZ7vJ9UeLQqqu0XKYaMY602eHF9/3JBIoOSt9P0Lj0AeuE/tT0wq3HUBv/0yD3Q
ZNEsdu0v2WFuImzSviA/BE6olibiSLVjOprwySNJiWERgWeSp+7l8roweGlBot2f
8SnwLGLAIQKm0KsXz37kGDXdgimzjt6Ayo4If/SqkG1Kv0h2ZYoBEtp7Pq3b+/ys
8gwSNFY7ABoyrINWQkPWuIcEuWuFlRcLGPerd5i0CeblCGim/KeLLbb0/Qv2V0yI
tlRZfRFoJ1kOXFbh3EiG6ByU+MiJWebGyPGYS+NvSg78AnGEcWgturxWFIYWJ9d4
DCOKEEZ0iapeq0mXXD/uWJtjHMEIOp5n82z+I/d/Idp08mbsWptCmfAeKbGELFMG
bg3ClzGcF+OyJDdmcD/Cox27kPPLVwAdfwjVeuc/Pq6PavA1laMzcHj/LN95Q9SJ
ZriuKgCecq8VdLikYzkaGHyn/Mqxw7ZKzmQYGNmGk9EH2p9KwFxGyQhkSoWRIxE3
vvR6WMZEMsuSt72hIkzvowFjvWIOX5JLbEdVbg1M+WR3yDe7CiqWyP2zH/rIvxD4
1HqBlwOQYIyP36oze+0SGPl2018ny7QKVIVjj6Zi6jC+tFzWgEFTgN4Gr1sLZ7Qx
3lVo+tI6c4Uh/VQURvt39qfjYXoDLJ2sBYaVvg+GNVhQi3x3ZxCRR1olh/z21unS
zSCuCNTvfdEWpDWzMeQr8VQcndmRwp61DduhZMRYZ6MbNbVlihnnaDBiP7+hKlrk
BnE52WcssAvIxGmo149ykjyGZkbCgwomN4aPSlHWPoRy9ps94rxJh/VdO4EaS3Rq
qqIEdyS8Rysh2siNgS3LPTdd08y33sDUtYwF64d449feCvNg1KuVOhY7MmqRqpfH
SBtldX6bSQUGkZbhU36tOSSB3cLVdtfeNLcUcrrUZjw7FkP+bzoFTVCrbLT8fvPk
DMIlhXyx5izbpX+XVwTDC1xTQslanI0VrNm3jriD9UHp1KIwmrKXoPlY1vDcjHrf
es4NJbl58cIoUsj8RHgUl4MzxaJwowAL7AMPkpaXLDfThmQNrpG1mXAQ897GteLo
bYRjxagfvixSfoKgQaNzuflyzELUN/cU6i8Z6KTe/f3RBIO92EFc5Xd/8ntmmX6u
uIPy9mosuG4A1Tz59sjvwhCGOG77+3UGVyMLDquwRj013FNWyI04mD4JD9Gcx2eS
nEi+u75lCC9FWtohGl/TF8izWnJP5ikm8CFzex9BiqvvPxHA+74HhirMshqrsJZX
7dYM+8v6uP6Da1QKMSd1tt+3a8dvl/S1RGWg4xBm0JK5PKc8OllfwdlAeJe2UNhu
/qP7++yXGjXMw96jztkpCGdubE8x3PzMdXtqVfAyMgTfXwEAmxFeQSTL/vtLhz9X
ycaIYoIsrxjsCRcdeRGbQGi6sd2P/pcj7Sw1Lqi0luV22d54AimOiBPfFEzE5ImS
IzV0t4U9Fe6r31QcaFilFiKP5P9VuYwUf14HAVThCSoH3cb5Erv4FmnYcHKHxeJ5
+ZDSRldhZmbVp4ew9UMP7xSwoDszHK0ahDxD0YUa2pa1420rYtWIhdfrzE9oNYKv
yaV8EDqzfQonGOitgQgpP882yWePlsSTApdc7A5sg6ihBjTEVNrtu9xza37tp2yi
H5C3lNJO0j6W6nJiqX4dY+cLOQAZ7FlU/JNyUllrzYl6qvM5GaPzGaghqtOizRbK
XSv0KQnfnALaOvvscT4Dtj2gDfT/ikb8okHml3E0AveZTz5jRFheyKc9rAdHe6Bn
skAs+JU49ZUIIfsoaDtb3NcZ/ztPRa1sFWS1IOPBFxTk+p3zqpFJ9VXLDnrUBsZ6
VKQzJIXCAt2lcUUHL2TYXPyJCauFggcj3CEUE8lfa+V4m4vc5xTcuY6CGs8Vob0x
DK4fUNbc/F1Lq+vqifR6lmAyyG/FAzAw1+FRszvaLOYNxhHfyvfm+RZHAZvJE1To
MTu/1cBpk0boCfDiD7koNdXMmBxMOZhcE3ASrFbe+8ux5H4Xw8sN6qntOJwNKQFD
a0CWsUEBNeUlIW8LcPtKLy7XclLpyygXD8c0xsmvLazll1u9zJiiyL5qfIfkr4+1
QrJXtfsSzmDPrOlMR0Q3GefIDvJKARRdKvR1GCOTXg3rfaGyOV0rfKLbUp33RJlS
oNQ/IoqQiUEI/2oNc2/c+ccD+fwzOyEDWXrsnTwm2X3KubR1WNCiq+Fz6wNhFh/C
J1FSfmfV5UQrrIDq1p9CAuHyj0PXak8EleOETpLSd1OAiH198+JDWsf1QVFdTppU
MluAeC92JadSFd0KLKmULvipmCK0SCYjHjY6v1x+sJ868NolLUvp1GnHxXrSSh8A
7ECvJTDe9+cRj2dc5FMBqg9xiuDmQsGfWtXXnrA0dQQaJgMcS+Qm0EUqQBShShG3
HWyV2IcWI40tN4aP+MDEsP7xcgXPBfxRKETBOIqaDw5eRiL4TKmNr9o6HrR2GMQc
c8RmfB+Hq5uaUdUgn3l8wA6Z/LDGDJfhJ+mFaGS9ZwOCNkbQMaXF4o0AQyErZGOo
WUny0EKsI+5HDlJyi0qRS89F7fOk2J2G3HjZGeeYU1Z3Z9a67Of+aYlOPwwBzDp3
Oj13aQGSnwSs3EbnxHUaiCF+qh2486UvG/T0tC2hbSeaqEydq5kOPZA2iNtRR4ax
iDnAzLOVrancKfUgvS1ZRsatdboOMz8aRibVVr2rNA7uvUrvZgEja24nnO+kgMy7
779EsuROQjs0JFGY/BoM2I2ZCnYrmL4QcY1BrgdLpVGsNrJrnhimPHOQdpFt68Vg
zJLWEcITARu7MxR078F5gxGqVG53i7KwfJ4v+YYHF30chcgzEa00XRjKkYCw2M09
eKA6kyrjbEN5s0N8L1ozPyuM/gw9j4RdW2kMG1zNowpkL32DEQKUvNEhkBgqfZ/7
Q95ROcCy7JJR3eEglRYHzDHH54RKB/Znuz3H214FHu5ygrOKNmO3xDP9vtXVsVJP
JmQzuwSU87YFMv4mVMeMJyBg60KbbheIbNmrJfdzxScS0Cp4h4jmf4csImpFeMO/
XdjuUxuTGFYbFI+HCN2yO0yl3wUAaLTUMsdiBnH9mCxukymnZHoBrTgT+qbrrGMr
d+WyMEzMf4I0aVIQ8M903ijAaW9Ynm8sDekgvRHnNFwgH82NAJ3j9Q2MDPK6TRYZ
DquzzgLYbHH+SHrFVhyJzwRCUiis4gXlyhHwd5YuyDJOvztOInCej6I3KGQ+OFh5
MFBC4HDz45Xri3rEoApY2DUtHLAfSbUVGmmhhpxnB0qziliU3P3Xrib615RcnwvO
POV1y3olu5xvIr+IsG42wACi+aMEvLd/rSq1uoDgMYseo6QdKpBZBkGlw+uQ7rrl
Znwwj2ASx1NI6reBVGTMxO0KTThKfiuyfJ/vDMweAonH8aqRwijqLyyl+Cypf9/u
oxkG5DH5Zk3rA2C5Qp7K4WorePp+apP3GyIySTEeTet2LPIOkGDDmBL83l1oCT4V
UBjdtZitEsozlI0w9wOPgyf2mDcqr26C+QiYZ4O/iqqY7aUf/7NAleNUPTbO+KVE
gOr47nbR+chWdpU8Tgp9doU47ViRfKCBZ+muT/XEzzITWXKh48Y75hSvFgEiMZtm
ff8ccGYZaLu2/RShn8kmdI3FE58wuac8iOa302Jy5HqOapUYUJ9FMxfBhhlC2Kmj
gCEReTR5MWKCLpzaT88whmRJT4+NA2NgqbibIjOdwQFizmdFwHsnrY6oJs3+/GrW
Xs4slZ0We3x4lw9tf+UFyYbk/whj9r8w5qH3aUR91Suyn8QFvfE5FOW0xqqEPz/T
B1NHepWH7bdhZ/E/Uq3aUh71hmcaIxeJjkWipVBgOzVRbrlPzfNX5QQS6dHQ82Xg
SVQFtuv5cMHSfKjvoZcIapGMt+AyOmshlB7PbRkM7KZBWLdp8uh/VmK5ae+6A+s6
GRiPFl/FIOtWMW0MxIqt9Kb/N9dojnEdRQuYESEeO4Tydt+nd5BLXU2UK370VYTZ
sLyIKWk39xbV3oto+SJ7fKd9X7AmChR6vDoQHoSIJbfAHmk6SiV0MBurMIgAF0x8
+ASgTjM0Tv0bCvzw1gePIAuCjKjZByQydn0KBXO2s+jIoqCvuQPzwBXC9prvPCtH
h7ZUGgnDVkjUgeLmowQjCKpE5CFOq9eqKa+bY8bXZeJRTsgsGhdDJ1gzQTaPCtgy
QSqWHypCp+WIHbl04Mq2+xHoFcUdRj0uloFWYv3c/it9Y1ytaNC0zk3jPrMQFYfo
+66xNFL4QegWzsNpoGG+GJf/TeJFpxZWumGhUbekOKPxGZeCh6u/Xy/jVZHqolq4
yhdD6KIzbbLDAP40orPW67ARcxHQ1Jkca/DQ+EuH0oqXgE6FvV/Lrt1udA8aJZir
+jJyQfZtLj9GggKnHPVgE7PPKiX3nLf1nWShyHB2IpiGg5A4Ni/UEJv8yDO6Cnha
T/lnpB7VPbUtOC46qDGBRRBh8oOFsDniKZErvqRux+OnqGo7ZruK8yL+XoN2ALHn
iSk9PgV0kSmDZ989HYLxxbHcuAng5TqPMvcm2BLSurP6kZzH4zfzj9qmVVd1IJsU
sD82AAjuzJd3bDeANXLAVt5k6RSVinrdvEu/JzIlJIlY9TaW+n1zBXuAhHkI2rEx
em2/3lTp+4GJ95gaVO4rcUvmeEOoMVbVRPbSh4Ts30+b7+/mVGSVViUR/ihjQAzl
PCmJBKrSwX9SEdrehdii7tjjPLWHRq4jclrOTB0VTeDr5qcYQ784MORDcdcAJEa3
OXfQcww9FOe5tMF39NnLMgg4ugDWwIuLpbCDcRIP+N5FX9MEp6EtGN4IqROIKD/a
Ysy3h7O8iVxikAieehh32Ac1jqZ71nUBFi/mTGJo3KHatUK7hB/MeXT2wRrpOTjw
AqLMHc6OWgsh3jFrqZ0Oc3E3j1hHjXwilQuPeqLn/QtTVJe9exRwUUm5Iz6rIRDW
aOD/nMQ5H0o3S2Blifjur6ADUQL2Rt08zJtCPwCIHTd/zDGxWRj5E5f/HnW9Q1aC
Sh+QeDxTMPUwAOKdioh3SxxR5U80kjGG2WLflzwQQQY5cp+f3kd3lWP/NkW5LOPQ
+3g5S7/3P+1dJNO1Ici9CzP7wUEMgc/CTR513rjT9v87YXFvn+kgwxQQ0QOiBiBT
roh/ePtxINWaLTIy4CZeAsFyxF2C23uGm4ahWGzkK0Xc1S4nd40vsqYe5VAuwVl7
Rr42Fm2c3UNHIcQPP8rzMXG2dEXzpdn/DWF/3u3UJTNvRX2UAgI7PIscuskS66Y5
sS6XYCxnazwYdrrb8yBajWz+hZcwImObzY+QwOsCgyUUngYwXcfgTg+qHPo/gpxS
DCZGkJpkYydvCvLar/+2HRpIEW0N5/27VlSlfA4wNQAakO8dYtfdeFWcMfbw4plo
yQSG0D3DFB1xqIhV+Bq4CGa/lO1S2wgzC194sa8XwI+fN88oRWEYB/7XCk9qIUSK
JK8tq6/vE5HZSf8STUt+Lv1rPpa7egN95Jc/EeEX8TMxYlVxeNZyGbFj+Zz95RJx
ixJuGghFJnzosAzj+YJ6ZBoAB742c3j/u7bWFgAee01kCTKS4JAXKNRQmEbLrmmQ
MUql9o2lXiAs8PdlTNM4aSdEfTYt2OatK/lvzZ5mcBJ9XnRMaUNu9MOcgB1WaRs1
e9DqTZS6EMv5OFn/taa14fHwNQp2ABPt/XAsHDP00Oy9vJu0cUNHFBTOmbyD8L8f
DM4v9ZaW40IEWanNY6nbTzSqhicgquuBMr3Ef05UXEwdFRpvKmPyq6bShSJ43bXD
EEON6kC07yAPDHmVzDzFj6dOH52/2TpiFsjVBBs8ctzJEb8K37xnY2XTxc/hpEvL
DZETAUvJCLlux9bQ22K9zVFrJC97NiW8Z4odn07DaNG+OLSFPcHC5ecZ8IzPfY9K
I6SPGejsNEPvSNRrEL6Avemi6zQ745ZAA3e3EvcX8fQEnqkP2FJZBIbGJZiS5rKq
m4I4ApGkedQnJ1g0SRzIWMn50NaJzeRa6YeEItSY0WqDcKfhyGKzQo2pydMSSwST
3/DN39GdFGTPmuRqPXXhrpL9iJBDGCDEkydhclXPcgNYcSklNlIb8xTM4S2lsH4+
9iKRjgVBcUGQcbR1v23GH6kqn72Z6gKT5bnZyNw26bP1mCiYaYpMfdzk+khUDg2d
GjjUKr7weyf4zJUXAfeL7uYRdzvrgokRjajz/REYWh/5IyjSUfKtgdsU5xS+x7r6
97gi1fSHQCBZ4Uh1rvRCs2X710SWJP66I0hPCeMD4ZMareOiQPRFPLvImCVo7j/S
srws882ceUbEwT5h+F3Ce2NOMGGT4MpikqvPLKRNrwZJi1yaLL04ZXva8TW9qEJE
nxFQ/aoCHuNcVYzSaU6HKvEPuXVuAh2aBC3HNrFeezDXNO18BAlllrU43o5kaozR
rhf2WHyfImcdtRNwq0aCfd3VR+tzHGKpgUXLmlTwjGdVmT8qGFOMMLJgpNlqsZWc
5QkzmKA/KOoGTcCSCH1iZeBi5goxn8U7rtLkY1eBFI7Ji+PELsnXRVtF/Bib3tSB
8UZMNKHTXynk2G9Y9xXZ3NBviSBHJUtFuO7+oxRfpmmcShNrknluAMpfAcaDEqIc
Z7Kw2headA5UL8OncThEvr/+OLmc4DgdcRvV4hlSDnHWtrsvGfxSDi3w5gBYPdIo
74hRzqbpDI8M8VtaBw9WJl2Bw/Z92lCkKcgmLD56OA5ODlB56AH4fVLPqSsR7aR3
8X48c0LvRpORvqLHXxUn+XH8yFl0OiliW616Y0VK5axD5xwNlHZuWh1b9fy2AMjk
97LTsEGwdlDESVaTbuLIYN2yIKyNe8q/NNU884SLPlb1OQL71U5tDYX0EX3VbzxG
3D/BxUC6dE9AnPHO66ew3SR6VJZq/7X6plxFQnBWPOzoOEgLgtJ5XexNQJQrhX5+
tZDvhXFxfBaHwlAAs2dC0RDie7ecJMExrLnk1Q0RZsLifUdOnInI4Vjb3qdGyJDK
01KcCN5PCCR4ixLDZy3aeEmEVxwR9sxEDLFXQz17LekJC0iqEwEc4kDDDDJpgeIM
GlGjsg6bT3DuD+af3AbrLsLeejKftpgcm6r6PUxU1wEAhtJ2NaUTQYhqiQ/K6kjm
BUlR0mqoGGCV2W1O/TChUPjBDftQnpST/CEhvbzJfvcM+sFJ3cCrUXXHJ/S2bsOK
63PllWjk9VruYbox8WU/oPrgcJ00UKDFzejSchXujVolYbwEMqfak5k9H5SmRkte
3oTgaXhokuppnVOvqAX4jFN+hMTSYtE7z0h4PDcb9IMYBSQD3Tg6XtW9cptBNCZJ
hMk4Tbuevl/iaVg8hA+nX7Vieo4SuJ+PIX9SY7lzCUFAFzd8Di1+v5eUJd7tY8v3
d3Mp27Ap2t4FOuh5MBmS4rcTE5cOk9VuKDUNhK8sGLw7MQZ/NxQ7XkgYBxwdREeC
6zOtVHf65ZNvraIeEtN2RbNFXFotxcScD6QLun/BEEKYIO6yA/feVaLUIn4WpzBZ
7UFCZ1mewWLLKNY3Nqko30bNQZ229FumxD4fHttGVa3NY6Qbh6Tg4x0OlUmnsPGN
hJEpTDWE1VH9Z5tAVL1CAjdAffiHhRGS1F+hc74rVJjsmz7/d/+nu0EIUM2+bP75
1W9+FUaWqswm9ja2/tpqRhq2K6zCcFxBCPqcPM2Z0K4chK1Hb9okFhPG5Ysl4IDO
GH8TIFNY5Lvp6+p9z/b6P03yFV/0Il99OsXTtnt2ceZFvuMueJchb6Cvy1jm7uBI
zhpbzDqVazVe3AsEvmXqMkxFqzPyet3+dTadD81HPqCSzVRJTVFMpgbP5PmMwHcU
EXtcOCpGmQ32MPWYWnpGBLtYE8CQNYh6oPJoapxZ5Mx0FRrNVG9g2tbgGJB2fwgW
K2lJpAmZNsnQ7h43XFrFNyfPvgDnAhD4eUI5ycdTT87/JcQxqDJe1IHoi2k1qrT/
4XlhzosBeaBGkw9lZjird5m5/ZqzG7OsjMme9iQoQ9Lo1lThyk/2wXQU1fohSB2F
f7asEMu1yUmhWegQC2UKnUfuPE6paRrHMa6KOTQuz1UKEn7q2W9nyXzdyjfLBRPn
iWiFUQKc+hHMFpKK/qYHhixRllucXW27YxOzqX/+sDeZQy+onuDveEIroVHyEdyq
AIk8Vern9wYVWuFmLsIUKl7AWExBzMH7Rqmg+RcTqOwxTut8DfMyWMKveNcR+k3V
cWEha54Wy75hcVmkmeW5oq1utryxEJLUSu3KjdsR/f5PPTDSsNrlxjQ3bc2BJ0Gk
uEZB3IJ2bd+B7rpjD1iTyXISf+ZjJXKHjyxKKSaSYRQranbdPBV8z2DPoH9uLFDQ
/AP7ilJilOc3DaozixsFgqhADFZlJV1x+VNT2YAMW29hOdbMZnlTlyLUfoLSVGAi
UeSuzdrsyvBr3PD/mEY6PCHM1dUv+qHBBCoxUh1zhIPfCq0WWbF2MUatyO0ZtESn
ddg2c915H7JW0WnK3Zgs7xPOawCZPygGzyjwZA3zvqpKc8fv3QtyD3c1H6o5qgXm
lqhmVrGqkbK8Q7wpN+CgX1pp8i4lL2HoOWgafILdpWrx9SImDQowV/ubsl2xbHet
gesR8U37oQtby7ZiBYaVOMM/nGbVegHiapAmJtfBfQMzVDL4lMhW5/HVVcm7vYB7
uDMJ5prhSOlGhkk8OdcCtCRx3gXfdoYU4aIIGUKZEPelRtGQzoVXQyUcYHdid51X
IksUM2AVlsCgqrH/JCrQuQGQRAuUoPAyEkqBBRgs7orsYupBOidFHlAoG/8dtm4x
qPbibDyt0j45dQFZ6i2O5+SPOL2ULZOaGzIt1YDqAFrhtnQCz7Jc7Dk7EGaLkVot
VBwvtvG/Wudwm3FcgKDzS8K9l5Ri5b3td63bi+RuRjm0y2pB5Xm9WEojn0ATEKQf
SC9H7Zt5SOCiN/eSRiOGyANnbjpAFlyYLHYr7WZrY4Cq8jTW/bv+ParFtzUi11xZ
ssHUq5ZEl+Ysofg0SB4EPpSI7LrEMNyWI6R1e0+U5pbnYpjLkluv+ePZk3t6aN4q
gbtx2b98rFam4iFm4+m3YG9kzA30y4V6CFM/RkJvlLo1TOmmgi7CmvJZfPu2rKaz
2ZIHvY5GfOUEECGQ1cmJj8kkvXqyZA7EzzI08DpceK6ciORU5OggiVV8vb4sqjix
H8taBaWU3ey9CEiuEMe66lMNdezzDTq0Hy/U8fOmywWElzPsZIf2fM7DEVNXxT90
w2hoVFmfK1vXK4nXLS/mv2j5qCC8XX28bg1DDsein8ftDlpnJIQu8dTW6SA4MKTY
uFsgqz3TrbqrECni6xPs2+6ED5kjbCjSJoonYYvAxgAjFkHU0uTYdungN9w0/5Mj
2CIBoAMGgHV6BFbtl+buG/Byr+1wvanfj6sfbHyDsrM=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:26 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qv/hTOkw52EBgFCOplX132GRagW/sEjYbSRHeL5VhM60+NrR8SDCBif3i0Fr9SwH
HKGTk513buajE4SP5HPbkVQuuQr6FLvrQnrfsbPZMl5fL0gm4EWLXGesTWE3vlbq
rEucOr5tEHtb1XFr3ZUxTlKpkw90UihjcOUjvGFzGBo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5872)
rB3wlz8yxXtXoBwvGngIKi4a9ZKiHghETak7YqsO+VFrn5443i2S+8bg3pimBAVY
hAreXlIpNE12avfgLp5R1gxSGvQc3uc8Khl50NeKs+7dIGXUA9mx+SeQDNmlbO+L
jaIfQKJ8kEK1p/gYEf24OoYXRC+ZEcfbdZ1JRHpbyOO8gPLH9mIgLdbdxCO50XsD
jJSI7/c+Cp/gw+AnqjJIO0CStInZoYCbs2aR29yYA7tDt9rTMMHrZndETqxwYPoI
CYb+ACtWxRragB8VF6LywkMxCZl9M2E2xZAj3IQemNhxotqo//V7GpcTicDo9yuC
HFiu1B+YIz9Idbaovbf8j+s5+k/XjSUYN0DNDpFXoba3ZwA5HLFyv79iCwlnOy/O
VMCYbL0W6lJYwJ06tnJ7jWd3szI203313u2famvmgkefKOjr4Jcmy1EoE6Vip8MU
xsg0ps6UHphirNgG3nHoqdYS9R/ObYUs7iIHJAF2LPpPaKHWNxepK+1WTN3gWBLH
zUvRz6J4fsuqlI6/VROGsUDg2GObE/B3IiQVW/z6PRm31mfA9NrLJ9UAs5auXtJp
fwNNOCN+65ismBYfH0dyzez5G/HwXKJc9y0+DI9w3MP/p76ZmPqT8YQqym8berIW
2tCYa2a8I9iOILyTn3nQmGX9OBvCVHhRCHJdl7HL4h7HXCHxk0eGRZ34q6Q0UWj3
wHZzMfxnoBIfitnEMXfj5JlXDFAN8NtGno7KkrqJazS4L6Rn1HGf/RS+1tGbvPLV
Cx9XZNml8k52GR3i56Ul59ymQArfORGkz115AtYiZzMpueKUF33iERL2IV/8PsOk
Djmwwuy+PiLrqs0A2EFX4lUBlP5vfEnLI8Jod8Ufy42daGEhntNS05pMBuedmECg
nWpR8lHluOE/8Nvi3I6bYxNy5N+ppMYcwsmAYbxq1giE/3Zvoh0EvXIMfHu+dzsL
7C+WKgmW7S5HqXt+d3+8CLsp+7v/AHEX1EhrFc1kbYe9uCLKRjrjHixKwEVo6kzI
Dj/rScWDu1SqVg71MXhan2W/eGbZkJ1uYnLNot7L+d5vct7jSIfcq/yptoTPtCNv
5lglFKf93FTnDmOeu0jYEadAAal2rYmGzNGnrLilAU/slLvNYIbd7LdnfhjUtTLo
6ypuw5iGsoRyW1vD5q307v6G4JJP8IMlW6T4zY/QJalm3+i5wg+Lccc69Ssuf/X0
A7xW7v3Hpsy3Zcg8eOph72qSP/yfsfJtAqQwQpRj1lTNxQK5caPxMB4feZMEBniJ
knRgLvuLyPCBEoKk8to59UWOuTgnl4qixjUMqp6mL8kq/wooNR7tQxY6Beav1ZjZ
M23BTR4bXfqd2qGVyfvw53k45LSq+nRBaIMn35ehfxAUqNIASM08d06OdtA6YQX1
uYKNxfNws+0CiZLgCP2ROLfidW4zqcGwdxKnrDCLenOpw7ags/BKaRndiED7PZ30
NpkkpfwhrMNgswhiPP/FZLmkhd2KF/5dB2mHJOQA1k1fOJYLOzEMlD39dVwmYnD7
Di0ejfAbid89YjA4IXaaKCaOZLzgf+KbfUXEz/fd/8WDFCVZeBl4qZyoDAdiP5o2
NrnRanaKt2zFG4K6wEKHGBq1788w7cwoo1lK3Wa5t9GyPqQDOMAohhgb8flS05XQ
JIOoUKEKpub0JFFAIkbwst2otRGHVdVYNPLQsjKQleO9+KgO7xunxG8VKVIe4DE4
exuq6472E6S8YY53cxQxugiXrMoUzL1j1AWREOIOz3bB2pmR79yUmtgUJwNDI4bM
5HyhCl1yxywDj7mep2mRkIQ7+JIxYMeujGbxDceMVt4y9U/4wSvmWlbbAy6E+Dp6
3XMio+rJKoUevGGHGSeUbzMAblpMxyLqPV0mdGPsFQsVjDyiKNI1nK2IDqFZ1y/D
qhdTKsvAiyDCXTlpEdCrD1YruM55APdf1Cd8wDsLjlsFljWvCvd77fV8AqaR++4C
+bx5He+LEh/fiINENFktlD5ep6sKNUa4FRDwhSn9+vw4pv8y3skvqdiK+JQCb3uV
r0KNvRsrKYaa6tUFd1OJ2ik2c7wb+YsZtr7XJnZDPpgJUfsGHLR9yu+cNeTBIzi5
LomW7JZJAMy5k3SiMsj3YXDOVtBx4/pHpYeTADY4UD1UZ2UyzYu+UTG7I5N7ubVH
Lh79dY8YUcioXeAquPUuuYXws3wnBXmwuLqQdpUC2jSr7BoZ0jNpOSQam6YkEHoo
qECoUBzMgltzVYzFtIJi9tsHWu/F87mxLelhyIgWp32YuIZl7nv8yx2L89DoeaNb
hDFANE5kIyQ4pMno3htaRIM1Mkt8EOxXkOZG4K2SOV8j/obdYPml0OQTW/jgtzC7
r1uprrp1t3fsex/v/xlq/hnGAcSTb265grmRA7IrBoVQ2LyV0YRL65pixo4ntMtu
q+sCtc6BJnDa/vMrC9Aq+fq9wS3V6IMPIlTIVQV94Xx3GwAvvq7QmWG3KudL79D2
h8o1P98ag9PDAWd9J8o98apwKsapBaXf4/bPB9GKcwOKpmgL23J9wcUGh0R7C+Bn
IUe7uyF6YfrbmTIL+lBNogpB1oTPQjpAp2qS6/SjcV0dCbgfvTOxokhI1PPoUdQN
4xqgGAGafL4mIeDrIwPOyvf3WW/CPs8Dx3M+b2f+gxwvNtDkiHM5gGCEuPRyQaJZ
Wz12sC7NJ347jWVy61BFQIWA2XL1NdCo6Pbd6RcGooSaIV7sVY0ZwCWKUlx6g6Pj
dTOIn5ZSrItWn46EHC3t8TsFG9SsYvGqGZkOVuTbxXYLtLLDr1PfKt99H39Lv/4C
0BWCFSXCZ0aCpn5ZJj9J+A1o3Y7veD1Bqjai41jWVsR2TRz2XS/jW+VWhYnUCVG8
NguRJY30CLEry/rv//pr+odui6YxXgvOkx8vjmRZgLDIltzEpa7UR2RB07CIJFet
n6IWKNhI6BsnZcQsFBCqA3BhGvjhuIIqhJRHoFkvxdMzCQBPzs6BeIv8jUz2zQoI
fODLVB4+42fFK6f2qs3aaotsNeVtiH8SSy1Cdc7OUjXpUtwpe4Pj8pG3NginSRt4
VKC+3c9X5J9v5Ky7kXcxHHJVSjT9cky8RzcFg/4bQhBtXB9Om0beWmxg732vxkxl
k36HPl194lBBPNRFEpjD6nJ+RHDUDPJ9zO6d8YIQuyGIcc6fed8kmlBjW55jRhaw
fxGjZ+VsquwB1VeSUtQ2OKtiI1DRgDsp2cUzbIBisorpFVymLbOoRultom8Sj7Fy
CaYZzE6IFQEAZr12B/NOWYkY0mvCgaR9/IBRQDjmB0LeMWapndyKMfTxwRP4+qbr
EjJLSnwrtB0X4OhP2W4koxF84zEK3i9uNUjqhyVNk+wt7auSSgCo5V6NydiKmuBy
lIJrxR9d0AVslmxpdrm8HkOMdT1Vfqbb6zXvtCu8U51d/PpHNRTBMcDnhFm2tPpu
D9ytJK69P1b45bT4lBprQhEVkTXTKyt5r1MaFOsQy0Q3BnKAIaSqjxx7T3YBBIdV
dQ94tdG+17p10zkWqg4JcKpi/OtWuTTgZjR3v4bszLLBxYi/SYt2u8GW2yDwq6Hq
41lS/hjzz04bMUEWrdQBPmpLNwiT2r8nzAgCvMGWVhuDTuYUj6S8M29PTEKSBAZc
wfWx1hwmOFEhmQdzRKEl0pS7xpW08OjrefMi82NDS+d3GgHWN664rzPSZVTtg7ch
ts3JVGWFTTr+65bm2rhipkJDx2GowG3kXU032pFhCZvYS4hhX+pzUJzPTUyNdHcT
7Tn2NWW6+lZS0x6DmJ04oKERb5ewHAg87+7HeXFBiRyZVNLHY8GNKY7AhSHUeYdC
w5PYBEKqO43pCTYLq7JVT6XThNCedp8QmPb4WZoO5Oam1gBncYAbTyEFbdwA1k/F
5GnMnJPcxwbRQhd+0wujMBWRthqh8ESGOyh3FhftTny66W3No4lpWR/8dTGDMIqx
/oRQGxNw7V/k9iLLG6zfSM+N3n4lw3JldeDETeoESMx3gN+qUldRO0Xto6DMlIP/
ARFlzLCRvi32/kFYkUlCJHAShR5T+T4QOKpXs5fnats90hyF/Gx9arlLFIkL6c6z
+Px+RDzjPF5h6wTVWCAEgJzjsoQTsbH64UlSBBVgOxHMfiIVwDWlDhSkD6yuPhRj
CxR5JxT85FYyvQ6Y2XROsDG45NDzZQrsDFFstsQK2lkBgoeHtXeRRS5LhD9huaQ4
NA60cd4zU4tDnQEfMjzb/2xdackkzMt9ZCL3kydB5goFaY2Q62Hfr/yAyRgxgP1B
hOYput176Rtf7WB1T58DJqaK6TAsM/dql+T7G1Mw4jLsmGa2O22WYXDSdcfww6Mb
Nl2pbL1mTsrVLyj9WI6lnQtHU3JYWYuaA2xmKIXDFmV5xm8ObALoa6cHx6qbR3vt
45GMHvkASB5sTfftNEb+8MBONDasbx8/yZVCVi2OQyeGXq7AHENdMNoMm26yvVBV
qy2VHsudtuULVEA2jdQS6S8LRGADZfAXmpB6RCvOUK2gR+hVoVvRuFffer5gQHyN
Z0GrHTHye1xUimg8ZYHoKwoCZYAbYLwIaoTaDtl4AEm19Fpn5OZ4AzBw+N+3afKT
rKl5pnp7BiviG9ISY3y/fBrrwdyNadvllM+2jtU3nqbYDOM0ilJ09Q+ZBPmITtC+
eP9WMG5u65NxNkKXSnFpmhAZI25GQ531QGPu1Ao5yrx3wX5YPN3XfFJEqmWYazyy
C6OkVEj6jrQUQ6POodNug//bwVSYtgtYXQs+5yc7pXUQuF0k7R6OMv8qVEmF0iZn
R8Z3k4qCqZnDBpxh9MMu3M63aO3fHUXa7G+6u669UdnVlnO2yWCudnNZoKHHZsDB
+8Bpr5zm+h1b9aGWmFHcg00uUuywvssDjEvCg+NvhOSxHVU2m0AMDxFLIShnALp0
RtstDjv+Kd3bXudBZyd0DQkkquVwkSH0UXzaMTLWy3vaQeQlcJ97RxB/YE1avoCm
k1PwlJd/Z+kg6Q8t0/xV6/OW7l/JrF9JvvOO2T/hXZaa2u2xvqztghV4XKre/TV1
SjhRv5LnXWyCJ/2/MGdYF2AdZ6ceM1sAHKy9481Eg5GYMtyts75s3z2XxghnloSn
cvn62qZuLNxpU+Hb0gI+jVHo9jNTe3zDwQfj8yc1lyx4uF6dMnNuitXuZhzg/ykW
NraB+ytUtQF8z91IcBkwRKMkY6x7c6bakqJvY78eLTbnOKjYK9mNVKY1nGbEFlR4
DIlJdziCGmr/gMrK15jLtQovVtzxKY18RuI2uUiVJ86lKlfpnHTg7ipv4d3q0Lr+
0DBXUzk4sxHwRS2MxPKjszHUpC4phBRJbC7q5houRa2QgWvevNuDBksJB29qrhUt
ektqzDy0qzVlRn7LZ5ydSGoeIIlkdj4J/+fN4wQoiqyzlGm0LhcZ4pJB/DYpJIkH
PZwsuN/vLkIQK/BsH2UITpGhf1KvY3CQGrEc4pjHc8It+x8XKweFxp0P04QDYy3w
oshax37Hn3ea1hD/XoVWuLNglJ37Mcy3gpHbYRL4k9DwIyzlkBAfO0ZghhOg/kke
YXU319L4pQaVes/1lTSVFRBHV2YEfWmr4mD0rUZ1q+XJaSfdozPyqL1S1BkH/EW2
k64kC+0yyhS76ShIWAI+bs/WoHrCQwtJ6jz7SWXQ8xHPmdXnn3VPghf2RBBZtOjH
lmSavEKmyWrmM3rD2T9axqIbfizeeYvK2hEr4foeWWbebSs23VhiugABYO5I8tcB
th4DNO5rNfmmrucTo5W7RQ+xKsemVjbjtpS6rQyvzEfY9ymtSYcMo8rn7vtF92qF
9zh0VSpHbNL3Ky4GwtNxJ+77ZFs6hgcme1YKreuLSwV/r7AYF2W1ppvsJwqqWQTA
6GQRkaE/uZLm/RAaMQWOUWwTpZcdX2rbnNXOeBArMx1RqstIX8vWkPACVdn1O6fM
+kcBnPgvgrLaz0JFhOQmYBNQ6s9Or/T6ns+0Ut4OuoKeVDktbgPy5Hsd620cEQBA
Ya2FdSVd4MhMJc38MfWMsEMcFH0angqF/eIWU/dJgAAg47ML97RN+ikG/HHeRlvr
cv93ecxBhN+W366exAMMWL+/UKxCHefouypAz6HVfdHgT+oNSa+naGBBUYCv2ls8
IF8JVBSAgqhehtpP4xlBlfrPtQHyt1tsAlYhXdZc28ll8OsE0YwCAvuN2RgWLrVg
Cc9avCEriYLEMcznUmexjwunTZJ5ycYY4TXVPnbGtnT3DVQiRa8toKGrqZXHIaHX
+VGjNQG3xmgm2NX0IhZXmQx5y6D538AQ8PTKiGyK/bwWHk6+41FhaH0oMN18cVkP
uUvt30hUZ+VJUcACzJENXBuXY9l6HbR28o+U0vy3SSvkANZLS2UHbpnfvqXStYIb
gA4xW/H9rM93mVqIMQwAV4YsqYOjibXlKPojNwSIDm45+o+YaBXgdRXhP+EMbSk2
b3yCYZY26RQ76+VTzhW4GUB1rZbWSurMhsPPkZ9E1wbK3oTJ4GiOkSz9Kbk2oPe3
AcKgeNxrwhDolGalB0IbS3cFUl1CNDhr6rpzCOJXGIQVmIGlBlyDDOwud6vQ9EqE
1gRhdHsge8JdbAla9P49eDKCLPFfQHZPI/W5YWLOdGZ5yDXCrzDQEvnrdjw9oL7/
w05t1peSnfFONM9MmnmDe1S4zHVHycAU7XXGSFZP7QDbt+0IqQRQG9aFf3d14l3/
J8yoMDKp4i1286HWpqAP7nyZq0Kqo6OMAIT5dHuPOI1I/X/e2ng9Ik5gM7Tj5b/V
aM9tbT6oO8CcXqR7hjEjLIdlTLsFnxZcfAv0qip8aLeNy5ili6hgh/03B/M4tFIw
/BBYc0IO+AOBmZiX7K+i7dyP4T7pXK6qxE4aUosP8yZYBAGNZigxbNf6QxmZ/D4I
8BrLqo4kT7ihQSzhrJxw8E6YN64EnfLavJyOcm1xdoSd++j1bYfuy29fiAlziCdv
tK26Wp6lXnSN1ukOpDhkz5MyjFrBD78R3ZCA/czz34zP8wHktCv1UtGISfBV27if
flmWRHejn7uWVpmjw8HUP919okEutbZ9L9wLa7drcYy9Qz3ro/XWSsyK2q+vx/Rv
zIfBOlcu0DYANAxN8ka8ukZ516cujMYdEBU7Sv6E/0LVY13QeJcW23iRHQpDqhBt
ufGTeRSrFXCpaE1l5fE4OHUIegrvmNBn4bC47OpUm33yKVLpHdo9eTB496tyH4+r
SPT/XjsZaVny8Rq5VJb19Sx1u7W4nt3mNIJpcbc+rVavJ+5cktXJkANtgm9VhLdg
Ul8/QelbmAfwsCOe25VWtU6ueH1+mu9qx3mhnnb33TdHp7fksWGmxqDUWHCnC+nL
aad2E3jOdZc4md9GTyPboJKxoDS5PvPKuKcwInaB63B6oLM0HvfrwLczbvg7YzSw
IyaOp+xeytWotiSsL9Ka+V0MvGLnOKt9etcmcXVVJs380zdZ+lyOGQ/zoIUxa1vX
CN/lJhlbUfN5ADl5TbCh8K/eK6wuNf9ucxnX5zgOz2Xer/BbqTJ+tLsGYd5AbtPb
IbY2N9tGc1PQ9HNxr7lXCcPf7KSZbBhB6rWnkS+ayES9GpXR8LRp8Ks+lDPzP/wX
/3QrzW2xv+u2tEXp2XWMOoOcIA/is+IUR9qrd4sRwLN/nTaAkr/lK6fbu0Qn0h5A
TShYWSTw7nlIGl41og2hceQ8yU4s/hFYbWtkGkkYZ8k1Sp36P1coJx1TMQwO0vih
lpuVwodYaRJjhgcbnzbOJPSNdICxX2ANo080uCGXAJvJUWQdZ799x522Trm1ZSXQ
rLk5Sxt3QlX5HYFDgKCNng==
`pragma protect end_protected

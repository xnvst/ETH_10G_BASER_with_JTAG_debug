��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO��Ӫ7�)]�Ln�d>j�~�Bۍ��n"�MQ�2��fb�6P�j���JM�/ɂ���	�w�T�P��
N[�=��� �d-���gK��é%��!�&.�d�p�β0А���Q�V��E�7�S�=G\��V7H{�mY/�1U�Bub0����l<�˄�Z�&@�#����m�N�����Ι]N�%
|V[��/�C���tE���UK��dL_/KHX�n��S�-��^0 6����y?֥C�$��1m�ӥ��[��R��=��5����	5����]Ē����*x�5���]�D]i�RU���ާ�a8�r�2�F�e:M�m��|d'qٛ �%"-X�%~0@/0]�#���X%F�Q8���(�c�<�.Q��^�*<[��h٪�5P�4
�Jj���%�D���[�p��4.<Ԯ�{O�l�8�ø�bH�M�Czֲ�7�B��	ܫ�\y�S���*�q��M�pK6���.U���1˘�� Ϝ|N���w[����~�PO��+o�?����Lh���*Y0�Y�z@�5�R�%��W�
W�+�>FS�R�ש
P�멄:[B��1�"�����{���;�[V͠g�PH�~�m�y����@���x�-�IZ��;�[`���ΰXG�_~�_�l�>�#Ih/�|=I��Q�$�ԐZ���v*s�o3��h#k\�.��i�K��x"?GEk�*Ed�|�_Ο,̔������@%A����vXlʡ�U8���}09��������ްfJ(攳[���Gj��"�������
Y�/ug�x����?���lQGc��,�֜���;g�ǴnA�i*�'E_&�Sq!"�����/u�!s'`n�P�&����<1�!��!f<K������-4.�v@�upӇ
���_2>�A*��&�X�e�F�.�� �	R.��cf�X��A���l�a�;.E\��i�cbh��Y�x��������_�S�/��0Drԕ��>@�����һ���{�iX� �#h�����6(~H���M!��4ZXC���{��y�WS_󦁒��}��膕p�^�p��Y����ugy-�'!#��SR�A\�D����.�(��B-D���v���c����6�k=��K(a}*���7�7L�:��Q����:���ͮ�?i)��){L*��D�'�~kz=d�HQ�j�
�����`����-y�������b?�!�) ����fL�K!������qS2���$��̴͝I�Hu����E������dH<���@0[uαJ-��Q�+�$PP6����)�7&2"3���	�����:����}����9m!o��,�:�~J����y�� G�/�*�&����4�|�_�O����8�w�H��2=�[>��n����^��Z]���֖+�s�N1�U9�\��V�]J ��i��WY�����A0B��pV%�=�U~�oT]�Ĺ��l���:PS����E
͍�����펍�m��Ez�Un��5�_+�A��zߌ����,�y�no��B�!�e.�����"�҉�wӪ��Z�|-�֨�õ~)9N d�*����Rh�/U�ۻ�#��C�jOI>*���d�B�T�5^:Љ�B("~G����.�ғ��^O���Ͳ�/�[*�n�͍�^�7!�J�i�Wؒ�@��]��oh�U!�{��MW.2�U��@��R��.�Sj����lt�]@�Ț_�ڡ�e��ſ�F��H%��C��S���7��}�3#9�,�3Ud�l�qR�+��s�R#eD�����R��N�#n!��A�w!:4EA��p�����n��O��=�ھ=� �ل�!�\�;���(������Z�by-�fs6w� �m�DC���W4��db7:CHmq����߫m�(m¯�R���n�F�H�Z�)�\I�] m��w5�@:Z
���-���`�C�bH%]�o�PH�@�����D�/��"�qr$R���ڄ،��&$<(���!�Dc��͜�?��<�'�>�au-E��@�j�\��J��ƆL=�p�F(僛����e'f�D�ܷ�[jO�tW��0m�2{+3E�|���|�Q@����������f�X�!����?�Ɨ!���"�`�Ԡ*n���&� <mF��I���]:�	F8 ��`_���-�2�֚��otް�>�ӛZ��c��~Uco(�i��x��F�I�6ER��v��U�-?C����+�B��`�9���M�k�RWWa���7>����V��/���74+���1�c>s�2�Tp���!Z��d�5��"`���e�(��m�AK	q�XC��ܘ:�c��)5� �u2��۩���2-��{1=4�)�[4�j;�޽��d�c�"	���'�RF�CE��[w�[�o�vl]�'����x�k����c�Rn��Sп���@�_��)R�@y�e��iI�4�|*?�z�2	�N/m�OY�w_!�L߽cĸ5���7ӈ���1���j�������ޞڃSq��Z������"d|��OrG����B"5Af�IԢ�I�Fa����J����?�mS��X�hT���^=\���>����N
�p�$���򸝆����F1nӃ�&��I�.����tO�$+9��1�`��8�����^5'3�wD�^�Ԓ�A�"��|α���1�}2���ݜgIޓr��,�w�k�l�I<A�����c��m�Y�)�����K2�+��l#Oy�<:n�3)ZP�S�u�(S- ����@�|j�,1��߭��\m��{&�tߒ�(�ڛ-�S�� /�T�TX������TdɊ�R�>fw5�֋��{��S�^e�������i8,�?����Iu4��J�2�	��h؟�Mƚ���l��]�=H�ğC��/��:��n�|��2���UR�j�;T�����
�Z�r���`G;R��^�<
��ڠh��9��i������*W[����7]q�ӌ ����b�����-qK�쎭�ؿtA1��$��p�ύ�Kj5��d���*8��3^	͖�z(�FP���}h� X޵b��dKN:��~	��-��;|�1��A��h�!��ꀣ@\�CG:ct�vw�,���_H߻#n�=k�g�����]2B˻@�-wJ���"��a���N;��]�*�1��X��lC2�VUn梴3C�tc�0���I�T2���1�N�f��(��N",���@r�E���LjO����o}{Ӷb+*�L�dR��x�)���D���K�43m����M��h���O1o��E����6)��>��Ɩ��|��1� d��\E%���ve���A��Ӯʍ>q�&y��7'�e-&��ER����������EV�[@g��+Z4�.J}��ط9|���a��ٵ���J%?I��GPK9��63����(yz�S5a�?q4���(]e�9e=���FK�p7[��h�m�A+�A�hf����ݥ�����[ڙ�Z�;�d��P�Ls�w׋T�:�p%���NYn��U����.'�F��H#���Z�Ni�ݞ��cNz
��<9�k��9�{�՝����6����*c�<��-�9����f*������-��g�a��`�c*�ϼ�I��Œ���l�?ZDJ0G�S*�����N~g8��jnb�"�ւ"���:	3�`o��!)Ee�/�56m�6_�|'��ӎ#��<b��[���bo*}tH������6�,](X�����5XOl��Ϫf��䂮��jN�O�j{���0�d���ce{<�_���D�r�!vE���EA˪�u�$ ��w���E+a�>���l"1��xJ�S� ΃dA%�X��K�kL6�����J���J^f�9u�g����Vt��$�qnTh���v(i�°Ar�H�_��[Fz�bU���*�+WB��G/��ζ�,�n���F#�v��y��f^}J+���$��65������._=���>ZNx{�:[M�A�s`|�F �XB�z����L�� ��	��\A�@ߍ���P���@�F&,#�$��D}���*��4쮋\�����u;�0�K�?��mE$,��?&آ8�?#0�y�u�K�c�Vk��zT�ii%@_t`�[�j�ln���R���Ŝ�ߠ��.�>`&���4��>���p�A�M��(��2�gF7���u��������uQ�i�VM>~��&U_X �l^(++�j�Z������]��#V�Q:A*���T��9s�c:��M�6��V�$��L0��'��]:�������;]X�]sf���T�������&�NW��/��ͱn>���/�9=�  �0zd��U�)�K6�J�X�#YD�Q<a1E\^��A߁[]ܒ'x�^:�����3�O�R8n_)[=��Œ�.Ɩĝ#�\&�D�~̃P�%�bj�� {,�����M�v.�;�p�\<r�Zۇ��g�	�]�	k�ܝ�I��c�׻�Ϸ�h�!+Ȑ�yå/M������k�M�$�T��u*>{�S��'U�PfU�S���������)����C{Ϳ����{���8��V��"{�ԏ �M�ʏ�Rœ�>����wx"o��T!R��j��U߻��Bt7�e�]�c��ĳ��L�5G�rp�����`_�PhHS�kqz:č�$���?����kq�蟹ή���8��b�r���L�Ivy��<l_C���~��ڕQ3:鈕��N�{�Am5m�)Ը����g9V̜����z�v��;� 
å�Iܵ�G�f[��s�]�� ��@{��������a%�\0�z��3�R����:�}-Ȍ�v�Ǳ e�1(؃��G��S?5#�~,��F,�*���_��C9�=	�C���w���I�/�6o3}:�ۦ%b��1G?�@'���[��j�����k B���͏�^�v;S 7�ݐF�[������!����G���F���H�,�q���K�����O�����ɮ��tG���eZ�Q��nz�^�M�deLlW�M*�/梉������xq���?���C��.���� ��S��p٘ܫbWy���v�&L+�]��R�>��J@|��o�-��ufi�P��v��r��
��uТX���%,�O�1+��i�){�gJ�;��{B���f��&|�xm����ՙ�0JP���>�(2�w�G�[��\)��l��ӊ8�B��G:e6���Z�8�; �FpQ����A��m���z^Wv���j
;iFV�t%��}��
 H�+ߘ0�9�բ� eg�c���Qg�0�o����� �M�:ٳ2-��S���T��'ڀ�
".׍�%�� ��b9?���n6�O�vS�A'�^�R�W�Փԯ�x_`�s�⅕ozf��p�Y������ ,�!�}Y�SK�U�������V6����IGwh��W���1�4'��HI�#'���NƇ|P��ܷo{��c����`��b���i�u޻�j[�
�`�xà��r)��-�_c�8M���","���z��7�.�"е�%5�����5���	WL' ��`��E��5�
kߑY�7���ļ;��Q�L/���`�f�(��U�y
���vbG��.�$�>Z�b���N��v�/�*�E��j�	x����W\�q\3g�U�Ji�\��y�.�<�+���MՕl?��:��R�^��.�ŭ��`����qaڌ��k��u��K���Y;HL�G��;��RC�N^��O�@��?1�F���)A@�ᬎ��,	J��l�l�x}�k��(������Q�,��2�܂��k�>>�v��k<�o���a�@�+�� ���ʌ�o�n�E>�95{��%��������G�E��F�8)wvV�	l�w
��Q�g�fA���䄦/B�N��UD�x�����]�t<N���ʐz��b��ŀ�n=7y���R>{ky��Ӓ�_N��e�s�*h��#u�/�c�Z&�Fd~���%0^I����z8m� �=��+���Jy|i�W��Tʶw����`_��ѹ��k��
��钄j�HT%-s����6_岍��@*���%P  !T��)�7C�u�SzeL	��fYnv��8�N,H	Lf)ѢF�^3C&ld�OV|=����o��'�S^���Z�omMR�sϊ���A�m��C.�,�$|G����K˭��ߘ4 ���s���Պ2eq�(��1��3��+B}(5n\�z&=�,��]����$��4>��'��
// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:31 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YUX9pzUbL2cSQzDQBoDMcN1WGyOSpM86cHO3Xbfy9ZyezjdD33jng1YIKA7A9CgV
iT3ztyq1x6zdvGccGx7/up4jG29Sn2z0+0pXPoACUszcATDEBAYbSHyUO+OZiAz6
IJqMPhM476cCbeuvR+IrKbDiiyn/w/GcerS5WcnEPLQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28160)
UL+xpCqzjJ6Gsahpbu1p63aQ8ct774yGydcUj31A5tuP2MoYAC/3uGYKqlCMMxTk
mKGx9H3njFNcCNXC2k0XPByZK16LFn7+D9WV1SYBBR+9XHARL8MIscmmLfNTOJ7K
JykJGyvL9TRBi8/iqUdBjGBihFvQ8QZ3GckO08pGChILOaib4SW9nH7yqc1WRE4l
1MvTpKApakcEZtrg4xTPkFXyjymV/vSvbQmD045i8sw6xDTByPHDnl61l20dwh/2
NOow1oWZPDwL9akmfsNEnr+3gWBfkiyGVP23fd4wQnp10pLV+PMgK4q+GY1eKmny
3+EsZT4+3BfM/itPZ1uWBgRqbvqmbOTjcZ1B9UdaeCDI43bk41NnUjYvYuQ/ITSC
wCz7OOSU4NtipiP9RTKU3PhcE2dSfmEbhDCeY70DZ/c9PvCadGmXnum6AdcLnJ6l
UqIZN/84ss2ylpzo+2tGLbZX35On0bMGvYqGPi6huSBhW+rWysRPf/GhYs6dU7sa
+a2kOHzCBfX5NK+X3TVflyzJY+5HsoN5O0lY1Sk5jj+RCo1V91wAKbzE2eH8wjoy
pbSz/KYR9UBHouPKLCu0LU/bjii5oV3XW81TpbQWCMaJMZjyOJ4ln1Kb8ODmdLk4
qyxAqP2aFtuVUiBiqI5LsAZ7BYpdn00udiVYpW0FORoHph+AJew608rAeeqjQAH7
WiDA0nsKu5RVhA1SVBywStXy/QMtxgzlAwEvZLFnCTaAkyLGyTs7k94MBFachu99
gJYldKKQ+KTBfeTGWMjM7tsD5mmnQIgqrK5m4ZQOLBXKJ8YAamusChF6ji5hEjsZ
7yBsLKXQOBmHK3uavYmONthOFn2woWQo/5REiYgo5TEmIdRhCWsN3bcbcZzgnUhP
TKscvc52DeLKn8gJ1BIvgAxJ6uvuZ0pWMHFFDo2O5qsK06J8ppdZheOf2wKWS1yb
VYInk/kbD70Ln99/ZFMoV0hZFF2QSB3OqJpx4f1ILYCy54SdyvUJPG1QwQCjh6Js
J28t0iUSxzwgTdIDnBZEJnc2DZitZBXJT6BwljMhERxuKxhpdLDZLy2rh/eK3G9D
aiDQt69A5vo4j0Zvd9KPYmhDT2fi2mokqT7KwE39su0TRURROwpc9HqnEJ/rqhzG
dhrTmtHOI5AkavPll5h6C+EuGGvz1VlitVqv/4wRjzLSHGwE8lMCB2IFc6wb6b/u
kPa0Sxkn9X6pKHtdQaPV5USiYOeaojMPIhihW1INWYssrzMV5+Mf3V+78hIHATEQ
xLaY+DD7BinMEtUegHDYJoflIoG4Fb4dkmFMToiQRNJsU+FDhxe2Z7FykuiQRkQE
CtTyw8lNBOU96tBl5gpii9HN5IPJPqFsuaiDTSbXC+D1VLbS0Dj3muBKnsLRihda
6J88BcUcVMjajD0fuZyYyWLCc6v6JetAAercjMVaHLtQjdRTU4NhHagqD7UZSadD
zo1gPjYt+qFZMcL7Y1Uy+/3OTZv0kUQgFnwANOobz84Du0QcnauXzv7yME6tz/RW
2z26uYVSK87+kduQ3FwroBG9CK1oNE76LIOZAHFqcp38Lht6CDbpeRMrl3fowEEs
g8V9rsxMaHNbEDka/13atkewSQx5/r6GKJG9+qFlEOk0MmR+78OdyWAZO5nt9+oB
sxOpVsHsaoL8E7DNzlkHlL3x43+a24hfcs+PD92rhmY5UsyaY2I3iW1yspEYnLxX
o1f/nd3JUQrjuHxlNL2jh0347LQATAAywjSTXOrkrJ3xbQH6t3HtuT9DGsuzuO6T
hJnARYuNzFpzDYp/tP4Rkq6ObEB924OGOAodXm7KItTf3nHxPIVq3y4luTlgVKUF
EdrLtJehKQR7/0bFHeA5hXLXff9lm463ruRL7bb33koWHO0U1eJxqm8fadSNN2VD
2owAWapwD16rIA0K87bxq63YS613B+ENf1BcTwgSFWTDdCM4RlW9ds86wq2HWC5M
Yzpi3HJ5DS+Xz+V3afLPN7TSZErfG1YQsaPQy4mrLelnmy7AVHn+3dVIU5QFfyER
lMRWKWNOD1K47pRb0KZR0W1fEUh1xZ6jG3B5MWAeuycKiHDfcr6RpbwW32JqcF36
UM3kt1qqpl2N9dHUeBddSM+1On88BqMFH0txRCL70ZHtmdTRO/IKOcspkDYumcQO
8jNAiHUUByAFJr/ElsEZ3i02fWzpX24gKAYsZQUvusYT20IDqeUYhjeAmI35oJXJ
/BeDR08a1+QXK7NkCeMRtlU82CNj9Rr7Ii9X5Nm9WZh8DhcDaA0EtrfJjUDdENJH
O6xNbfkoxDLf7rUYJTL4A02QflnjurSYJaxqFtDMhXGec76XATeEhpIuNsD84SgL
O2HAy33k/C88KHuIYrwJDKFWLN5TEtYwOc3RjzK+vKJP6G5fvqdaPCVcV9gft05P
8eUen0Mcw7pwLWQvfzIJn2MUpKhpfmgD/r7apIQdbHkU5ZGN11OkeRfn8+RWnoaR
rO5VUzNRjf7CTdGF8NlmHEvkiXXhcMPVQKdayBAHSN1MtgOstCFPnDVlhsQ+/la0
oynTDyFnyG8qVeY0UFI9PvOXSxitSGrvR7HbnwfxDm0WDnl/4Xz3CXzIqeUxn56A
SP1bFUDws9QIBZ+6d7HEmEkxUW/dJnDmk8CYNoIozP4QjLVOA6VERDy0nvXhDh8L
hfDoGWrK2lef4FLqwgx4WA7yZQZJGg7pJdqYM5zSKaM3VA6BolNhoW31NWJsv8if
kDDaYo85qbuzFSSXNaXyxyGqGIX3wv/Zcc6lRO9n/+Bi5jULkwVfBBCQ0ylqJdTX
VfTkqTaFFE3j1WFn/str/5+O9kLM2Q7wslS9QNFw4q7uBmdfKJh+A6gdNGvlLuVJ
0LzbnIOQ53GoYWTGmp/ANmz9rsD28HUQC6wy65ttBf7dXMrNGO8a7ajPa8ml3XzG
rKQX1R45teQrZtoVfMEIFr2YFXnKhWoyA46VNvlUq4H1CRgKL15W4laLVoTWMyZo
AqEjKvnBIZ/LjkkgCxUgKbI+nppIHy1LjvUvHoCvi2Rqf8+P12BYwqd7bzV9uoTM
hLOFhJwcT8vubsGXkqNYwIeVZCCSucoHAMnfY8A1NdmUgpRMdLw/8/vZZOLyiOq3
z0FPiv1VTMRAzOnEQKrHzZc5g7t3B2S+ARtNBcExNP1O6WSnUY1EBnNuwOqyNluG
zZNnJdcMUxpPUyvqjv57InHAFRWbJ4TE7lCxIBGJr8mL65hSXJJjdpEHien8EGGL
6cx5UEBMFJJYgpS+DvW8pKIA9NND1H0goqo1/FBhYzSVlU35WIXLTBHYCHFscgSG
aZ0foKQe9NBs7W4arfmxz+F6pLAxjK70Yf2HmcOu1bOxjIRfuqSV14DSBagKsQXZ
qp018AYag4xgoK4Gimb1u2SlYOW4HHiEbD5x3KqOnWMEs4jW+SS/NN+LoU6+hog1
KNvXWJw+KWHZOaHOGytV1fqIIUvhHbLdf5Vf6soo1Z4SFXojLXDFs5pA0gtpfz2i
w1ww0UNbxBCnewRWse5r1pBRvZ5kXytvTCkkBUrlasMT0TIA/+Gj1M+MQgCTm/QG
YC7NpamFhfSJzV6KaDbId3QBGk4RgUBfty7m/gYK3YCAZ+VRaKLstX/iZdbX/YzL
7l9JOhRl1/PcJixw8Eq044NPpOKsEWjBl+akFSBvnKA+ug2hUO9sFCsIOn0RTV3i
ZoRyw1Ddes9Targi6tzvrfCLqS4Mt3+DXgAHjg+xJDC/4HuDfUxuspJesGpJH1y5
L9WqObIFLNnfiKVA4lOqyofRsRV1Zm8XuxA/Rqu8T+5Dks6MJNoddk3VwCjOCclx
3dec8lgi74F8L2M4GtjwpmAANoHbcEWjrulvYmczxJYC2lF9CoIdSRVDGYyWdx/3
5IDffdKy8JjHDBL1sCedejv77yWquRbECfrw+kEWNqkQFpSoblzXwZ9fXT2tTsku
/hMTDwVU3O2NEwuZd7AVfNoN3bKGpy2QI2dTLIY6UWbhh2yYXJ+BX6XteG45YayM
ss/kB8Tcam1PgjtbEYxToaizCPkEp38lJ27feKM0k8xaA+v0O/QJ5t5dqWjGdo7V
KTZZilorqcvYeLrPCkhGVksbzqKc4V7j6V9IDQs8V8u9wgOD9JYbrywJw+kLm1AZ
nKrjz23jh7jx/M3VgD753ZTtLkyhQdlnVss0L5idHepgErxhljg0eg+6inix7vMO
06c5wBiuKXENFK19XJAMjj308fsCnuGWoZgTn5TG9aAAXGuss01QEN1W5ZY2IbS+
GmESlwQR0H50hL8bzuhBvni4UFoTlRev7d80He7okn6OTe8ZZeWAfpZcZgcXUHeB
PdDfbEiayHbl51QbjLSWoGcAy5C+JHm//OWj9sQRVI71spe2pb1tNgVhm0v9G0Dp
DicQY+SS4VikcDiMV7qIGwHTSz1dTK6qlfsketGBAyIiljgYRx53ydc5QUHGZPIA
0KUt72TpebaVYoWy4/cJ61kXr6eNDFYq+/pRBW4Rlt49pnoB0eWvA7qW0U9FpM5W
2e7jSQplnR0WHpZoK+6lmUnZkjR6+YM4C2E+Bi7VMPrwT6IIFVd90y8h7LdNpi6f
+yvyirb2RboUjFM5b7OhZSfuY4JD6qDnb8xl8/pAn8/h8uR0P22xe48e9Bl/GKTz
7Snv1ED9ifUPE/YYSCLCN3cgUA0iNiKHdBYjizn6SzRftK3Gn0UGLPpmpRTbreRV
1lBT2b5d7IGKcJuSYhBruwPWel6H1IDPpikNd31ehqmNHcUTOY59FOVT4JyyUWtg
QdGhDEr5MpXTOJKYIyl8w7ZG0FoXS3wpqYyRWV82/NLZwURu2X8jcKvSAoDfsKnT
GmtTVX9Xs7+YEMXRG1LO37V2jLuh4LH0ZGF7/5+FAeEje6yt0/iFHVxkuvXI7ggU
J1jI5dVKIasGhmdE9N/J1iFujCzvKeTBYOrsoq5tUkiFzkOnu0Z5IpYDJSChSayz
OZZ8bjRHrjwmzM4n7y25b+lQnF9uE8JtoahQtNssWOOY222hZ1vfKVMNW6Bcu0wA
oBwnfLQ2jNF4IZqyL4mKsh2TAnkXP2j8tG0MSh8mAwpAFxUT+EgmHqE7dhPh4EYL
RQtXfs+zL4k9o2ZuGE+r/NdLSeZu72tZeNpyWzxDdRoDXtsR/AKigG5wu0XbatI0
g1g7zME87WXUgZ97lxTmhygIhjNtEZVUat9iva3iCUy9tIubdo5kq3autTnv8We/
tGqUxe7yEXow0ELd+XvFCpzKdwHlbMmNxMHbvOOTG8xcXey/IJQnQBX4JtW+lij9
Q1PDTPnVa+pXo1oDrFMWEETdw0vHx8sbOmKgdLtK15xNjFqz2Aw2Q6IYLc+bjr84
sadeslVpojIGvBv8t5TUKBGxZ3Plas4Ar9W7Vw6UgLRbcsrTLFjo3AsAr+WRdwH3
w48ZYP2NJCaAdOsn9FZ2K9BUEjnb1mwrERj/0U/rPSPe7+RnzeK1mUbFotap9R3F
/4awOvpjR+vj0wB/FiL3REXNbHRFo8Unop9OxIXMpMF4VOxelrcC2XKADg/VNNq8
MfqKYERYjShsaFHPf8feEU5dCuNvdO0870/DwLXGhbOSIQOCtx/S8W6Lrj2EAdAQ
eLFC/fyZDTwgh75hri34j6UAM7SjPkPGftGJEqTJkV7IXFAe8AQuXRMi4sn55Oqb
I0NjaOk/GP1TAtZfKxd+0xQ7OPWto5fZtd1cSUg8G9WUXdgJ3hZ/BhbOQEBbx6dd
tmptfhylGpFQZ0EBTNTKJpVIb1dY5UTJubmpDOaySzBiFudGgJojN8Z5Qq+b0qfZ
i8AWdP/rfAu9R78H4gwe3BAwJF03GlHajpRY2Hhr0nJfSPWeSE4Ovz9rYZqBD/4s
a9OFN4ixIleGXZGOUDZSbQDHAiOSJpJjP2x51uBNwmOGpLvK8PcILNf5oKdbuuOw
LQNbNyHK/gmXLxjn14+d8YzJ/RWGa/uocpFxAl97lgkKOHBryBzDJYeEX8vWnRPJ
IyZr4RLU6xeFlxjjfEFssOvlflKDOWesUAM1NY14FginQkFn/i86cQmUoz3ZoOsd
cc7Qk6Gq63DoS3tjD9yMU+Q5z9ZWhrvxZU7NGaou1ir47XdhQxmHRRLt28Cakk7T
QrKjylOvrpcRu4/xOZfhi+5/sr02Mn+UKrcbwxbXEUmgs55muLi+S8Wpi7+aemOw
gwx30bxMBsvkN+yl2H9prrUlJK6lWZxeWoBzJ2rF078kj7dFOa5qWaN59SfQLnIr
iHo/G80TRqqUhkMe+I4303fnAS7j/Bw+JTR9uP1ML4F9zAXI+fzQyYIePfzxrOnW
rmhj4hUu0ZXHy3meDL1QR4wqjY81gQlMT8og/3UU0EROUMirfq6hgK/7IqZMSu0e
kDqYcY4mzUL7SpNHEDfL2Qk+3R63661CLqWjeHYp2vCBoa+8v9GlXLYilvJSzhw2
y83FyB+PWemxYNoFbMueyenDpm23/URfSoTSxG0GGrClwX6GPF4ekkqC6RpWgQVN
I4jqR8wTGMaUq+mQPYU72EpQEq7Yyhj2/jcU3QKOrBsq7KA06oTa90lQpwPdCmCy
LeLgswXUaORCrIu9WkqQiYpJxU/TRSSkwh+pxSELPa/BH9f7lHoRuPOhWtLxg00d
2jOWVQ1gRYLVhHz+B5iDiEN2PzmIKJcqh58RE3iNTMhArG/mt4IE+dTj8oV+V8h7
chBzgCu3d+6ejfz9OFuxsJhA9AWRXk+U+4DNmOHAG6M8OZue+pryPW7/wpCAX/I0
/IAD1cdpztM5NF57EJwwUDudDIWIKX20Bf+Z1YSA4drLChXORs55/dzmphDr1HeK
v+vx33JJLerH/p/a4I39GsNWfgN7Wgh/SlTTA17dNOjP7efbAz9O8ErlCc2GjeG4
2hcBMuuJ4apStAoCN2ufXhYgEuvksj0FKalhDw1Vzgzas/AJGjoNs5335sSgHF3j
MfGs4PCXhzS0BOM93+Na5ca39ibj3CDxXiX71zbmZjDaQSUHtj7bulULFVwxJbRY
8Ui00kLKxcymd961YekvDeAGahDZERVGhffO7d+LUYwH3at8LqJZVuIwDEWSMGD1
QYvj0D1XsTknK6SkDhztLTOTmu2SrKyy2E0W2lYSFWnCr31CSbpOVLSH07RCmqkT
1I+G3aZEnhSYGtAT8GWa7NwRxBWq8+7RQ7T91oRhaA1svDKmYinjORxI0lRJZ34M
yJ7iYjz9DWp5vzJ13+SIb5U2vbuQ+KzA4jWKCFnuW3STx1+l/EaNT+7MsRAbIUZR
iJZ7OJcwDIBkhs+CF7ibqneCQO2OqrLvkLjrBBSvGFnNLXxQXWnNtp54CxeUKXtn
qTnln1bx73Er32HsR7STzlSdtxh5RFN38kMbv59CCzy3bXYq/yPY9eHXcaoYMTN7
hunHLRn3HDZuaoiUl++dZv+ILamUnrPM+F2hi1GBB3vgda4151ghpmdzn98L/Xbl
GkgOdyhqG1WF1+7L1lc03akaGaDG95slOeYE5V1Ae2mDy8oGgamUBDGnnr+qlPO/
IjbXoQYP8OJAdg/D6X6/NpxevjZlJ0F/KOy4JtquINo03rF6kvq2q/2DAwkH/ZEY
rxh0JHrJQeFObsgFi9A/gmVhefCqmuKHA3sP41Ky44h0olVI51n4/ho2trxMLsW9
0o/aKGNGLNTbP27KOCA6OL/BEpdxe9+ZDAvJdJmMJxeXMNQjmFliU8plkScrdBe3
7amC23TZw5KjkVXNVLRbNE8QBPJNeRZTtwplpIet6GVV/FEhu79nXcdrFPikM1bK
EzlcicGGWq/Fb/CsKO1fghSUx7d1grv9JdtKh3z8bhSMTu18YBGAGXhiHvtQ0NOQ
uQizkYz4Cc7uQVCcBwaXOjtj6WtHirsFlZ0TguSniSxp4FDEkwvNV/yEJ8Q41n/A
+Vk4mrUOXdYlWdM6n4Dd/lu4Z5jLSJe0sZajIgAK4IG01wyE31VKpsuRKs9Bx2lF
rKCquFtvKUmN6Yb8xvqprJctBclVsX9LQYrTmRZKsQV5z711l9/OBAmeNa9uxEN3
Nux8ilQz63wI6wm+ZrIgRaehXuQX0TU79U+N/zyGrKkdFIETzVVT9MoKNPJvZY4E
VOV+rxKGWoCz80w/JI2yspV4hSBzYY4iw+hA1VzyXSrGW+hmZTcm4yMdSEx2wj6l
9sUbUs42R6jl+7AAZoSUf6ZrteEks+4yZ0CYZUYsj/uLhYRLuJieIkzHWtal+rXC
BZTRp9mppD4qFX+1DhzO4Rf/lWkG7VTWwYxiU0hcT6IPHWfZ11MkcOTP8U/ZZRm9
WHnlpn35Y++vVxkL+LrMYQOrH6Nty0Jw7hEnxDVOsk59XPL0K6OgwUwIho83RVr3
rTMUtEWVVMNUDPbugT+HpGiWEVWPSzKo2FmIG48kvuiItTZqCNUDgzmppcYeUe/4
wVixBbum6sTAMdD3sbEoCbGwvAql13jkNiZL05ChN9p2P1EOxJKVzgZKAdvjeTFE
Bi4yZIMaxF+sChu66ia4rEgErTz1e8dVQjpTDSXgSwuFBkoP6Ug6uGFdyDOuFmEf
0qLYGv72shL/eWbugUzRfzGrLScepGu1kBMsa16N6wptQo2yRuOaH2kqhD0BSAL+
J0A4stTn5H5z9axdGUGIuRF2SZby/LYLEDIfR8XHw0GF9jnjh4u/nWOV/Ci6FhoM
qepk/EoDSMWFPBzA2Po+NMJqxUiqNpHOP8OSZ4itnzNyTqd9vqlUpYhnygh/Q/Lr
U4nZaT5ckdq/m4yadGXp/vhpW7a/HiO5DGswDePXbKNvbPeeRDIeq7NSYley57eg
TBQHBZV3K3GMyryKcHI3lOEPO90yc6n4HyNcAeaBWcb+R+fDeRdmca4MjAvMwJS6
lBWMYbVZoFfTWl1v8peTAlsqqBsoILiiGeGVa38z2fsxTtbZkCZCFDXCiuGeAP0n
n/rrQxZ09aY63pYcw3DrKXo92x79JvdlHmB64/qrST2goS44zpVrX0W4JoC1WaNj
kn32fbOJCm2knkq+AT4hZBA7zQSwLHkFzGGMmfx5xDYcE+6PnjgU3uVZZJQ/hwhM
LDVBxAPwvpSqTCYtflFEQjIobcTv1/lLewk5pcXWjSgbjech68byWjoaX2v9quz1
jGwaiC0YIKw0iryftUuULxhDo+fcZ/KHdr5ON/YZcOp4C8Ze1+1NSEsr9jtK5QTZ
Vw2qj1KCwJqzlOGnqmZtmF9oXTP8uduAVGBl9TtywwYPW4OPEY1Zl8i8Lt8vf/+/
Tu08ISbE48xZaKF9Sd+4fQIaNopPzLutxnycbcMDule/lX+cF27Xvt7/E13Davjp
KTSwutWPib8nTMLUfyoCZCwRnEHPNacFRU19rnoM4IG4OkTLMPLUepMDd4XmD/Gy
h2EeiCN5aIn4bV8mIVHnhwAq3XcRvoz1LE7ztIYvy+6FZFkJHrWrIDc9eqHXjw33
gingD1Mo1qtOd22JvZ1cw9Sl04qri5RBiY90Vs/9ZLjgT4eiTLHIvVOTVywAV9sn
DX34Cj7/nkdTJOwn3zsO7tenw5OHVkLK1kZg7r4mfDmbGR12sEVIutGTcI7GJp74
Fr0ZfScgnvkZIf99yob8xLrjQae1u/YCc1zoUmhCc35liR8+xiipMVoaI3kbpzqT
4+KvzbKrXjD2wFDJ9tKEE54vdNlq9ZyRcfrh982E1XBTF9VapRixZzMI3ZAdlv8B
w6OaII+XX2mcvJyN4TTCv0y5B5m2Sb/La8vDW8KDIQ8P6+kJxaq6eZtjQEv7xiJy
KLdmPNEDpyKqOJDAz9OiaHcA5jeWMacaq/Gixe1SD8HzS8ETLvhGSwjhAEMp3IDj
nxIpJSTWe3BDh/bRzBVVgvka/9cl4kLUUkyeXdqPyauw4ELjBxo3EL1joYHYzz76
NSp+SU/WiSa+qaWALkTVQgKMOvDEh7CzL+4pxUG0QSZNDpa2Pxo55jcSSAfjLZrt
+yhM5++ek+iGJZw6BshOYLwKGZUMuie80LFsWzc73DFxsyG+3SJFIlGHg0isrvrh
g0G1JoN0WphvIzaRsXm+LTAYwRKD3D5ammGrUNjHAo2ZR8EWqbEIkH+6Wb9Dj7Zu
AJO4dwRP1la+DFQZdV2UdbyOnyKRrP+j2+NmpF6yOvPnnMyf+hBBx+KJvFjmvzML
2dWaVvppcYQi/vX6AG+J/ePl1KinUghX33bDfEukmzcXaQDoFLcWIwitKhogfKrQ
KG4fQjuObL5OAShPlZLQtiwvOi8j2chyXCqHbewOjDbZjaW9YFMq5+uq/TtDLdU0
JiFp0LqvFD1LwNkqSSeA13mNCRktBsUuhLrDQYWe3+R/eLIzeqS1NDYo9GWOYeYg
7ciC8opb98MxQ53Cazb7KwGFHkBv9c/nQotjxCTvtYw+4dXQrIiPaRTZVYvJ1PMY
fDMxlVOC/KvERCuQyqbYYWJ2oWjJP3OpTUv1OeFubFpl99Kn396qL3hcIA7Cw6e7
J7dwv5xm1Mxb6PDMT65xavc8t0o/OvfhOcb8yp+1RcpgnTIEOFZPSQghSG3TVyNg
VgqBQnQ1ccKhxZERWW+fGJJ4jmm6HITi8x6FAWvTOBnZJfAHu1gB5COOf3Aq1NML
o9hYMJ8t0WZldHp+gdUSaL2cUP5aUMpVd+Nh6vLpjaYk7BATEAuVcoK10zlYuxfW
5t2sxwBwcAvwYz2gBDnjsQZYDK/CVfbW8erOGBryeA/FeU6aLJ8rbfZmedGZvqOR
3WkgZWc/oG0l4uVBbuxvwZGSqVLT7BoCb6ENVRsVD5ua3mDXUD9UB9Vt5kGGy4zL
BkJDOvBWVRp9cdZ1mfbLT7bh8sVo2Fvb3YS4ZF2OmIP48MeIy+5W9jNzImCh2GV3
VMnfPpqB33rtLo4SvxrwseS9mtwrc0CKQjBs7FoVddgVLyj2c21ggws/9iU8tASL
EBcij7xLEqSc11LkXHhgKKwiJ6unqYzTMUcrnszJ475pbu1HzTd4S67MnIQdlJM0
bDz75b4K6eFCzJBnSJFot6RnD2f6dxombcOIv0ZBUyOSRQ7zAfit91XbQmmBp/u9
t/vSEvNbfmPxVj8gh8NiBHqV6t1ajyyzw18gJyPbgWQIPvwX3XQDun+r7DyJEciX
+iVhF2+S/xGCrgfFrFfpDx4JIwscWJUKFoZh5kxkFcU2f/rp8X4QDVTAN8qRumyl
yIdSgoLZhCiBf4yOknfaH1KvmOqlEjzvwfnPfDmRipExcQAAjgHwxQNrvFi/TXQK
O+SWl3pYcdJ6UMujNEhvE0wbXF2ivjLdDeOn0FnaNH1w5h/sh3YBx/MqYpCG5lq4
CLuDmR2uQOxLe9Mr8L3fzlrmM4A5P2u4CSiA2Zskjirmc16e2u3/QK7x0Phs838/
fjfoYPZgzrv0REhXgNLqSALqbYtI4QYkoHxx23I5kni/+6tjwbfqqH5cSu6h3Ptq
qDb0haXWwJ0WCslWZzgDvkHy1fFMzvXhcbXvCuDAl8Q+zoBi6sj8pFAIUtsaPL1q
8jJsEcQt/0oa7lKk+6Na4KU4sA99syVg4hq1sgJ3COhcW/1mDAmwGfbZGaJSHE/3
kPi38Pr4Zo07GTKaWJgU4M3VxBmmIGkdfoW7TFxNAISn5hPLaDgl6w58K9gmgx4h
L2zd5q00XUdBfVZuadWptydMfvc6AzFXZgxxCVS7zTN+ShV4qT3Ux6TM+kUm8QdF
dfmZQI7JT/awibal2XzsoSTwUEK03RWlcroRyCGGUFf/USfNToasrr+RBuiXbG/D
ydLjFZIEfuu5+Bd5upx1WgW/YEpLFX2QPi20IN7P7Af/F4knnnFzH0osyZkcTT87
J/I0WkUHaQbyspg2xfP0M8Ln4HJEyRI0qq8fiuqzLFC9sur8tb0T4DtHICwXz/sb
gcWvPfILs/sKwSj9pL8sk7xIODRk76CTf5msCVYVt/b30gaAWRW1Qh6pY6nMIhLD
jeHEHvP8YCI/SJCFyk+APTpljq5ydamVOiNIaWEOTKUxEP07bynJ/KLGiLdTTu1v
G3tiUWseJDHrP6N9/PeDhgqS25n/+l1NTQDHelOOSKmNshkgak/Ce/Tv9Y9s+LMs
0aFN2bN6k8WmqxsYfDP9N93dneoSyGz/ZR42Ru9rRvg2yUsXUZ9bdE4YbAh5Klg8
/qQmEtMk7zKe9cjNtr9LMXPjrp5d4gXWQ7gM6oASBw/i8vZiQ6Bt9PFuP0gggcV9
kmxLCcU7fAevb46um/Eu6sha4ADGFh9dKGj9Ifj2KcTRdJy5IT6dOx3yIYP0fKBg
vUuQU7GUUUfYlj/u1eO4FHEl0qIj37Tz4HVf6C8JmxZ3unfUGxitlWJ+wILF8A0o
3kwhLLKJJFXctsf7eMVmdEA7ri/q3iSKtr1EeEAKQCANotQlOOn7hvLyJFBiNjUU
LZM79JqVP5lMGTxZd6Nb4YXiLunWW7i9pxolDcSy+VHJFZAZCvijD5q2bFzy6JQl
Lf0LCiFgpKUkD7mLgrRh3iU54VMiL9TvKKH07OpClP9e0UFIsjTIKeKySA7AcH6q
uqMEVLSHs0/tWYA7CcVl2FElLkdhATpfYEIj7blA54BUnoacBOzQkZ+vXcN1n1Oa
uV0yMF7OEDLqX1/sC/l29uz5/rzUprI91/GGvi+I94CZ9jNqxBt0kJnkSoKexibo
EdcDBmIgLEW7px6tBF9rI/D/j7FlFEZOKike0/dwD9yUDnExLnvFP5RaCzCj5azU
NO/C/RtwxH6QvAEls/LGpuY6JVORJyMnVBnitOegcdhhhVFWpHyRRsL0m3/8WMrn
XRibEzgtVqUIVF93lHyTMzgzZwIoHRoKS3akxavTC8yGiUXivxSj5fyJpiQix4Ez
564q5m1aapyW4YQ5fICDvUsXIzllbhDAZp5ciuaJZ2XcixT4rote822tEb9xQL8X
ELG3lXQEpogEKCyRMBsUdFvf+4y4D7a2cNRPTQDOUf43p0fDnQ/ciUr8/Za1mwJL
KDhkonJaaaxZB1FbCNoKSkUORh6BWZ5Sd53olrgZOicAZW2rj3NzbBvWQL0bIdAt
EpguFISyHRIPa72i4SLjhYRTdeJAWzd48U67HJ2IHO/a0UX+fTXpFWAtsBqzCipi
UiBEtg+wtcm/b0WPepNIZN8jAD8/QtZvnLe2qex4RNjOj5QYCYXZO23pS7ZGidiy
YlJbVm5Be/o58/B2yQlz6r+7LwC1GfHx5NHaRH2L3ZWpcE777YNMrkpo7a6JLKVj
YQ/1uSroNXhuCuaDJ2Q4FtR63y1XPBzNPWQJ+ZekUnE5F0VPLCCMOXu8BSStxBcw
0U6eOsUyaY+dHJAeaTB+Q752iwyfgMnhCSHOyKHgoNY2gwUOJcaKpxiyt3dgIVVU
Yev3MOK3jTWl4LZjM7eYmSfb8la75zhIFo0o8gJronKqoDKgI3w8ZsJKqkgG7BIx
6uIUPJzbfStkaUp+RhHVTZuJl9wnYPB4/f7YVjrmnpcCgix5yq8/rBgffCgemFw/
tUBO2d6rBqfXD771Ar8n3iGBT8TXNIEMsW8oOEu3I/3vjAk41+iFkqtxYQ4xCQh5
FULu9drqQ49ClFPrt1hU02jb5tR9OE0MGNb0Vjcj5m0xEWBLnkx0UXtEYWqP4zAq
Bmq0CKBcA/pheS2MtsrH3rwSUUMv9c8t5TFe+hSjiXnftu04ql6mafa4lt2VhgiT
MvhsQI5NPhwP4ST9qwvFJz1HMkTQJkuzRgD2PFeQpK3W4dhIR47OUjrs7oA4JA4r
yl1X4dvRcOhgcm6gVLIbE5WEZrYTRmEF/7tmgwk8pwnLgYPw7HabjS/AtNdC7706
S/RbaCczvnoT2lKaKiZYeb9CEKfNIxAe1gjp4G9BRsBnjLecMr7cg6+pZSnZ3n8/
i+Wdn8dKi0lNane4ibKmT+aizgGC0TrdsW4k/wLu8sT48X9eavOaFDcic8ikRTrA
bIX7YfDh+JyxuHM64I5PxWmec10YoDl+iNvuyN8QLUWRvlFVxfW+7ua8CunAp5rk
3gcGG5hCVrdZRItCl9xDOk2BScZ89xqTOzaDOTQU5UcqIaojlXTa9GKeU7nytvWB
Ms/FxaHFfDAktozspeXxNitcrUTHz6UOUGA1aE7HQbWPtwghrj2fvB0OuConCoPU
SXK91tdJV0Or6AgmVhHQTEr0w5kf6hMNavbvtJsq3Zp5V+DL6Q3pYt5C4tnzSTG6
/lP/LFb6rouQFKEYUECydnzuXemJ+wyBC3KF5URR3ofxfL1trvP+MIVJKzn111+g
OSl0oN2Q2e6C8fQe5E8QYT3+rIjGW7CchkiOrfJ9ZW1be4n6dYO0SpHASYN/RKoc
VRWAd1lyqF6Ncyr0JmULv6gWYbrJ5GG5H/o1l9f4ueKXAdFeGGM3V78po4rf4cPi
4ySRMQ6UaSozw+7pjWCkbXewA6JAYT/S+GhYL58q+jW1jBCVusf7HTsnPfoxQsMo
APBPtBG8iWOymloPfYcWA6rgQ19/ZqDl/T1mpr6Qvswzku9oGvZX1qUl0oZ0pVaz
h8UL3i9UOqJaI4iU6m4/SaUitcxkW1sa4Tt2fJy+b1oPA5tbqJXLIeXTbX6EUhPO
M3R4ZKwjmw0PFgURoc4OI8pOn+lfMYZTKAx8e8yoxH2f/ae6eCW5Rdr2DVArhic9
6Sa40mcGqgVWS0dTbCgGGrCpb+piD37xXmSNyFNdSM/Dk0Py64Wd5CsGJgezSJDt
isZHaiE5j2KJSnuZWDa5LPcp054anLpxR4QP3bwLbFoylvYtftwEG2KHJDxnAJca
UvTkuNuvcc8p1mgoBys9iVfDlYEXA3Wgspd55Wr5mPNvnptSSpKCZfVUeqv9RAvX
Dgy2FOxC17DDC0pE4TQMWiD0nPFUh2dU6KyfB832Jc17JAZgOdy8OYlQYHS/bmYM
v4I0ssXK3hUvl7oxdU9qBZn/hFnQBj5sQWviv3a2GzIMxmHmsOpC0rl30yxOLtVB
94NEpLZRV7maY/9vjiGvPaNimTiY7nGpzyZqwTn2XQDi36G8dp1DdQm5P/1v8+Tc
hdJvwTAUr3M51OF7t64fRIYxDIviJI/27fAborSaqUODHgcV3jb4c/trOqXTkfJx
fFTE7q/7P3pVsr8/gRrNordzg7+UClVWheHbiEJSf/GxhCHY8KVUlbl6MWwIiK/A
v+wyVTZLz+dyWLnd0MNIva1MlUTAx1r1crmS6RKvdypeYy5DqMtSmEgLXx4Dg2tU
P7zDs8Ku4YztgUf//z1NKBinjRfpIxl8McBzKv4Nmq9mhbgmCIjNI0yjz4h9sEss
tlYfxFrrgjikNVv4jlpmXDyCJXe+hZHYJVetvBHa9KSuCpQCcwX4j0ChE83kGDza
uty0ECCx4orj+AUNZfpQ5kyrK9XkXnsllSteR3q/3xIgCj413akOAp0ddqXgeXX8
OgnflVQS1+w+enJxeh00vgwq8ewxrpSd29mfHdGU4nIgWVeOkIcJ1C/hqyrKxy6Z
i+R6DCJuxT952WsTcVq0JmH5FjKwzwpB+BYnajmKD9BF0J2IUbFQiX8JBM9YXvWa
fG7JALaEsxNzvWZCamKtJxg3+ss+yA61epJIgSY0Q6vTSN8lAX1rv47Yy8KMMz9J
Zg6jKcXVh0NiRbWM7y5U9o09YtWI30Vf4LO81Z82cXX43R0bzvn3emPMyLQGViKs
5gbwdb2OO5mMkQlWQ+rXStv5i5B6qIqSkkuQScrq8qdQ7FtHrEj1EvFYxBE2yYkY
vAmZD6lIrVI4WESv81ZlXacDzVBV3VhXCWLJxvLJ9aLXXIy1ahM26nJ7wqU7P18O
yFqT1nPxQH4T3jWWd3rRp5ItJPd4+aNwvUYHy1lbATtIddJBid+b79QV2qatueFX
DImUytEV5UZxUMmfwV7YKgrFWgNpxIrLZ9IwBTI8Pl0vjng2bmOyO8zEXW6jtRZB
KMuYMEfjd4YzHuIZLVxjKY3FX+TBeAnIC+jiCXx3+16SinCqsHhWc8kgtZSEKvwn
+JaDPYpszprljfHz6GIenLRrM9wsSWinKW0GkkhPIX6DH6QS4DPYF7e1r41HVOYP
CZLNgOI5Lw5M9wXj8jp4/T30ldfLWjFXWpbq6jLsnXiZEajIRcLp5us2IZjMdTjX
pZcNbf0m3x/J6l1o0Q+5hPWfdpQxGCXF4GUYd3+D6AdW5EILRZ8s7JnPoQd5bo45
K4vSVYYKqwtCvUdZNJw4uW54k7t3fZshWLC0sIVv9En20EK/GyrXuiLeKQVkw/Z7
sQVbYdeqdVwO6oj1G+T40sKJ9PN50mLwzw8f1ZS/7tVztXmMefT8dLQHUdT4Naos
Ztt6oysUEfgt4u+UXOwQTWj165beMJXaBQZYAFSsIoPOxAtEdtJYrqa1Q8fdocSo
nKN6jxHqDWp75W6LocvhASkrIDPWXOz6nBlQXbOSbPjc7K56KfLvMZLjm3hza+MS
BHVVnyFVTo0KDKnVuSs3PGoxLjgxkJ7Q2ys4JzWnBuH5O4s/ORD+nq8WewYasHho
BhKXJTwWrnwdtnCWVRNwVuT18+moqss5vSWSCyOmdMnLmJjlWfJPJsPkkWlAqz0K
d9i7SSmDqqtLNlAKLJlKIVIVQ9v+RMNPAT0iaRZs2Zg7IwU7yDV2jF6/1QdyjtiA
QMs98WGCdnuLbs/x3cU+5hhOjFsBd+t208kYvhgV9hFg3Fgr5fTfy/o6OWadnby3
RgheecdhtplFZOmTKIsnUJIXOUTaRPZ2Ffwl+/nMAOF17+s1Atmlig63bltbQwDi
FUxNr3N1tzpDUPhTRZh9izI45fCEGAgu3zsHjxa20K6wRcIDOmyHf+iZnngO76jg
RVAAPHSekOvmKiK3y+KlVgsBEM8kBRHTF3qlvQyz69OuCjmUgRv2Q0cHLgjsnTLY
aYPrtlD1u8aMKea8fCjA02BUIQel0fxSVua3ooIIh1xWtiTBCAmLSDZBT21OJ457
r1dxFzg/Dt56DHcXKih52p/0/PPjdHjXbKIwE02JTdK/iS3Vetf6Y/n1uuGuqAze
OQVRjZT+pdi19uhYmHt24hC8KEuQkFsoRRAIiDy5Viij3M2wVRTRbYhOYY+qLsdP
Mm5VfwCUbrBKLUngoaJ2xFQv+kOkioiQ3WST9+D50pGcEXiLxPv3qsinOCPUzdmW
h9Vor2OCfhenvc4WmEPK62W0inCAgyhqkITRtRlHTWE56QSkzJxMspmhaNdRPJJo
jdDu5+h8fu+0q9ZcAQXFi1ajEbNiuVn+l/mSTTG11euBupR/WEoGeDK9MywWMkeh
CVqcFAWutgpN7f3wP22LCjtb1CgSOgbdpOCojNPq/Q+oTIos7wwrFMmoul9HZaRH
TDsmQgyFiUmVLBrzrCtkBs9wrbd6aT69W7kZAn1p7MWhFdwi51QmgD+yUYWL6NpM
NNeAIJMdbReMkRxw0KoSi66ySGSQotlpfIySnVosf89T97sV6u4obhO4Jty6dr7g
xbB0F78uoxhfrvCMDPgQMSa9dqMSL5A503vSIBdj/ycR9Aq/uxUG9kdvIEhHlJZr
Ooj4GOKUN4VVkiKA4SbmiRPrLblUw28DScqDBGgkVp+u/l5f4OrW3tLoSDC2ozif
VZqpLYfDtV5d9khy0DeVMXWu1YJqkN0xlRf1A55as91HwjIxkwCPYlQtcqhPb3nT
GDHUQ1lmiFsOPDEcUhJ2pN7Fkq3t+vTk1uNaPpijFsHVOHM4FbSp21IvrZbw2v+2
WPPi7J0unWLwT6+disSfLoiEJBlz8//6zjREgJ/cUWt+JK20gUjPE2ZZFfsn87Jn
+41sVJIBtgLRG1m1U8vycZn5UiD6J08GlSJxB5G8xvxw8/0wNmJv0btGwOSxIYYy
ghJ01aUI6pj02/RISciQWp9sYBwNERQrCoZB9yRRuYG0RJMxTzprM4jCM5RoXDyD
kn07LaSFR46WZi8yJgi/Km1J2Vk3DDNXXu+eMCDI4WKR2Gj3HQr64+3KU/sIIIWD
lhDt6ZLLFyN1UuzW2P1ylCDLihxDf8NBMCpAXXiptNP2nWmuXOCqHDxjtx1/MLwk
W9M1EJXgEJOxBNrRIlgNfH6kM8gRt/DUk1z+iGpRE/LAY7vwrPv3IzTf/LGRXwDW
gWy1yQ+F/3Wqg/yF+UzfHLF1ofxr2uyq+ArPqIHaBWqjkmPCpPczycgB+eun/BDQ
rg6LQm7O45CK+HlHyXCg6647rfGkFAkP3fsRWkJm/bYdB6EuWKKBaHKyNzpxAhPO
f8nfXs7st0NGHKDhkDHPR+FaeNer8f6rWnjnRXErvRhDKJv6QtfXnQ3T8UNRCuk3
M9ZbgwoxYaytVY/WJ3cuCFlmNMIOmX8ezDY0cMr+sLw6ClMdlFbeuOgUI3l31Q9l
FKt8mqtlhAOg0nMZg6REAwTneMxUbfqJ2E1040uJ3utJ41UqTl3NF6fkasAErSzm
6wH7nbRdiTuWCaTGeax3qm4dkpGB44ag1O/RkM9UFlkpC3Nbh9aN4Hixf910rsyx
UpH4TS65YG+EKn1rT3epbbIFL7L5PRFKYRiWt896xs56acW+N/K4zrkTShNaMfb0
XbrIDvs4K9Ef3CjjNtsBT8IEjQ66Bn7ol8b1OXE1hFva6LuCvKORAG0VJcCicXGg
LVwfgqYHwytwOKr+3lwprW7FIbJtbH0sXnQRQrdKNiANrm18tAhGHVHFq2BfPkya
LBWUnqOwInsPLh/zNIlJAPlzjcqpp1zeU6RcYRYJI+8ToCQtsT1kGYnfDCV9v/lN
K4Un5E6tNb/W9yV+Sxshy8JsKV68Pgb4PZV/DlfOL0PWXAZ/H3RYodb/tx/QVpXi
qjCh9fX7e0Fm4yQwFSOUXbqmr1aAwndHVv1IZ9G+9mwXmcWdtGaf/pJaW/88EmEm
BXT1u9YOhlEJZKbQG/EHEwxKZCrNoMOxlXhgrD0iXz6Bu2gKwtE64mLL1I/hh2yx
CwduszzjCZVzMZW3QSbBDcX2Hgks2kcIlHbhVI7qjxJZZ2DsIb+X5/XinsTPWH0O
QUPYnSDEduLSAwV+eb4H8h90TZVVdkrCMy1nINIdEIDWVl+uyV+sx8dKkw7jdOJ5
OLAV3h4ZVq1r5hPwfOxWnedeAZ4kMhYLWGD5IatAOMAOG5nlBxNV+bk9U0sz9J/v
YAUAUqnJBjHymOK+2MtYjxvhRkB80SQC0sKdkBug4++aS5zD5fCr3r6H3QY3CV5Y
J5q9NhzScieYnlKEghXQso6tV3f7ShRAhZwkXfSml4TzdH+X3+qCHjJGvbU2MZYX
Gh2Nc+xwGnq4J9h33n8gjv8Q6L5Az9JVCYTyOL4Nlp3ZmC7sChoVkYrLC4+I1y0y
MU8znO7ulknm8Y522Dy1UStTRPgERG7a2Kg509MTumUkbC2gFF2MflaCqriUt6hF
0tBvunBzZyVX3McE2Py7dkiq9SEkxk3V5lF6TJ87FHS6FU/OfqfRh7pxCZcjOoOK
+Qq2OmRfZQUiKVoOUDc1SGed7/VNTmd2foDPHn7m9FBpQvruVM/3KYs5GUwji3F/
BPcd7jqHEJ3K/UwGHOTHozGXzmyDf1bPWvevt+2qd8piq8imFZp/l6p4U37WuGwH
yuvUMX2bRMalwGlRlSj/I1mZn8KBNX5xEzXaGa5MGj/crzqpTqlYPmU500lpcp4C
+IT9sZeWjjHvpXf7OzD+QMeixEgXFxInB28ZLw0aLN/PgZgxeqzLgfFBDYSTg5Li
m2hNz4XEiOG3sUHYiZh8wiXFNfcBcmaKkU3KyOy0K8wi4Xng5CrGmBLgILS6au6P
lRUaeVVv6dC5Ov8wyW/u+Z2Vy8Q1L3Sz0zXKh0GaffFUI/H8ddT7MV/wrCsDKCT9
7AUWiduLp0PmGWUQnANDSZkBVtreXzIy0LiUZpG9l9p4CDawUf+zREOt5/r2PL5u
ZwgBZwrgsb9SynRWPWtuFMggCkUIHz4kcKNvx+EOT4GwKw4TuM60Az40GoIPvwSA
3Fnr/Ou8KZTCrCiPj3t+GqZFLREtix0ZyRvEvUtU5/1cshsAAEmFiorL1xPyCPEG
RxOTsajPGzq2BFTwt1kANqoFBrMRqy3bXg6pPW9xGUmqyCOtDNYOY7FBCSHDw8tY
RMjAo8w63ysGBiZw79HUsThvyAEk78mxi6k52v1wxJZaQZn1NA1ovlDzOSgeUOvH
uzjvs37o7/o4FMWFgd/tUONuhiQ9aL2ONIAQRMzwECGA3uhNSfFqInImQC365++c
PXZpgLSZcmGHgUJxu+Vgby5pBJ4A5jVXUP6ojbA17qURNns0tso1d8q5C5orPHP6
nYeoEEpG4QBRIsKC4Wc6F6MDX+OodQQ1kD4E0unRxfV4TXKFhtRNaxIzzpTbC9nZ
OScas2BSxsobmeSxEWIhEPzTeVmmztpLfSIF1ZPCuKmN0bz8fwL1vc71PQtJ8zOp
tLCppj4r/hnavdUQy9gYV7wUfi3zCTD5WAcnvrmE57CVUNdOiPlMUBtXA3xuCwEh
aEUWmfi6gdYa80vWKikoGu8XRQahZr3XK5Drz34pAELLnuWE+kMadPYJkLIr64R3
rJrM6R9KZHUGXnjV2GwGZ4oPW9FXwiE1D6Mt3tbumo86ClMtm9+1qJLHeQq8UNmc
5fNR1XTnLJ6PuBDaLLWpiFOguh3hGwDZ7k2YitZJCiuo1ElOyagBbAUSpuN0V/dJ
yc959WDlXas7TDzsA0jzetRCubn7ddZyOWDM6fWTjtQDPd0nW1eK+fsA3UfSDt9m
srRp/d6N+fA6nwNjIrjBa8AGYPlg5paA9YwUl9cUWQq5yHOp/GBS778g3FVaDe3/
xHT6F0p3pSdqED9M34fj+ODjiNgTJ01Rc1b34UzrIT1LljeOo0YmUj+zE9CWh/k0
ydpdPf+aRkE3lFABCoLJdUdlWeU/lPk3TOd0W2/9xjd1EKd6nLQObE8eKvwcvvUi
JnrB1BwTzJtA9ICOKFPIvegnQKRU6cmQilfdrTJSerMrUt0R2eVR3GVwK/XYsC1m
ZbU47EaFhg22tHknUtavBM1Hw6Tcdz3n7JnugYle/mDHyU1HkL9Ur08RhjHcZwFN
w48pp0xYUIFhsi64aM5iCaFQ/+ql/cO3QrkLgMMe6Togg4ut/P8rPzgvYWrhnNHo
IwIoS0/RB3eE65Sr1aHIOJbL2ZBFpuMeafPROm2HHXlIxjsUELyZKdf6ozaIwBYo
4wCy7y2ZN73Lq779bRdBFGtsKh9FSK2KVJsUakgj6khaWnYAb+0e1EAIL8qK0Yse
X8i3xELlCUqyhGWN/Q24HuryexQ3h9gwZYW0APOJ6SjnEnuZxIStnIo630YGciu4
Winv6b2JcrnaSH9hC7ZbLpEkUJ4b1/GRxImTCY5u7183YnzsdDRDap5YLVSMHXsY
vIJHcu1PQrDoS/0t6KDO02cUm4McQFpzbJKZlMS3CG+Uaigc2X6HW8gARPMdBXfj
FXAsm3d9Ifzgjq76osBBkck19Ka+muVflFGDQbICBuLSzM/K+AqZw7JNF/AfUya5
pxg6x2R7T4CNpnpJ8Zn/3S11qkQnAAoGeh6nZtpuYl73j/fQEyVTczY9zN95Obdf
nJa4JBDm/MwbH+lrvjdIU6I1Nhl8WSf953KChG8v7vJ9I2c2vTljshFmqRJTS0I5
jxxUV2seU1XV/tzKaLPJQ9ipjyvqmHU2ZBOYg+YWfk9aApYqcZcDoPtWdWnGJ1rH
3Vlv+d7bumQOxOwERoy2He65PTQi+VjlByHN+b80uSKWmHqtqV+sIHoiJy3DSu60
PQMuCgcBzQGZfnsozfMvyO+HrbO139kKHHeV9/PvtQBp/64BLcCKaKYHjm8f82j/
Y6Xoig2uDLDX7JpZ3sbU5dbEAxEmeNIYCAAO/G815+4S15zguVkTVtm2J7y/mOgM
KMIh13ySXt9wfyiqeKhT0Yv9Q11fBUp2f4ov6KBBuM7GM0mGx4CUMLHAn+uaJLMb
KF14iYpDKPkzswOzAMxvPhtJE7IJTNrkjgZppddXuOLgDlpw44D+5xKBTCihW84b
8elxfNpNC99U549XiKZPODAw2HDtDKGPKvf63rz9c7CrXoauSriIfWYgVlmhVSEl
5VjkhowHgxW8y1YIc1JtQLjWhYqUJXXFjWQl0h57wBcmJDaqmI52DpyP40uJNlSv
3nNcNO94pSXNxeZfc/x3qgHzEoph+VxfbBZpBnGq0YffiSHiv6W7SCUYV14GIFAr
o7oN8P5sYMNA348S55AJ094lk99Q0qzpbHROszY7MsGCI9QTC4ko0Qlf3x45AvQD
Xk3bRt/yO8oBWNwPfa9JodmY9ufCeXoqCKmzIOD75BPGqoJo+8Dr5OS77OMGVA6v
TB6NcLoiiU/YweYeFWrWcLO1e01WBW94BmHQZhT0YyTNMtt0GWR1dsrIkHSEzsP5
hrSnws75KR5z3fRQochyCm0YW3mY/R+I7qdOkcXW1nJ+O0/QVNHhMirulwnCr2eP
o5t6+3UMwsP6zgedhR2ofxLeemxkpn/WHMITJogDOlM8xY/7Kwsn4qG4ye/VeAC9
F00BT7M4A29OvmpqZ16dv4eUT3zHqMkGXQv93eSEeUukTJrg4XzLXFQSEc6L2ouU
H2aC/fyHe9mVrTytomdic9lc+R/QrciR7GAFIpNbuaqGCt+Qe8HbLkQNSIKi1d22
wfD7joDjKfBjoigArrd0n6AvK0vFkxTh43K1aQ+3jT71kTGa4mllFmSm3aHl6lcs
avy06rqw1mJfcp2FAf2bhJuH2vM95NauKgxs3E0m8a7UFbJAprGen+BXCLFL0gU0
dMMoVJhjyuyQbPlFA4m80UuJ62QifCkgR9C4R+EJrIF4JkbBJiY7L0tZ0T8tFh9y
Q8bvBw0xmuAKQHZUnTsxX4tTQ7aHBLZiXAK+iMctZfcG9Nef4QuublmE1vvjtKuh
fHjeKcTEo+fwvXFAKPNnyyiCY9mlnZomQIUEdM328eD1xzqIjD3CJGTMB0GYMI5m
QU02Mw6gfgcXRRsBmORpE7rQMS7DDQlwWx6jXDtIYbSVBRupPxQcmDHzsy/2X8O0
WNpvW8j2b2ypmNyowqAIm4JXgUZ4tptlp371kX74nuJs5by0C3C+VBky2UGkASxs
7b0P/ZJZzjHk4FS+YUD8uMYFD7dP+nxVOxY3fksnoCEi0pSQmumnxw2d2NfVXuGX
boLR9ulJDzOf9hv66+RcL2WbTPuTJksGIlSLrskqk4HFoNO4GoZG2Av3yhJlus0I
Cmmpo5ePoI/hqn49a8CI4lB4P7KLbU5zcIdUFT3vfBS2McTW53ZAbW9418StkDI+
IM527coHVI5U0gWU6SS5sDW5aLB2x5AaQ0yrHHK4ZLu7ZqjF5bFiYoPApPpxA4Re
Z2iu4hfqkJ/LyqyWC0TWu1ZmzQKlbj2rnJ2eGq1+FB2bRY+UseGkWj2abN+ih3ta
4+CILBhXUaSZcV/5/eKlo/Y1s+K5Dmatt6+IeM4SeGGrxn+okW+5oF2PWoeurfnS
aXQKNwM2+U2REShyy12Gc9TpdwpSYETIRlBhx/0BNw3cwcqqCyb+94hy/r3IqFTG
0Og+UZ3QfZfxhZmXpkIHlWkg1fpyPndbocpbVXxpH/wmJXdbaPffCPFm/mumV1F7
vJwroSpwjUOm7NjeT8Uy+UJknVV255X6ulYy9/3d9I3fWR/fqhv0ckk746WZfLGX
y7c9d38gSP8NzRAb2tcefvuUn7UN8xAOYu9HgGh+N3opl8FhDhLkE4n58X7X9imG
XFF8TjkWAEkys4qi0Wxi3NbmT/qRhYMmuCnk9BLStXJAJOse3NYlIcJ4OdFUl5BU
1V+p6/sZNmw/nWH5WpI/EfD9Ir5+6iwK3av+IdhOjnAov3Tepn6T6UkJ14IEqBtn
ESfva932ct2fLGM0+jVepjV8wJzZBSjqTFWz/MSWdFqasdLuPWEx0B3QBQ8WSEjN
LgNA4vKHNzdaLYIJn8uqgo5e4SlYaN6vtoiKpP93Yx+nNYhce9Vh9hE161vOW2aS
36m69xvE7phhaX90UaocMw3hZ/C21CC6SoVNIv9BkM33eDmV1NXT13uKhTb6nIXf
Yyq7jLqWbTRN2ikJURxatOg+kCAkrIRxFudMIPioZmsFBt5zMNnBUpmW4NsK/3S2
uQ3eXq09YWaKQ5Q6jeQkIl3iiV0WqRH0SRQkuKuCsemxlpgYFZb2UKR0Mlum/4KQ
hQ7KHrfozfkdfaVJjkg3PXr/ZVdG7xt/LP1xINZZm9xFGHJ66hsl0YsWZrz6VI99
AKhtWenV8aNNHSYfUWOSbQy98x2fAjYlTp+r8+7m93w32aMp0sVYG12SEg3k9QZf
y4If1M8IBoL52AWvR6axYfS7JOaSWEbxnvuT/alOuN/T8zgsNtCjGLucQKOyXitM
7+7u9bGuieQCswl3UtijuB5E0PWOllf4LjXgMoPMAcdho9tOcmBpH+j/Cb0TBYtC
Nys5DoBAqOlhzevZ2Ju6eayJ3TLi8M4yX5PyWQF3aIJOPjG9AvV8cfiwR9+QfPZr
RWvOsaqJDLWqePpmK/r5QuraJTBlQwcpFb4Fb2rNj+u4cApic1rrC3J6HGEjOBCW
EWjKRwBaRDu4Zu3P4Y0qBhvptf4OtMlaSQM4GJQkYheSeYT6sZel6hIa/zlLhWJd
h+Tp4abpqeWl7c5eenCt1N25LakFs0dB89VikTVIjULWSik31DPcDUoZw2et+0OA
K0ukUJQhthW7sk3LO0h32yPGr+4Wl3xlvP9ddIowdVelnOiFgYgZd1UNvwlPnBVt
CrJNbJ1z0ufVgkwapRaTzDU7Z/nuliBUK4TmN3gJIa0lQZ7E/PI8QkUuk1hYEZiB
uAoRZQbLu6QJkYInkagIxPkaItZEd5Y9SpimKtdlf8Ksml2k4oyEVUsURyZm4EMP
DZJJ8tPMM98cIpGhpN7sR9oXgWQVhNdGQwbqmCc2YuM4cnSv46je2CVypygnjh6q
pceOSxdKb9jy0YIkV4Zw80TMqAH4LDnbx07Qc0o3jMFuod99FqOsEAQwVnbyXgLX
NXMt0IA5/a3y6lWM/SNlzNYM+b2WEtD6SULeo+Gh/DEmy23FWa6VmpeFal6uYXrC
Ceq/PY2nVBbgSekjnWR8CGkiqTTcTuf2L7+HODaO8G19i5G7NLXaZRnTeKP+t2dq
X2XhYJe0u6RuOog1+JfRZjIVhwvuBB9Kl8EeCoZPWE9Y6egf+N9j19OTEA8Z2nke
2lltAwsW7OnuseJuhPMotDd+HWmsVeUclEdb0Yl3UE49hzyvBuW49gVf/hI5yG1T
Bx7vJpMvJudDv4uhD5YI2eAO46ccWnChmA4gZgaq0N8Xj0/Ws0HdwapNTLqykO/6
LzPRFUuJMGgrpq75zswFpsf0WR1/ELz21u5vRtKmvwAja/AU/809E4mNGhFXevsJ
0hoF3QhV9zbOe/vWe8fvgbdoWZv1Hh2ldQYnXU8ZQP9nr3sVGWLjDqy9SKJFYfhw
jaJgfccuK8fqPams460DR35Yci+yjprS9YG+44fJvWIm5leYKLtyuHggWZx/3qzR
PvvMxH7hiiueqSZ60//WZVSQ+j52CstWMGFgoXFjq6InLFigqMm2kKqRxfDi0u9w
6WS3UKwQiDpTfLw8eyF264UNKL1lkw7VQUAwP3R/1k71yH5DdiabEWLoh3NdJbIk
akPu7SwknSRFVPq0fKjOm1riQID2JVl6xy31aHHlmpVbNy5GPdIH0i5LVQUZcbin
Ev/4+9oY8u6D6c7nLMvsE0fD0Z0HKUMVFID4D98MYTENEkDEi4znJ3tvF82nleUZ
BFdi5BpFRACAGiv6SUrCIlI3PfCtkhcgG9HwUhVtsBujDFFJSRrhtFhoRQFjWfY4
6Rz7NFgtBCjHhka0a2ZsCTpGqvRMoH3dOI+qF2NcBARNaB1TGwvJYB7jyAyMBrlj
TrKyG8cGvkaRG6C16MinmBQcqWtH5BKRq0G3Qx778Y4s9bbw+jKzehP/IkmVEI7k
galUTXIsTOM0myUrGtPhOdBestD8PJBuiR2U5xw7QH+npdCJM2M6ZX5jadu2bvs2
Nw1hmyvTHQEIh1FGlcqnNw6h4Ex+0BNMKmsssC7wXefu0yJunrmd40lvGduaKVx1
Y0vFvz8zI356uwI0DV6VodgOXmAdgUHLbpeaT2QBGEvRtLFr1s2avKkNrwy7M1QS
HrVDHhJZ9GvcXbaimjPXIWgA0yszNEU78R4JTq6UcMXBmjLbAJTil+DK9P9ltYAI
SDHhJWIjhkglPrKhnEMvgLl7sVOU//sbL3eTP+7Ut/72JH99S2Js1BOQ8KiqyHjK
eSB2JjIwqlyOAEdaPqYQFVJxvjfqZvlx+hBCrXoUpI7wOzBiTqoWHhdMnHs6sBTU
rTfmo7zKpgw0RRiCDm0r/pII+FoXaZH/PHsIvR3tW9KPynacINsjjhRpebQu371c
oF//4nqgCpdgkABRSpHmqLBBRhKwAbbKaT2mblfT2xzcWGWwboK5s+4KYuhCoOtr
7Fid54voh/eC+rAzFQlTcb2KLEHY39rYqA9fvkqOuEPJnE0z5Y9axXE5nbhwrTDQ
pJIJAtsvFgYGV0nW6/b4TVm/UvtD7mr3p6/xwD92kaaD5lbkbZvsNLg6y18JKn/5
FelsTtOBfvxbPx8PfxyoyfYUTKAZe7RkjbAh3gULnzwDmUdUXYceCXjJ9QWwldbL
LOqEQNuN5e160oDHV9zzBB28lsX7nRBD6reckUO/k2RYJzds6oPNmf5YKreuFdNt
F4WpDXMcBHGhlktEaVasyfGagP89P0dTUSQyN+tCwIhy10K1heMMtdcysQufU7uV
kKj2nKFRQjTOQ6hNYYC4jXw1YhPGqoSkgudqzM6CJ3zBKSSOE2nW81P/+K9eqLJZ
Vpe4YMW1ZfpJoiEdk3AZlC5nwNPRG4QOELkpLW4D8oG2Wh6QPECiAuRKTa+59HJG
AAf7AR+JXe4y7XNJ/raiVzERu7VFmMnBf8h16AXChsGvrt47KLTxgqLo84IdU5rA
MoXWboH4tvDHxPFiXnA65mtXS3AhrRz3Pc1P4l2MSFHluudOwy3uGYFwrmoR6DYE
sbds/5mvEGweC/NkADIZFSprQrcYbS7DnJK5jNuO1sb7WIHb58Mwil8zeMTxuS0q
2lmV3toiyxwO4o47Kj2j4eu8lAVrLUAyPGKSD8t19MZk1SH3sFcM5yHeg6eO1KFv
LVkieVrdaDucOfu4WZwaMCV2uuac7eU++KvP0Utf/NBxdMbKz0T3iKfWVRqEQyMu
ls6Lo4wozVdmGY8Caw5Q09niUU01Ku6izFeJRGPA/V9fLZQccB4kJbVkT8hzVZjq
v2To7TWr6K2O7kgxenjz0TRmhMuMNImMVVLSyviccZIhCvnAX88+gYu1o8QMLRaf
jumlizUhcjHdIzx+ZHfCvMLt/k3P3jxBL4czqe75TABb7nAoQvXh7X05De9IBX5m
EDKhhD5IcTx9hdBSC1NOqagSbPge8lsh+I/71jWqZT0sqh+1AV1xT0P0GVjAveYW
uqnpy+O3q7bvKiD897Wnq+a+aZ7PA9bqvrVmNVQgvAAxKzhllVf6/mtQOgZqwqCP
pSRib71nV2t/dbAqY2ACIvDpMk84Pp6w5s1MmAl4k3tEOw+0K1KVnFQt67dkarv1
X9hu+PwgzG3WBGJIcMhUxXek7tmCE3AV5yI6dq+rCH6tqmLhLPSqr4l/BNvdiEds
DovY8tIK5F6we3cCFajRkZ3pWqsCHPpFu5+fxxCJLH0NihFJSleCT8Z66R+HB85h
nSxGZtZ4CDFd6lUyDM4J0eNoJIjssySHVi6kcgc58JnFiIOQ56dcQbT2ixCQoT3g
IfGBEzpi0c6/rdPXHshp86SlCSJSNWH6SJSX8FI0snFjRcuCry5oXL2tkihOX7ix
yC+DnbhrvDpMX3g2ySexvocqfOwLMuPb3Kd0qudD4lMUUlfKJUDZShvgL4/t0TgC
eI8/XoQUcqSaZGRXjlMVHF2YCoB/2VU9mPIT5ypApsVgIpiezaIVpSDv7+eYdFQn
XKZWZSzceUfEsyNm0HshjFo4z83iL8/Y1vvN/TfQ9Vz5C0Ota1GX68UzOvc8cDwm
5yLrvT9+d/5GUCFk3AshDfTRyr+j2Fgo564UoM3QeR8iT9CQ9n/+EFMf/A4jsDK4
WQf04Ll8Dw1HKue3ZQFLkNuijOiZEBiojSxvbiIn1uynYanjwhaSA3vfsOh30YJl
DuxiqyYAmhJbdQeIkU/4z47SUeHVmtq66NbmpKl3yqV1kz1LLXxjM7XY9bTkxcHr
nD4K3sZiKx75uYziO+9ibzojKysBA6LS3P55hsh2V+3W0QGIiQrLqy3QhNakS+A4
BNYqcOmUBMpHauWm1R3PE867e3A4ENmkKU9dSzduczWxiMXFG2nhRPvaez6YV9yn
23w2lgIVuiUj4Pn0NVma1S28rwfwfic5mc2A7b4QrNGvDXfjpWdMecpOYWIag7mq
inMF49nvWW4tLgSIRwbJfqIHdSDj0Hx9T2HYHMzVWNDvJFk4eKrQO6/QjCQwJKX7
D/y6SVgXTUZ5P3XXgDWpOKny55WVm36b+C/nywEtfYjQS8khRcYdf3PdPoIv1fDI
2jTIoCGPxxLtlYeWwDldwfmSmgaXP/9yydAHdR6uCU9ltFNVtzYuMuFFPo/zdjwy
hPgqoDBVvVwJUVt3vRfphDgtXm+nBo9LKhHbAdrxkwltPe7HAeNnbj/bKPETY7Ve
+h+PauH2XhaydIzfz08HTtI6bKoIM7UAK1JL6ivZrkRUtikJzxr1lfyWlZ+7A5Mi
ndkDEXSsH5XFkJFXewIDj6Ojk53nrXfXxPdVWeaDA2u3rV2D1giG4eHCRqLeSk6w
uN9Vtsp4i78WS8wyEhk12MFrk9cTPUAAl9JqGPoiZIboYNOTLui6GdWoGcy+OznN
QJqon3hDkhRV0FCq5Pzd0l0E+ZyjofVX/IpFt2bVc1ViTZQ+M8ZfNl6f6RO6ZLTq
huQPYj1oo39+tHICp7FPKa82kZdQa+wtEDh4T8UKX1H8fAPz8bf7ouQpOYLFRkv+
gN1277ounNZwTcKm0gVMpTfEz4oEpzKWqdU8l9nGS0GFky9K+z8qwySrWKPCc4W2
cDVbhkd4toKTTEcL3hTeHD7RI7Qw/FOOn2ee0Vm7/E7JCSlfAcxtc/1U+4ib8qvC
c2noeTBK3B0yqP12t+oM3agkdpKxXmNGBZ3DTXiyR2cvB/fgDrFV+m/nfN3wT/qU
Kw/f8J01Q14e2YuR3oRU4C8F69S+kFXY1VxcoPzOSS/Rp5aj3yC/OV9HAHU5Q4T5
2CtRvxk+4qk2Fs4UleNwVJ4cU5XwFBTdkbD7hyX7In89u1w4wXn9vapOZiWOSYHd
m2La9QnpBNFnBsTN+gWEtHgNiuctKq/f/KdzLe4KJuILpfcsGMEsKiDsA+F34n17
2q0uY4X0474hWldDS/98Q7rfKThZED9F5b3tO0PgyvrvCQySHWZe7eaYaAGWAIBJ
xHkPE4unki15TBFwEXJz2B1qWapDW8cKq3czaNqOiibapTXFF0VYIhhwxSXHC8+2
mXa0h89MhX+wjoZdw4L9mCmk/lkk5iBOzw6DSDE9n3zw1Ll3pRZ2M4PPisykE8UU
NJXE4DqPWNOqb5XYEy17+V5mqTpcnUJD7d+Xyw/XN8K5gUilslxTf1C5sf7o9z1T
MdPbpwF5eormzUMDLMLEAEHQdjWQ7sUfv050DSxZnEuvbYfkXcI31jUKJ3fKwZRh
9opjUdZEWso4rsbo1WWsRlZYzQbzDUGfF1Vvvf/mijeDLjvxB2MzqsKqrgvIMPbt
Q694/d31aRlbAHkHvsnu8COODZwzen2Z5wAzxHlDsvg/cFRWG1oD6Ly9zu5v1Ans
hfFJecsUjrSb7uF+1BK0jMMxaNcYyyJUJk3u7u0C4Aondpe1ogaMS8m2YuWREuW+
yAKiOJarl2y3D7uIuJbkWkoe1L/YvIAPU2WVuRG/ArgdIMNEvc0j1Y+D8zl/iUK/
GWfGii209gEMrVYC8vSzdy9Gg2htCoLPdG19EZtlBdrY8B/btOV+s+0pfuRyyNRL
TUq2r6G6fiq/2g3jS5aakqQyD2eA1sLCgR0pJwOSAgVNfsHGxAB2WO4z5LtI7kf3
ruyoevr5EaTd2o8zFyrqd74TM1NoLBE64vmoVO1cWiQUcc0qC37/s6uozAk3ziUi
H639nGJ0bmVlL3zZA2tJhFXjeLCdIywk4Ng4lzGhunUn88mJdbKCV9Kg2E1nqaYN
Y61GG+EATBKc8jjId9geeWHDHV/e4g7kWevYC8MmU7n6Ul6S/xT06tSonA5Ih6cs
0JQwcCK11xK9kC/2TXl6WBD8TfNzDXnhCOQgV7bDU0vL6kh5AyaxucC3Db1cgc7n
NlFWqQ7gzYcHlB3h3WFDL52Xq8hgFfBcrhwuy8fR6KukdLI3SiTSd0vpmhf8xkYb
SEZO7A3scXdlF/1zyKdhMueVCjk7QQ7td1Py8JNO85noVc/la8UIKkeC8Ra4x0sh
hkpaQjhN1idctTkcV4iRieU1L253DCiwDsvhFxtVpbAqSKUlSVlKKN/kydOqi8uW
q5/DA8ynWbs1pIHMqC/K8G5LOy1y5ECwXoHC7hvp574R7ZYxyhux1HJUuNWvuP5V
UjvAEsT75nGDNKulq3y7Ldl1a6N7MdVqUvPyF2/RLBd14IC0OX5Zqw7MLwclLxbD
0J+nFnSJO34KiWD4+tspp1eckb9fLBDSLtmcZsIqBAZOzolU4CwtXbuOBGuHbkBW
tqPR9YkhTjA+K2bT9+nj7r9aM3RxmiEgqCjT/y2seTIQW+f7RmhqzTzO2aGqroy4
OPqHEL86pvieOcPfO6v2+TLY2xVjHr6T7IxbvHYTg+ruwOSlH2mpLKG9Wmg+jOb/
Yb8FVvY5pVI6WChEs1ja0Iv3d7DortASgaeQrAEBx6AR1Ywf64JjJoWByENaP4ye
Us6viuHxYWRKMgrz6Xd08gfIfSHUAjrf/jPQpgRFDPzJaVPkvftA16Jjc1WLayoj
bgVn3cI246p7ZvfRYKIDJ0gO5As7Y7aWeVMxUyhji8uRnOXEib0Hz0CElRFZKpR6
hCKdFUvYx2X39MzIbDEkt0ddKW245reI5NmTHJoPl69+wCl5NHzFPSItLUj7oJyr
8C6c7Zb+4E8TH68xVgW6WEXYFFhQocN9i+5feiUEtxlB0+Imow2/t8j4OYuWojCG
BpDdNJu1fxwkIzZw3UTBCDL6jgVnRDeKDDnzPBTvoOVmqwA/0bKsYsTTmo2idczU
mosZJDfl+GhLSRp6tjA/KQN07vMwiYr4eSjhhnJA9TDksxPigt7sAwE2BIX2g1tj
B+M5cwlHOVrZz1tcoAo6gYiLUUE2LGHwqSPDqZI/ZiwUV9P/n9kc83ZWo6AErBoR
Z0CXcGnHqvhFrfisNa3NQZteoiYEqj7aUt/dT/z0QX+yI0LgioLLbAlIXyzNW1Oc
gX/kMfW9kricc0mGJ2ri7edz5RhO1mdtfxLP76NrKEfLymqbeCyGqUzH3GbeB87x
iPOs2ovLo2WU9eVGttZKYCElYtvuTzGTkyZ8WwzkmOK4DtmbKJrm45rMysDuuLC2
Z6OKJD+egN02o4CvdeVH2gq0IO99E5Oh4md65G8P6V7xi38MBzUznS91BhLMi/wS
OE3EExpoy4yZnfMtyws5CIcu5wFo84xmTGIK/qTincVbVYKdGlIqT4u+k5r/eVS7
jaVLWrIW2Basj2KXw9aKsfMNckdHfpEbpn4XWday7OFnW5gSvK1oDjkahfeDbMqS
J4cS6SKBYvp+jWcjILr2n1yesN3DNf4sHQ/lzBE3yDw8NzH4JygbMnblUnm2bndd
XcWGEuvgxwZrz2UOECpftjRfJwOoOnukoTLquy0z2aScnPCkejZA8DXeZFx1pJR7
eASEB6Uko9tql5i9yYaVyCMjaLmpztMuMDXq5LIkPHReZyUP2l4MywG+fTT3pAVx
SR0LQyBdv0s15zHdgRafnjCx8C7+marWtgRy3VoDRSOGGM8/5yInyqMfoMJUBVmL
C1YK3fvGvxVCtAO6x46+9WR6PXp5ByOLZ3itDYEg1aMa/AwTu3o8IfG9NFAU1/kv
Fu3YCm/pcgBMv3Ja9W1hMMq/NfLRXbFLQZwZEzCx0O/oq2mHuqHRh+let8LVdp55
qu7PiKTDK86agukBhocjzbCTW9fWHeEl5fUjLH6QatOKw2okgcKm1jRSHpF9zrGc
grBav9Enx/v0UWPrG/Y0Mq5Fa08g+9eWYcwBLvi4BV4KVbvvLRgmy3QjzIsg5mur
xEk4OIPFnnRbhPJUX0WY1U4xDhOc0OkW2rho9WfHHex+x1s5DKIeb+AIBcCM5OPq
elupv6CGW6BSiWk06Sax39Y+ZfIObXgdvDL6pu2TrHFF/nWRcny9VTEJHOBjROge
xcUdaQhuhJePFEDu9uMoYTFl73Otqpcg9o/Esm6dm7fQcTfL0syXBeNNGr0tmohD
XT+HTvE+ygxJB8VTSgkbQfPNa5dIMpY8/qxYFUArKR/OphtXwnby6xLylmfodwQX
FYjCBtGHeKvlcAkunjYuZ8Ild/lAxXJPYQfTaIovUEpoIYvyRywJnCz8Lys96Orq
c+IIIp7PVMSIOlz4a4waPNZtOVs6DhH0InVlXrmHRuQIzBJM5UG8/c3ha6oyHwJx
6cX8qgvdIpU0Kf/C30PqaStAz09veFYqN1gcl92dLc5HX1oB6VlJHU4Z3IAeNHPk
xpc15RL4QI7FqDdKrNnDTXvC2wC7KY670OlA/EqTA5tXN1Nr+EZQNc092s4q+P8E
wPuz8T+/6nrNS6tUzHbGK9SrQ+bBgv92bCZ7obWMFYDg9RBdd13nD1XthrkepwHU
tqiVolx6R8hlrGw5lqOybaTPgjOVotE5dic6ZnfavAjIKbviXlFwDCl6GuCY/QOX
Edjfz+xQY4HrtODHnFm4eRUq/yq9DcspcV9WdCsn1vye8H4xlEJkWc84olCdC3+B
vTSD/a5SwYhHiUoMC1qiBkY4uxylcWec6R7OWqe73GgzLjZrRLZ/+joLlHWbC2cm
hk9lCKfSIlzw7HsmZZ43mByjJ4OVR8zbj00VeeqE1hdRWXK2oDxXezP5mtW0ovmI
rYYer6M/fyNfKeHHmmer2WPmvWGR37vHIIr7ehoP5BWCGYER2Wq3v9rKv5mT5Bg7
N3NxUMMFcX9l6EWOUeZMWLNgnED3+yUaJ4Q/MASraazUacIONOuejThh0b6rVmu/
oJlRucOi35Nvw6jJouUd2j6HRyqnDtmzcDUKWTUD3vccSVRmI/9AhLE/OGVBPu2Y
8I39xuVcC4m5skcdQaL/dBxgw2qaemQrNROTyOk7/jl6GUbmhGC35ZbHsrp54JkI
qYYcT2hFBI+Nc/C6JsvtJ9lPkYS0emY0QLIirC11+6Tni4jyF9lFJtcrjq9PXe9x
nwjFwW20BUZDF8FdZuI1rAJeHS4Ryee2nOHj8knRf+9hJIXSZrLGJSkb0C9lMaiu
uodbPMmVF+qksDzgK3nmaB3JoRyom5G9x9KNdqVXF5VNnStZtCL/uQHoBnuJqOf6
x276Hg8ak4JVe/z6oh28V/U9AO2vyJnFFrB5jWkHDjynm2aPyYWlGiZsFt5/iAUy
cACNlhw7ShoFS0vG2MSJvVMsLPc/8rG3Wf4hEEW2zXVDRwVQ5tqeV4LXXWLJNNoD
5Ct37OSAhUyTLVIxxqNNELM8GAJ4Aq1AsoKY/AAz9U/i0bzncenwjNfEn3jRE3+n
PS0DfO4aPL98ue8QvQdz0M1aXTgkCM8pG63gdv6ebDYK0Ii9LbIJH5AXCV2teW2E
ZjHTnjiEcNR6JMI28i8f1BJDDEH+dFy7NkLuAISpc9ogGtOixJmg2ZfD8oDML4R6
LmSJtUsqSmgGnUFDx3lnM6KzdLsohLFkCMT5VTrmBIexr+XPPrz7VU1WSg2ShtOY
NJO2jGG8SsvEMWG2H7pB/FzQsnrtW3/5fmsNx2RTAqwxuBUPkAeHXW1MIQVQZK2m
o8fk/3JLCXHfFYMevi2UuAiRkIkxD1W0tOZHV3rpQWremOJj6v3O+NC3VdcmRTpL
F6GhpUt1BXDpgka3UTqRF7/hgddars1URl3S4lI+aj+b1fL9gPJWoeWiPivjuE3z
V3Zcb6jrI/aTKDEGY+SfY8BA8fRdt86Z7OJXTzW0rQuOX3abFIKx8ecq0/c1KWO8
sBinO66fvcPQzBRvkFFBVELcmxcgu6vU4VTdhwqgKuh2u/EzqZrbEgyK/4SeQOZ7
beuWnZPmubYFtinJ3BxNNbauyza/oM84ASEHRpeCx4q5C9ybPqpzHVU+he/YVS3B
X+w6LI4lzt57HcifebVzfTwU5NK4yP9BgwTiGYAMdbkIH94KobQtN+FJ4JrpjsOw
/8wKw8MMLsO5k52JYyr/MGtehoSsJ0BTrLIAkU3kizJfB0uhJhKYcc8/MP5UV94I
ThilCUNjVEoE1XKjYa5WmubUeY2BGINML0zURENNsPueXXFf+ZSMrpGfiKfA2VUA
sIzUBaHpeYNhGJhN8r40tQhi6PdQNOrZ8SaBr4Z+3zX2n39uDHXwY1wvbpuI8D7Y
/ShYMwWnWLp0WRCzTYiVxrQFwcUsnmvebVKLFeTIMr35PPWROuZ6pXMHs9Dk9zGL
58pKE4FYZe1KHrVFINfI+lD2Nk/W0+qAWbTchaJsViNbE6rsp/Dc0lcNCjYZqR2z
fu15Z3J3k8pZ/YHiby4ei3ivkuQOGlHzX33WhwXhY8q5nDkjdBxvsNzZVEoRwPOf
Zx2ss5WC3mdp0WxBj0YbG1q1mEi9g4g7U8WcaTcZSK1RWrds6ek7QH6vx4anAHkS
vXCyvezjCCFCV3sIsTq9IgJy52fw65Kok9rr9VJ9zCelcNmT6hHF2290mlIt6A7I
OvsK8cYm/EjSwlC2qs4LzrpGCd8qlmqqrw+YLi+m0INmeWFap+il+5ya7LDLoXPK
+dZjBz1StGn3ODcFFHvvNXjk9JObA5yfVbtqWKa49YmTLHrkOBj7kWuC4ZpPMq4x
lE08ZyT8EiW7C/qbrhGnMTZGzSkU9dLGrbB5cJQWXW6948eZI3Ll6AFzOMlJA4Xv
svlSdYz30CIHcnVqR4rVO895q+CeTQPf7ZtzxkpJta32n94QXae68U4hzdhnCmzF
/3UAicP6XiHVHNRQtZNOsrkSMA/j+sSP9DY0+rwxHK//xsncC4uGDSKcJxJpHmx7
70Z2riMjNzLspd5ZUQ8pzf2PH07K4NMWJ9slPkdSSHl/vzBV1mPcHXTDvGTS/Cs8
E/Doyd/6KqC+RvlgsQH02U8uMVZKRudAinFyN01FRilI6DwnOiOfxbwAb9QFJ7Pg
04vjoFcMxAhtfpum7C0oMjadydHaQdRhsrDJJj7yP6cMTM+9R1sC+1V6xpaheJQy
0vYJG57uDwFibV9tzh05M+3FPeTaoNe9fBDzPIhZW85Q54/raiddIlmgrvWu35Qv
HXJECLCn831J3OPUiq1nzcszRFGRmm90UT37vzHN4UcgZ6VDhHC7EKf/uSGt1mOQ
YJqC4VjyefiKq+n51FKZelecvbI3/jhIp9ySwOejGXYiYEYsTxNL1hHstnsr6Fw5
aIyv6fjN6rzGeyS1kwEibeOBsLpLcVEF5YwI0naQKQeyuc+pvtsSl1Gqx+1TyFJP
jwHUag8h0Oeb+xun5gk49dNrg9rotkG+/D9Pyw+mzWlnvgp+aj+llNJa8gFIUPbf
EUfb5a7cwnqwVkxiaHevNiXKyP1ynYRX5lBaa0rLSYIIaYsEVNRd7LzmEjt/IY1b
6vpwrFRFlMQ5FYvoGvzS8kHMPgHFpV2tuKiI9/PmIja3cKy0pImrXvPoXzzrywH2
vMg775PBzsYk/Xh30iJ9B0y7evTqkz6j+V5wwmhmHrVpsTsuusSSBG+dErgePIGC
6sWGKQ413X/sLKZkzmUggLPGpGUAgeSzyYFbxv2zDDEpXTLF6WNp9CTIYVWhVTXV
7NUccp1Ig1HkCi314LiyW47xVAEn7WdX+kM9GojPYOJZkFfS3jiS7etRPyOCgiYm
MH3VkfmH77NOJEFhGemi2ztU9WxUYlkDJr3T5aQd8rw9xCQnK2Dmj9qz3ZGL0inC
If6eQTO6jgpXAXjH4a23HiK8lekYx59KPy9hJWfFf+Z6Ark3e2t6sXnF7BjEyCv7
oMac1ubxEyXhaky0zmZXtYM36UuxkWUT44FINGDV/sI39dI2w3mFu2ujteZFLzjF
aHdKrw4C0oB65hjy0OP4Ht9BrPv6UB4CI97nGKbTyTMly+FJaoUqTS5T728MftTW
wTzNlFsyv/t/erpvc9c42jx0eL0hUZNvNEYWBBcxXnahpbGL/BrIUXUulcTRWYf+
R0MOc/TDcV+i222by5sxf+ACPuhlq7UwlSG/TK/mkHXeuniGdj9SZvy04l+u7O6K
315Y3FRTDTKNSm2B9WVNrYgDFjyB3N5eF12tg3gE0POATWSvQL/vsJMTkIi6NJzt
3w3aXdWe2jmwgTGDbdJCglla705p0uv1X5R74DqX7z8/KcyfuOqQ1RRAjcm1NbPQ
kBSZSjL11uajaW5sexkxEEmDsuhtWi0yxEZbB43x9LKFAohB3BSwdzEuM0niISJ/
1ftHawvYS2EtNRQIcu1GoGPU1jt+vvly/Wi8n2+Ig6d4+0qaQJHSWK1QPadMbYI8
e6dln5PazB+ZN3LcBHdwau/FCXEmvicioOPHazndDD6Xy1rW5I81FeXy0WX5RuOZ
ycqEuDhpci5G4r09NIGUlLztehYaEJhUD3yF7e3MeBqmUtz7xVOXBI2pdzlbOfR7
h/GXd/v8ETC4YmD99ioCB3eDvKYMtPS0uP8sLX7RxWt3plaulYJfOASlOtNsubJh
3auxSbMlT2u36Xpe+W0bzp4p6ffJyYbXJ9xwqLoJFPQUthyaKK52LbFJq+4XozwA
OYh0hEWerJmk3cka4mwYVDVVEEVFqL57g3KJjA4iSkHWiIEBGpqMz7zS8xdem08L
GxNq0ybzZDMvi87JTeoNVCn9Un1x59iucSWRm1152/duY1KXl7ElkV7ww6JZw1vT
VKwSDncngSV02nsdsmmagt1OmlpLJbAEKRpoCmbs5hV7pS4+G3g4/shu13JERl/M
Zzxb8x4RmTQVP+L0kTikKMU8YyDGn8T9nJm3hi+UmNt7LYclqkATIYFkWZavaYKu
KQyJIF5aBkQ4kfc0IWpqdQbeClGuRgUQhT0tMspBHRuCRwsKfr7PuL0XiCAhMPGU
qh7VXH9k1Hczje1ah1ds081Qj0FPgz7PpH71dAELhjRDVXxyS/catX7VqgwCk88P
k4vPfbk4cChcz+YmaLdfyQuzZUoTA4Ny2/SLcFoo95e6pOLJKsvF/5zx6icm01ON
9IQ95mV6g2bVKeA7dGmCxne3oytxzR3YdJc46/asNujQTFD97ktDtKUU1LYPFAME
7XkirPd+fYQ4mmqWQhMApNgXDOnSVQVnwiQrrKypMvE=
`pragma protect end_protected

// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
hVNItvBct+ztViN5lARjXSDlXmtP5lYhPTRd+FlPxQrHMBLnQI5MpN9eo51gwZ76NQFj7tF7lzBd
T1ccurz3+9ohwvW+v3aiIU7vQulmCNXEMdJxQpDKQ/snvM+G/ujbsFHXLqmZIs8c7xIwvOptPOtB
lWfIRN3GR8pkrDw3TSv9Xrr/Z3vPkNV+joLj3uIZTvgorsmdvBm0aOFc7hp22HPIxVHo5ZP9bduB
/Xk5usuF2qN/i9P5epaqJoDorEjuTCortS16/tXotQ8SW4TEzKqHUhsUYQpMCVzzZ6oe/AyBVQKx
24YIo0haHtycFiQjR91HHnfB9vHHrrxGihJ43A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
AnxE1wwaAwmx79ifmsc0Rg0Ab2wLQ5oQmbLOWdspheWBq/q3xvbfJmrCXMKn+W1D2hmoDYSEOxv2
XudWqWYErRIx27RScIiUNRZ6dR9U33dzfBLCiITG9NFp/YMc/zaIshvpFgojpSqlAZ0I/JPJ+Fti
wvtRsGy/YFYFaxAR7wuc1s0EbSH49s5rEeVsoid81j61zYCS9K9gwzMxk26mSNSwsJbrcS2w5M/t
gSXeq/9wdEdWNOsgsIGdncIjSmH7f4Khh61J/St+KFtUQMDpep5GEWPn2/nzpQuamoYivkQYGPdB
sSc+FhD3ZrKlumvuc3cWPDuANWmYso1O4QbYoygdfLiwdWvquHAukpulfgPj2MMKiOEg3Ko3CIKb
Wki4DwlFTW/9PCHubp34qjYEYmrXJoR8pGOHLVu5f61XrIqk6YEllMlzSpEplIt5j9cGVcpLtgxc
dSebfrJXy/0a7ptNj1NFI5Q9FeVzxVjM+f0kjzhXWujv76pUyARI9L5/jGhU+Iybre9iPAh21eMf
10gyEJfC9wdc0z5op7a4AFoZ72atG96b+AlLV+pV/K2+8Zd87yXkOjdrIuKWOhORXDDcmdoKVpno
FO1N6tErGwf8jw4bvldW5Cx52Znz6LJ2u9hGRdcwLr60MNih5fYFa+7IGR8amVw24P+9bMHoSkhh
PxMi4yzSDJMHGeR/9shvbhAf8wwNycS7QKlYFFXcpGvD3k9VXrx+JnhjA0Gdk+00GPk2dTQJ7krW
OWIndJmFOz2VczrKl9vpnM2rbTFYl3f4YzpM/0KPGRb0Vo2Uv4WmONVw2iaidVh8IYsrLaXb4H4f
pGhY+2BLTTa5sIfj3MY82id5DO3VageIFoZ9sZHVNJGRQtRiIl0hXuQap0aPqYdJ14sz9StEBkZf
DnwW4wgCygEmF/odnGOGNokRvS8DHYdRVSFcEx1FZ5ij2rVZylQ4VtjTxfbpkcltlXHc5cuqK5X0
/3XbsrloTRRSpIMWstM+90+biSZF4NK7pR/zqQiKEAOla4Bz97zofR3JcrciZO8dyWCdkGs155MQ
v7t7GYUjDAOyu/b5caccCBk2Py6n27ySpTrlKK3fvMFqvRa5M8rBfJc2MGebqK6BGuY+R7xOMIUT
JjjdWgDfpkNN04XxtOuwW+C0hOAKTbNm9xz/7vmwjS1spF4/G/zRRX8t8Z9jNhCSNdyh4jdeTzJC
JeyeOnSLdgWz4/VNE7EkhjRGSS2vITebWDN7kcBJ0TjcPq7r0/sgJVYqsxHN9NPZtVM1/FCRFGfY
XIGZ7vfKStmEMXumxUAX29DMY+4I31V63vtOFo8Fbc9omXbljXQr/Vk6G/1yG7oclAkFhU/hlcpe
6mYuyr4iKnsr/OHMdCp7JJNPUW0syq0BqoY/fTfq541T3mZOVZt3/tZUGulxzAXns56LHjr7qJPg
ETKlAGMSs8QqfNu+d86AYwd77Qt3yZtugUNfL1UTpGzBPbED6Cwd41kJ60xXvQCJkTAJtdRk9MK1
Mes/VyATuTUy53P1lwdS3Q+2mV1L3Cu5BRC9ZasSYGeXcDUokdvBcd+l+mY+nFptLd0Mn3Vm1/rk
uSYlVH349DlloBL0dzhQgsqD3LC6EWVFI/s4476Nl7cTDJjhrSolOmkEHE2luDft1b2Zy1IfUoE8
GpCMnsJFmxJ8k+5L/KIcdaEDYJwqcSjG1tCXr3emiCJ6tkpsEgX3M5g9SZwDOFRes3DGTIAGhOdK
tSZOKdNhTC/7CePlf33ESuyNjR4OYH+kxaIyHzjGdqBXDMi+cmOxLWO0LVJo3bwuzv9x290ZlzWD
fYSsYcq/N4UsLvHz9ppyFSpfePbg6BQMV3ODsJBi+EHG2psgTlnArpo5kB9iQdpKu4hP4i6YUEjJ
TGJPBbT5hQ87V5o9H1D/N/HUE4eETnuYGMnwMUTsyboZdkTgbchvEw7pGf6YkB4vI2Bw29++BtHl
o83Dj21zWEHSMW6mctM10M9yCodCQxyT8VJgFTnfwltdh53wbupH6oTnK9lgfffyPsvyJKvHZmAT
HrxHqbOX9dXNXhW1r3hy+lqSwTjy4Xw04GHVEqGzX3j7Pbv1dxnJWuFV/UV7PIUVmPhqvvJ99Igb
aSVk/jE6xFmso5gCfk1StM3yHWTp3s4O2r1Y+eQ41k7V3XXzrCN6jchYf07UYOm2CshMu8VcgjR+
VP8DTvzE/p7UeI+403Wld7vXpSrNpJbZehRekNjG1h8IO3iyzdn+EcSXelebe/Fl2neejl8VrDXG
nWfiIeljIoLY2KMu87Dkiv5KxpJ6F8xaCbiaNfGX1AQvB0a0b+1lMApKyj7+SPL1udo7+MPHj/1E
6s3yUWc3tltRRSp2M1INSwuZHxOCTdSMqD7oI6jmREAYTS4x/hHe0zNndon6dZaMi7+1HUf4cXbD
OwODtP7W0AzrBqEyoySt33c9L/mWRNyzWPL5IoGdhwLpeFm4INB+opArfFr/UkMDGfgJvgoRJssJ
UUzZnMjUoYY44IFCo2xBHSsteslk3yH8GIcmrtc7kF8Le+Q9HOqnAequDFhqhKyl566ksPWEHn43
JKQZ1rxpTjw8G1fIy++yYaQqyFmFoRg1I6kf6+0QW9k0pviAbabH7BTr15663isScatd/9Vtdu7W
ae3LLFrQ2iUjEE837YjK6FvWm99+jXSJhqhQx6MVynrf0MnFkbRXh0lrM/U0+RU6hRbvN80fcH/s
lDZSBVqWp1ygv/xhdng14CKc7+ZTFPhGJ5zwWEGlyqzz43KYJoZ+ddh+2xq/qz4ZP7d+tiPNEZSM
shmtufQVF+NzVkewzTlBYeIxjRNMpZxr6hliPJQwI57oL8/R7wUHKb623umJatAYdoPU/mhbOEom
WPMuQx0diSvVh+L0JMOILXcfAdEYgEuJq7iJql0Usgqu01NDp5dcM6IbPzKa7lHDd6SBxCm274YF
Ox2sQDyiZ4aJjsNo2tauD7S3ESRyBK/Fh3Q1U/pIPJzYm6Wb3BNp7Y+r4Sk7tgGkcWqO5NJj2fqQ
cRLMRlR6fRjeRqLzuvgj3FqDn/mxo6xTLWBVS/JtCBrgUtKEUv2N/kS4o0LU3xkeWfIUvIuN9Zck
znGA+mWGaeePeWgxQ9Y90DsLBcPVzcmbJRoZGgTVtmO2CQiKks2nfj6805qRvMlw8gwodrwdNqbc
uoEJls8RFlmz1d4TWHVfOM9f7yfa4j5+IsAZn6k6B0MCvoMPkVn2uuCXakwsHjkIyB3JN9jJCsGo
8LgzMygitVFgMT+/6LXuOrEYs0vYkKn6pO29nvuPVkR2UwbEtC4Q4QCtF0if57UmTyAbNapcdcA/
NDhDD0RFzNEdifDJoNOT73srYiXmr7o8QybfWM40tnKVO4q+32gx3YcI0qD1riUkzXAudTdIKPxX
7QQ5SpMSnm8q3V0tAfNR0TyYzy29Kv2BuJ37EDXU42wkOdIU6CLmHemWuweneAuTQEDqGjUGlEeP
SDJCvTYoklhN5VvShpoQTW3K1a4tVHR90Sr0fHabkR3c97Hzqhc6McGmcg49xcMhPur8qU115Map
+SQk3pGF4c2lpy/15Yry5a2+mx1F7egdsgz2EnkUpCyFogtXowvx/XRS51uBLlx5tdCE68MySA+s
K6AtzuuiCsHAvSRwGCa93Fe+9+Mnonb17HDSPcbJS7xzF/t/FAqI/cS+s55SDm0Jtq5+TpbDv+Tn
YN4tY97B/NwdcXxFU71ftCzaPOLl6kkALGA9sNAf0Ucy4x/trK3YO7yN1IABAP0zgzNI8rDIQtIR
1DnGlIgJ+HUbXIYqey7SQ2N8iRvabTwEoHEgVj7mOTIncgKN1Nd4Hmi6z0bfrw8bMoKQjf3M9HMK
056BxHobfSXkNoAK9b9sF/kyke9y2kiOdz5/jj6RskGctP4AXnd/ARA5q2ajSefCRd8KgN3pEECn
t/1UF0Oh5O5+asWF0g6BqbNIINi+AKKIQf2tOQRaDwxID9Oget8WvP50hMdU4NLZCUaM0L3Xfo9C
qHFVwJMQtSm49UQ+oa7HG8E5bNkLR+Ng0ClfK0xECwC+02wYSTlYFRdpD/u36pwUQFl/hBS3qdgL
XDJ492qKsgCk6GXwxjqH7ZgauPQsmr4wqwLe2+df0lKHvuSGdYoW/Y5cj7yEKARCsO2sGV0OLpEX
ZJUCQjoWSdSLcRUFTJcALYiHq/fldsmgRNny5VZzPLQ+0u2NqIlJHntiM6GP6HNc1jCB5GK6QP85
de3VhK/SDRA6xOhRuw6okTRV9+ZkLkX0BCvJeSF4MHNdDanT08hit4cVl2egEC0RSSKoCykZKjit
4yQrFQHVmeSGOYc6ImAA0SIrm9b4adNIm/8SQM3zN1eLLnewcaUcC4FUV+QVXQ+Khkxf83h4LBUj
Z97LJsoKyOBIWVkCE7EvuFeaFeVS5NfCA7Wl2d8JuIAygZUhaeaR1/BQ+wDxDp8apaPYXvARR9s7
ZTeoRuP0qlTC8IsP58dHlkBXcqEklMwYCtGiH7c59D7RGsNXf4m6AL1mqebR1nLL5jQBZMt5inzc
rToWJfvqslRAqR3J3pazelXWHnkQ5/UQMMdqITCdMBFr0lxcdpSwEMLZsz3dAjDojoUjEaovUS/K
hg9RsUQMdg45Cjb5JKNFk380IV7lfriRhl4sTv/WzEJdhOophG4XCJrMp0MLr34iOM0oM7cOAlrB
nAd3dcY4HOi7Y42tafrSeRxALqEAXz7X7Ef6a4cTJGHiSmIEW6GFXh9JPFV5NyqKsVsdQ5sWoyAi
jZdNO8uWnzeQFU1haM14IQO5nS4HcUZ6rZyAZemMOnswsZc57g3OfA+ri9/Vl3hgrkANNskVvChC
IpGFunVAOfqdyFt5eAmmu5oz26gRWitON8TjDC4QoZktBI0nD5RpGE8SCK0NRpRwN1ITasTqssQM
yg2f0ojWwdWeDrNKuxd+rYVZW1YJlPCULlmawI8EDq6w0OvUmNI/w0XoZ1OTHDGWqmy7mdzkMLj5
1D71VEw50z1qEB3KWoTv0k0MdKXDrDq2Mo8OxzhLRk+ULE26MhjVlbezLE4u3DAyaT84xWLKHUqz
YN7fNXTGTjLywjRYyVJ+PW313Czxba7NtzjpscKQBvvIUFO0Z5ngZS40b3ZfO20bmrW9+NTOkZ5j
0hPF5b8scV+K1OiJ02f5OQNsVtFDChBUa1cJQst+E6wFJnvVQWmOr/hl1rKNh3Zr4hqmaqORIv31
MfAyUzT6+67HoC93jqQjcLhRkgYHa58087qInxgtJDTuEYxegmu8FaOrSZ+vKT/FRGDAY4sflNA6
r0IIwdlpSB7JYmnzuPcNgTiLHvYi8Ay8DDSzYmI9gLx3V5MUxtUc205jSoOUYnmaAkxxILM1xT8j
AKTRoGLbteQdSTYh8+qenpac+T0mNE9r+peJFKYHcJ8o6e5SebGNca6ff3HVG3ovPscFgDUJvsjD
XEGaUJ5qDR+26RzteZ5cKqDg9evLJunqSQ/PzcrIvrm5u0LooXe6fDe6KxB+DUMJEI5p6XE5au9+
pqr3FLbNuH09pIjbiWXphH6Zp4fwAQOHRDHgdEsyJVOjR0+MdW0Oirl58po/idl3wRER3cdiRU5Y
W2SFVetjyrpHLl6+Q30Ouugmi2TO7z9wt4qt/qksUu2ke8l2GGBCJQ6YJ14+bCG8kq5U6F6P0XaM
0evRY+cJfs3oekiG6RA/AX0qpWUpDqxeZfuadEzIX6re0cBmqwJa9Qd8J4XMQ6F1EUHJDpmbrpka
6U19l/rGNkdMNNtZxd1tG/eMNs1uI8qEjWHEnpGX9wqcD00VC1Rk6vyh6ezfIIwc2whClcqpjM2L
NmwB5P2iX0GfDClH50GJThvYzdeDVgdTWNWrdPHUOq07nGqegtrSyQOu1t4jYn4Z3bLM13zILpwV
uhAmQDAL6AIeumZZHpxqEXDQGjkhaNj6D/LMxS0aK9CmBSW7JY44H+/KQ5ElgzJw/E5pbxNt2NAm
2D8ijlIhCEcyuKJrnIY/VvIkDNqt1/XRjbD9dQCtrjeAZNtlb0VQ97vlPN4KlKt0ac+AVHglCni9
JWtcltiOzYy1h/ts7X6J4ReqxCrZE4NdLc8n2p54gL2BaUKET4YQfhNiTQysKsdsDvTz1Wrb2wLz
DCQkDB5T2itWnJrfYSQNfXecAr/bmBw2Iue2NnoMQ4608yLPuYqFxbJ/oAKmNlFW2kQANzQsbyXC
gz8Yyo6MAQJqWuRaDNRknc+yT98z1XVTEUwRb+YLqYrCKKLHwIYb+AOn6iSeBs7NrTBW1lDdyyQC
HtUuV86d/qT+eOMHiHGSYdDMxcE9q7AmEptLLYRfvuEvsSN8AkH3bcRFjOVM4GB2S0kXJOtyPCId
3C+PWZcEzd97Z3N8ucNXMswIp7smFkekfscll2wV8KiQEsDpz/Fzk0IFq8s0Ng3t1zQ0c7NRvfw0
4Iy6QG4x6MTArffKsDPh60axrrRThR0vOw7BPN8y7qYOwbk4zbNi7nwBOCLQD6+SAxwbUryUIFkd
RbkZoD4kIrYTrYtVVvD9mC37HBfVsQ2pWNGinBiaJMpdqIOEQpbYB2FmsCTahOC7cnPuLkM/x+R8
rilnqJWoSv68U9g8YSZxFFt2fhHW9C6/fKHbpViaPeV7/Eo75uuxv/nf9bb1IKoqseyj07qDxSFb
bWkC1yKYRIuVwZYUsz5iw6Ms87NFOkEsIr7h+S/ZN5utRedzKfyqHpZqeDFjDZGp8grz5yR+3nqq
u32GW08Se9aHea2ZYoX4quFNEytfcWvVDM2pvN+4wsYyXJG0qhTTnUPKj+YidB7tgRXo0d9Hr0LP
3nUmzhUtALgLA5mrodHMjHnjwJpcuvBTr7aCyQSF2VuloVioGaU/dvJCNu1PMIYIWdDGSdegT9Eg
LebGSX5+6n/3gvj501x5NtH0DHP2cPiy3TqFfEWVDb91i9CA180z1EbEs1M5u72un8l2k/lEQg05
n7IS/6erTHQsPs7kYlUZGqunnNs/Zb/HfqMS+1eM2vWZLlHgPQSFX/syGaJdnHWGgUDNMlxcgufD
rXxuM6Wn3g/BTPV7VvPbone7w++fEI9KUbSKfbOHHtzw9RBTStc3w+/8pozBBLOhO1rp6suB6grD
cr1CQSf7ECN8cMH8H3VekaKvS7pBWWar8x3iAIaTrlmVcNhjcaPrI6QKKE+namAPLjbvFvHMuaBK
x8MCkzBLR7GM0aoCAJjcOUMtCYxMjVYfI3vNsPKRrnfxmHVGkPjhz34nh4RGazxIkMvITM5zM/TZ
53ZO6qfw/fXEaYvCY+aHq0hYahMzybXP2WP6jbZxQBZdIKy7sYfENLgCMPcEAJF+8HxkH7tHKYqv
zfBH2mqOUmvNj3nxbv2KzskrKntY6PCb0RXAO1KYnC+Fxu5DRkHaPqmDRkGXe6G1BY9YXHSrOVIN
Xngf13u7GxKqFQM5DS53rkBMMWl9DCAJl9ecGJ9k5wE2KjDtNtCzfYMh4JCAZ1piTgPmE9P04AvX
gCxB9j4wTdIos0OQTLdQGEI3qCPsRDnUo9uLOVGz5I3ZM+hy0z/is/bEIgcPitozscjXD0RlOtbo
Lt3iM7LSE4mPUzwEb/1V0NJRp4yooAZOjiHSLSIEnU+sWD9SIT3ox6zNoaMsAZ4ph9mXRCEOPbSn
B3sl7XhUBgy+QCNpp1ag9Wz5Zglz91zSx5JHreEB+1MNWimvnB9yXLTvOMWFoueu5aWPwHVuELpr
dW2SmT8R34BY+rROjgpmuHNmNpG5TNiyf7YGrjSzzz4rtW6ly39nXwhvVgMjgUSsx5q1OYdh3hSu
MJ0ZoUdfrPpEZwsyiMAd7tBpeIotsO/T1OMJhx05kPzLeZ6iZK3j5Ggs0qD65hIMQTxHVSioFTkA
/sn1LwgKyjqP6cx1SxIXq/x3YF1NDwFJr4DESV2uOX1lIFKDeafjlJPSm2GOvREcXyVowcoGjlQc
cAxuKKuF9CcuKPEwfwaXUDCSUaE7sGYrOPaOWUw5ez8dXtGKHvuKIysfJEHK+Intvvh+DyxewHK1
EVKAmRLzJn2yXNAP4Qe7GSV6EMLpJMWp4yQpOAleTpob4bM+95SgJU5Zs1VLHlhyROdoKgwNFZoR
r5/GlK0bfv24lSyniKLuFaLUL7i3hhpplywUKeap8GIqnqh8wpa/2CCaX8opVZOJH03IUAiGJR90
nOBhCHjX/pX0aFgc4zDABbZTd/Qg0gG9fTyjtFghK4HITDdXZ5yt6vYhRBdzSNWXF636t+dbzor3
RDBMOvsns3NGQxNaBPLVZ6RUT50aEoQmB3b+ZMTlKFPTB6xZE+ybgiapfi64we+0oSI6l8CstPcu
lH0095JDNjCycYxVzsCp6KEfWgmyPRmg93Vpv7U2A6ra57iJDB2pdmMlnW7kHhFkl+Mu22Etuqn+
XXC7OEHdZH6VJvfE6UUH76+zGOZYc3iekhc/SjV4q+ORE4SvXPXTZ3eSAcvVXa7lvyckc6s5UFpl
raJ+3oQD8/v6Gf+Ua1bkyS3wvA127HknTRTnd4hH8GumI+rd0BCv3xkKy+TMKNPfyHzKQZLc0y4A
C5dN/whJVeNdMMAtSCMfFuxIZZZNzdQ9Gdm5WCesowJ9eSZ02JQau3GdxscQd6Z2u8fxJtDDRcQw
OKhRC+BVmRivUgjoS6KNGcmvvrz3C4z6xleMI8nj0OekeMfm2zD2J6/KUqfdBzBpZbaLaKil1pvw
+u9PAGlp+tnntucKk3Z65U4ybYkMizbj9hDLtLTQ2RjKFPQMbbBYV/Zcv0ZYOhn2eIWS53yaYXOv
HZpgrE2/4vhQscUZd+agZbY57h6/CBaTNktqdT116HMPz5cjJPLces/Vf2o3/fLy24DngL8rwtvi
OcK/mpkb6XDJtjzZ3qu1BF2P/P7vU18AA/t034Sya1gFOPCoUmxXUrWFtfen/d7O9MIKfn6vtCrM
cIpeSMbUz8qYqpB4hC8/zwZdQ8VCgdl5E34soXAGSoxpgULHB5H4tAhsbJM6PWu2Hl6kLGT6BDCN
qWUueQA4Zpk/R1e/pf0TRLJmHuOOeZXdk44+PP0HJTjBZNC/YDZCQGCCEdAMGM9c1mi8M5yiqsHV
5sZroe1ef9O5uPQ76hHJkFlcBfLrZL0qzvmbtsXgW3sQn7rPiMIZ20x90SXzjJ0FV4usu5hGRhfC
/9nDZywfbE9pOXpV82mWgnl0nYAoLDv79za8tcFEK23uH5hsdnd0qzgZcZf2YQJ7YAy7ex0Np+Ld
eEyR3yk6xfFVkqeWw3Db9ap6Qp0rHXhbeOEeTx689zNn0hmCuaaOAr2n5/LVUqiL2QIk5GBNwfN5
vaLStFhLUU8Wod8z+rRpHlMXxGoit9wsOxgGVe0m3JLKSxwmjAimZLeq3KRBJHeEJRUKf9QIUMVp
qBSa8TKsHC1AYpN1SQ2oLxi6XyPnDcIotPK6GvwHdqBHJUpDJmm6JZ80BE5Vdil7vyG9sd15ewA0
IrUmZl+7JJ6QgNOUchlru2mi/vDrOLLHqKja0bSeGRD3VMbdF5Vb1n5fzfxTOOqpu78ocM9JuPzc
I8dZAIA25ni7/SYDD4dq44ZQVgJoCkypK5ycyEQznxok3KqZvzSnI5bMaFV7ZtOEl1nTzRWaFCyo
6Lu+0LPHrDf6l119bqYJ1LdiHPDXFPr/Ai5oeZkHsnQ/ed+0YvYMBJ7Wet19tp427iHcGFVUY130
cyF1uuC5O2I0UE92bNpT7hYLtdfoVJw+nUqy+uC75l3x2itZV5el3KA86pCHaiFrItXn3NAJPThh
Qv1T0iXwy157LfaFMPDaSuAEc5O6a+xYY6FYGkzuDiTdDZt4jOQwBMkMA0Y/ie9Jwhk4zzR91kS2
ZVF3ZHYExQimi6FrbcdJwTqC2J1DhibnEZqOm7AtuO7y0FilInk+P14MSVCEkZ+bxyu1TNlV4cTh
nL81Tlvcf1zRmzmLGoPeu9Lbx73KaT3ghqZOOQsc5pc/u1nwIwEouTGIMxpxKRNoOuiAqSiinm9Y
UVdlvl18hEajDf0FIAtMWuDDOGjTudsIoi3zc5YLPWXF36at4JZoiTBHbxX+a7yyNQ0FcI/ua4wa
6p0D1cftuMTrEKX8fi79UkQncEBO8vZzXjqVLWnpOwE77Ki54YRoqN9jCXbaZ4xD8jQcKDz27HzP
e0v5CXjxG3GqDpobM7rpUk2VyMN73s7GhR4=
`pragma protect end_protected

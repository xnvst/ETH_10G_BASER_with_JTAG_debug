// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:20 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mlKIeiXqYYK1Gf9Qy5WGyLRIh3Gx5Qf1yqWRQYg2E0PeWTaAu5SVH9xM1qQNz+SJ
lY2gCg1o3VavXzHBYk4ewBB0ZWIaW4yLPKxZ9A4Y3s4Yhfc9kWtzIIb7oMX0OQao
uxUFo5Rfx51fVGHetBUMiiUbWKkYUAHqCaCvf00wl/E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9552)
YetrXWAqnsJDT0cIYLVOYnMd8Kgg44k9vrj6zbZPGj7V/4i47V6WexPEnz8aox8L
i1JKxe6kZ1MhEQwAbgR9hW0TuwUyfROqj4vFKYIM4PLcTgjYKfuuYE0L2Yf3G9SG
GsP+QgiJeUoTBvTr4UQwrgM5Krgxzax/4sbXhGyZY3FKdJ7NIiSYdh8oDH4ruv3T
4l6+jHF7QmdIujIJCRRa6StSaS4elsqTZF7ZvBSFTkVFo/uNLh7G3gLz6AiGNsiK
iTc7pX8FnC3FsDAY2fCx7htROcG0FTl96XOVlUEulv6h76rvV+xLA5zWFrZASRFV
q1W+JWiGhxMaOVtSxhZoxGt+xP6FHJXWiKDQJ78/dZnn+yRT9FXowJ9z6hsZ9cy9
5bw06LikAET+3GcbWFqkcJv9P/zwtlCTiujxhse8RId/8rxOf8opkZiIWqh17AGY
ohUVBjdvI8zgD4bSI8cAk/Ot1PgCepvu+3YhU0goo+UjaTxRDDocJ6C1QtH3VHOa
YQrAZiDV6bmY2tF1euZU9yZ3JHm5j8szjyE57PbISeAsjfG6nWb4/xVJ4u36hKl9
38HkT4wRxlW7TlFjadUu3iZ80A91BFkXB9Hy/fGVY9b2JpQpee9H0qHh2vw7eOsd
k98rdSRfE1EsFriPcU6dLcSYXHiBJ7sZ3x35UrJx1pEEksg2ANbN2LVi1G1zNeJ9
bjiHWZ3joNFNEppL908ACeZtRWiKKNtQgqc7lswwC7QQK1O8fCHNQ2T1WNgggAn/
j5+vjQtcJBQIkOOtjKhUj96db19Y4nCJyG7M5Oaoc4oMKH3KoxYXpOuCWXFw1kJo
Vs/af/5HG0NfrkDzEhzyXCrNJzn4ypqcyNXrquIX0dL513JOVzZrPR2OAo4UfQNQ
/6DLNZg8rl8drAVQg3DdZBQOAjYweVyLmUm9r047z1ycnJTJiBtjIzbi2ngmzNsK
Iul2kw1QfOFRk4B3j0PiJQD6qOSRdnegeZvyUt7vYoi7g2Hqj30OW8z44VqG+8ko
CQAdNDMZHnueX/deKi3dBcUe4A6MeQDPxMU1BHdB4nLZc6z7NAh41LDRXHzQM9EI
9CIhGDWbtzquq6N9TLvI3l8PvUKTFAq42HrAG2ucwtlaEfYDsYGsdvYHK6xT2ro2
xKkc8F+T8dE524wHAtASzHf4dyTRO/JEMijhKuprxCDelWWgQAFvbInP1hYTw/PG
b2mEz9Mjj3faf+zGgHsQg7DFJZi7xIhTh71akp4m+x9cHM+GvH8ytyQhDojrHrtM
TvGh5EsT2F1CWQNaAE0MxTMKaDtbCAemRHH+VkHjgaWreRRmiacULqDOKtZlDmqj
SYypbBJmzC401EttuNl7j16KLjiOQ7IOmLZy1dqgigQbOisiUeX82A7Ig0QWDckV
Vn/BVwuyxuT5gKi+zFlVTKS+NlkfENMo4DdNuvGzwgpv2vSMU9MJ4TX4GwYJmNf/
7tozS0o9OIySdJ4zBHSe0zRu990XLosXneZUoqF1F1PgSPyW//RPbIKa1FWMUWqa
897q8Mv5wBM7tTCPX0/mblImEiNeeNYPoDFm53CxZMQTcuofzNI3MmuqD0yYQu6m
xaandjINPOE/R4ImqdAdnlF1vi4tEchQYJlPx/q1yXASLBiLVJ08KTtkRZTMs1RD
7j4BwEboyu0NgpkI7Zx6d44G3C24ojpsBb6MoJVW84TpYnkxJtlOQvPR3LWRZHSw
PT67vTKI6W5Wt+DA7ZtXCYn9ZR+6MzqaGF7FChCjIyYuD9zETBtGhnoywkhjpBKT
eYXMv+1QKmm1iuvdoHjNyKzeVadCU/8YYv6z2+akMfBjdNsDv0l1EYX+O+v2F0Ip
lp7q+LRTLy6TJOn0tGTKLXKTCSMyR9OMgAkkCwRkMbeEKXd3rSA57Qx7wekLbWvf
YhyFiK4nhqzI42QccE8T378ZfNrD4pnMAfGFlKrUeXzyfHk416IwGpcb38NXY/b0
AtWwBmZV9M302kBR8yeBbQvNBSIFBICv+R4LnFIY98Yo1UqViC/uqVA3v/nY705t
XV8ChGKkEUS7je/z934/91Wj55MG4WQMh7Sb4LyQyy0h+mSeJRiyDZfNxD0NpkK9
LTUbeFIjut0ERSuqcENmFFl4d9lvDjaA0VGpUoH4ylnmKm21J5ef/D/bJaLQvyVB
tSyu9Fmyhigyu0zODzJ4iNYj7fR1YRwZ5+L6NGYjM0hHUJXHy0NePrVOq2mRpGo3
GbW+96xoFJfosu7iM3hrCMAgTqbxPcMB1LAER7U+NlYo2zcl6kg9VeoW/ocCP/fu
UGAHBkdJfl1D92N4sG0cuB0gtT82xdkPgDcWOy+vYe6FQdbcxp346dA6QZaJ7Eg3
nC5dPOeYuJknoFKhC/4WI4AaE2zUj6azMbFOFTxpmYTIT8WLph1cMO122tjzgKsA
lwkF5XRlli/7sofRHxXzc37P5IcFVKJa6GOpoe4GAkvG/mJKZK9zmClopS1Glt5v
5ZxUUhqk1+idYWqM2iDzbC/prHNmbVGaDgwYLnrG9E5jZ6ltoR5MVbYgFPadhBZ6
00j1wmvOLKcBpVWLTDQIO3kH73zMvvsKV76D6kkYTRWQRMM25IZhxUDuEjrDFkgk
i1soDDSzZYCbSF0P2gs5aJNObFwa9WTP+VUO+0B3EM/xXy5uj0Ccfv+v3GNUBuZz
DvlCKDphpFhPyjLL7ddHhZZaE5SnYqnuc0jTYp1LlFNL88cJR0RKGutyg6CvXBkU
C0kaaxw2o9jRjwL3Fnxat2blLvJgV5eVayKIRGL1mxYmfMYNlLGdf6Tu7qAv/x03
DAuZsG9rVAyfFhxc/D5WDo6TnfYJITNulAJORGJuqbOzGOv/kVgk5e6BiHEzRAv6
s6RPKD/R6561j08wwiXWFLRfv9HX9Ay42jlOXZyiAVcvYr6AqFtTDNaCDao5fruV
qg5M4EKwVR0TWgikbwwwVKkGOM2uH7Ud/UI+SfBFIIJdykKxwEjEkhYb9CM8QfhQ
hejD0ehYaXIdVCLD5ZSGpxpSu421mjOXHqnPfb0A1Lz9IqfnPpIAHBPq2ERiVx00
gDtYNaNeU08+SjyKrmyuCaGtyKqHETcETQNrnLyL6foHbNIG/ggd2+gHFtqx7rwG
3W//M0AH5mJUp8aptvd+hl2veDcMtp3UgWNPlx4lrCrm7L20yHay6m4xClqf4/R3
m3em7U0nDoxEJLYYtJRib1Q8SZ/0m/5nkzlZKOaalLCSmnaBsqsT47v479YzDDnw
Gxf7BAIiosYsPEgFJ3TyOC02wdTNoDyQKNB/Aw5BXG+0+rwmH6wPUoQo2dBLfxMv
HdSYZvkLU/bR9V6/JI6t67R0dXa/w/gC3MHdpIxyTkousTfSAFzwNdczQ9f1CsL+
CTdEKGmF+tQ8G9klMRisX+5+quNgktO+3KZ51FgPy89PGl8vl5CquJ3wsD97RUvN
UvaLehypGU8jcH1uLOh+Z1UpwHyR9fiQ4+Go2AiSDehsbzh6yAh5bNSUWsm7yblT
JZ6Smroxvdc70t4zL27FM/N9v/7Gj7XRaacz4396MCQcnPWVZu9vYlvjIqTMIpbm
FtuSi1Ss8q2LXl/RiWUboz8AZ2Lr7aQkKG+taN/4eXU76gsQKF4WLt7+Z3/aN890
KAgF3/EWom69Isy7M79avJhr5fSZPHH37fHPgvMatM9xvmJnEg+l4yuXHOqFK/7g
Z5WdnPvsJFbqH8Nfyhj46s+VJzIPUlSx9+qojv8PxZxcaOAPPykgDHr7Zdww1Umh
mUQDosVmw6QuU//QPvLQZPQrOjUh3bt0Fmrd/iVClLCcuT1M3ZHRJVhV5zvh8B8b
OeNY6cId2y3d+KF5bZiJwMfiO+LgXLikxI9IyFPJ5ppchqr/2CPGvo6x89c3AbRJ
STysBzbfqIlB3+ob+MVxzfC3JcydcXZvikzdaX/rDY4BqCOHRMfgZvdphEwj2Fou
lo8Lv4BuBJua0AVP/dqbSKSvjos+Z0WHQP8YrGIeKN8u71Gkm3hMkM13rt03FLVY
fnz9BJ7wrZp/V584uIEq2m01IJw5UnCgKT3CUlIxOrYWIIdPpCybCc0KtvrIn3Tg
UOFWppow/F+XvgCK4Qy13zsxaEOVd3c0bWbeJyyrsZUjcSpMMu82sqg/cu9d8tj+
1nynxaTzNYLB+qlIPCCq0FbAjGeADDH6WbYnxRY0DE2OY3pHZPzkdV6blQXVN+9/
780Uj9F7C0L6IMHrQDwuFzwRc8Ir63Fot2PxeQGsNxckGXHBuwlNB/CAVOUxCoid
ZjprxgKj58hD4AqxeUt6PIFSPCul0xgoOBLDQHs33BrTPcK7VwN1YR+foLovWZFL
iyqUeUBYUD3lZDXgRzACV7fRZQXN3CpnNr56+NubE1LOgVPLDEbObgxd/wHK0bVl
nucYVspoNYZ49kEg7Ylc7d3WW6/KFB9k1+tU5UaWHfbMoLXWXmtudYtan8ijRe2j
bs9gbuAEtqN0JDojMrFgX1G6LUH8bhmMLcSFpeYnEQgduLv3wlDC0cPhfgSoHUAl
6AeOt7t6h1I9iWZgnwF1IcR49xnde765NsNg5A5ktVGGRk9fTWXmZaZbPCIA8+Lt
hTtkS12tY+SW8K/oq9mP5BU+GYKSqzGyDkoFn8zAn7ApEDXDi7HZa0B6BkLpU+ct
vP3CqBHuRvBDtb7s/7+1CSQHJeS+k7hOgN2KhIGJaO/Dw9ckBhExeR/eDtI1x8P2
1gp7apjlhpeTNr8OMamQRBNEy9e/fOk2xj6PfTuW5xTtCQrQ0e4dJDHKs3Vp2y9Z
orjVERw7TbAKUSDhke4BFPjgQ2K8ZyAo+bsRQUEa7j2jbXUoR/Zu7M3FkFFFgauz
NBSOY3xN3N6i5MH6MwJpzTVwGJfjfy+F3e4nFmnHX9O3Ctbij6vTMVieqaP6hW80
xzv/SapcBk14mnJK63JHlkE2RJq+RdM4WWf2qzgrgot0S5lPKIht6jVxSHt+gTbt
dY+eiAfpjB2k78UhS8+EIfvq+/R8VrbuOafR+Tuf8rKv8Sq1BZCeP29fTNjCkUJJ
T6GRvXSB2wMJagaf2W9lQ+GHbEDupuHF4tTSlsoXAF9Sl7+SGoZoZgi4W2zTPbmi
DtTSqVzjPFFCQbK4Jzbx+AmLzZZRuyWGmcPp+KrebjwmKXwLmN9JisThA159QxRo
r4VrLKUsIB8oFJi3PxhXX2G1TfktCvA8IPDwgCZOB7+5PMmfVzn/YC4o5pkRc9Fu
ZNKUuVF+FGgXNmCl3WlNq5L9KWIjnwxetovxNU1nABPoTvVLyT7+RPCuXSJBs+T1
5lXGHOaGRwHM6Rmj+t61Iv3RgNk4z+7qR40sHmSU8Ctb/quN02rh1DBhlnF7Hswr
ZSHACEErsQHW0UhUlyq8GVYAMHC7FkmM9Guit/7KqGtVdjYu6l/2bhuCjV3+NpHo
QZNjfwcOQK18RgxxeCOQ3Q1hk7uTaaZXHNnVXJ3j5C2Pqff2d/uJP8tcuo39qor0
ZjPKBF8vzESnQ39Wi/6tTY76ARxihN6XCx486lz7cHAARx3d+HAp04lsGwsLGQ5F
yNYENjyi7kYvNi/6Rcshluxx/EoAUOC8wS6yWZJO6V9xOX3W4a0hKtErv66dg5lJ
hDLlSTE0Ol17PQAzN04totPhvK7nMWySysX4mS9Ws5B6wv1S6txJ9OwCISETg8D/
alGw0fzH7oTyjNSXRWl7n0DH2rzDFARgnOl/l+6bDAwrg3ryu5HOpXTFqw/xMJZe
NaQ8Xu1l1k4/R7LtHtT9NWv/AaouBel63ZyKBKzf6GMGBDlw3aYtzxNlkz7HBval
fTlkc05ZwG45YomOto6q3pf4PgacfdlrJF/5K4nKdPv8TTAE1PlwwB+qhCyl+/sY
lvRLMUzJvqKEUTA8jk4awLGGd6P9Jo41XXgL2HY3q1M+cQGr7iYxBJncUnOV3fI1
idhwZFaPSg818gf94vA2Dd9XplLSgPKZ6cce/P+6vfPBb1Sc0asPlYDGAFkhCah1
ivWmnH5dloJBVMYx2tEl1X4SW+7QEY+VmdGloxBrNaRmWhd6ybagy4pdcUyDugUq
OYfkPbPTjQlZy8cuWCA46gDgXuUWtBtH3ohIWgSr3ayWigB65kvbjwMXyJ3+lpan
zoqEf0yYnaWx1uQDQdFqb8qULrCB+wBq1zcGcRKBF/jF0P7VZBNTQk9D34Z8rfU3
nNmxWCg/zkgeVey6rjeqH7ogUo8l1K8JLNOoDYkgKLXjK7KYngWz1TkJRQZHyM42
y51QQ8/w3jilGCKc6tPx2nHvNLDmnC5qPt66B7XRDb8avrMUT1qNllc0Oedv3Sdv
ij3wTYngIzZ7KZJY0IXAR6rCMGR9T+KREgKWXmvABswlre4uiTHcINOYN9jc7H9y
XJNe8COhRf/3tNMAu6t5GLIyLWZf4LogfbISD48LRhjb1Xdm3MYbs0I4ICDrr2Jf
XoChaEJCepldagn7gS0gaqC2t3zK+fGE3yCfMlMs2yhNerscPmF6Q3LioOFB2Lr+
7GpSWe4LCD5WGTFALtsc33lsoPZy17JPouQNwWaxpeLn8lihHvsR+DBp8plfaDA5
Zbl6z8aNCxm2taMOd1Mgm2MKA61D/HpSZkWw0MKLmEzajlSQnmb6junQhY0rDVq4
BUdKzkov9a0hsrMUSGzTUVGj/e8aCQTdI6kT+mG7hO5/E/bQKlaE+4LlQoRGpaih
EwOiQfCgXr8BsG+n6nZge9aAeZX7JPfOwOCZqqQ+enW9dv0zK5WbEuyG55yFi+1y
Rvbr0OarzrwALOdTlerzeNZ3GERe5ZPPJZPYUX7HhUkAxWqi4fFU7EeSY9Vv1rJ+
af2W0CJIL0T7PXFs9O6GEdGXJmC0X+ZNVXZluCSuJxmuo8gP+KjfaqE3k6DLiFu8
NFoMs6cPNbUMAsDOYV7Hzg5VV2WB32WcBMXkp3CTQqbU1i3yRL9hhB0SZIN3GTYz
YcAsR0SQKVgVrOXPZXjMMwtPHDg6BeIAHHzqErABi6jsWe6O4uEtiKolZyjiAeZ/
ie0FfupjotWOdRWZGVbxRYSVXX+2puMB89V1ljzc+mUtws9t4z/SkExC362LFNSz
8Xb+5322aYkErbDZEYGiXUqmCy+NGhcDBlMELtU1ij4k4YAsAevjKSiSVVd2c+7g
ogRo4Y4m/XhZSBSQp9/W/ctSzqX14JjPNY7fFPU9fCCki4mh8TIqoRV3wGV9eCjm
TQ1/U/h0Fj3i42s7eTCBNOUqTzHgENux0qsK7b713PNGGIRpmhDAh44NHmJTKgpX
WYFdRMhg0CmZCF/KgbXxN2DnZ91bICTf8VPW34S1AcK4YgMwlcvjmaxfoFdjU0ju
IXgdAaI8zBBZDDr4On91HSF4fLewjaeNH8TeZHtBN/T50clooGfjQdRg04dSLEf8
Vc856QLZMvmR4qX3CGkE6WiCUQtbBuIP7go+KyugaLBVNr9aFqfqDJccKlh5qVDu
/qYNM9sBJSC6a3O+bshrQv/NUW1osVvmBx97Aqa9b6agU0FwnKdoNc4V8c4xo1F/
D7xMBjEzxkndDPY8ILdbI8GvSJP4Ci0+d1viyNHtuKe82rSePa3Oz0ENqpoVKsms
lOGMG0oLjOLQHwtiRs3yvE112ocfBHEQAMRCcp/tZ7CIdTXGlAYJUo8tuxjLYvxL
y18PgZAiGDorsY6X9j2Ca/r2w0teXAOLMppFdmCGQ3JuauBCtluw+zLAx8FguhIG
a4NTVHrEd37XZyuecUhnZhmLbUIQaU3g8bgVCN+UD+8k4h+R5O6e48No35w+oa/X
xw/7YiKgiemXijC9Mdcz515e9t6nuQeTKvo0vHQ9rtWqSZ0P59FMY36/B/nXml71
WPWbmH6S0m7PxkTy8uuunCXhBdzRR1VXOqey0ZTpZbt0vhAoi1115FGxJtGu1fQ1
MQ/NdHtv6fzA6KkBh6S7Mwl+94C257hgcYPo0GgC2bFvIv6dAApvFFVGzvOgp8Ly
ZiU8ySnZolbztiecAf/0mdQ5yo3INS9ru8qHybQujAsPJzx9hAT/aUGpOXXE+JfX
exzxslg7Je/YhdPrSZBMfIRAJDoXUqU6zh2pJ/cpRH2LrjqXneAtqqLMxNGYHuqZ
NMbcx1CikW9IpUXdEvIBg5vLQ6/k1nhOYdBGBCJNpwRlD0Rb4NN30NIbto42ZMrQ
qUUXc8VJkgPsgajHj4fIiJBxkFlx2QDg46hwwsQssGbE9S+Bt5ypihuyXOtYvhqM
BW8dWaP71zZS+Dg1T2Gutc1sZu8U/kckmvIneId9DZ3jMWN9xd5Bgq5oAQDBV6dX
OS7IlY83h5fB7IYhpeap/A9gszLFawbY5KUPC/MiNWSVaXoe4uMhOu22B7fKKMVE
+Ua8YSBYbZTKLQS6DqXVpaLZQs6JSuzFibnkAd/4hrMvBQKP6sbUo2S7ELWZ/nsL
NrIMrcTvVmkSVYOMerZssQTiNp0M1uZTexNxXKUc1x/WyIUvc1ncggaTaSPLPPi/
Jo7DWmQ46NZi1tmLjR0P+XnpcjbdKBmlGlknHhLTmowMFOvkZZxJEmuJbdyH3IF0
Mtfyp2L2lCwL9OI8esL5zb0fGsIfw+0dWjT26PtmWgzwMjtK/vhXm/Mv+LD4fXDO
bgfSdVPbAFQjEoT4H1/ACHsZuKymMEMdWajJVrx3Uz9uzRsxkvNBCm/2HTjwQSl9
pBB86c5uLotS0CvNr4Dxw/ZvcUioMoucCIn+epOwXs+fO2YYzssq1yjdfn8VpxkA
X68H5xuXad9I2x+5gnoZi7gCZLkq4w4ylHDSBzBabduVn7CPUWvXhQOSHwQ17Zru
tGFrqogqlPuhxrvU56WPsU/8AgSbKlMnGxZRspZYzF5/dXnEvSSySoPFYarHovfA
Afiv059dvLKDksD6qhPWNeuC7EireH6QlTwuYGpRdIsUubhb8FWdLgNmMbw+FR3+
bzEF6isDNqqFplIBkFP+TW9owuEJx9qkDPcQ40lKUdzIhDcRwYGHeRSLqo9zYriu
0Q4PKkwQ54h+JFjG6jUCqy1JIsRwNXpAIIo8vsgriOt/SVPhEQHlC7JmcDNnEyLm
EwMawDBP10KPi+r94cGoxAiKilTxwDA0mrNsTMFe+YUvlneiv+apkQhK7eBg9ejl
FCqwN+rnAIaeGGYeZbAY0+/RoaIwpJC1jtBSxELWiKR9dy8DNBysDKCxrwT9ZYQL
qlmzh4Eidi620LaWbzdILH612Lw+SnTSVVu8ENjba9QGa4ug0Tt3ah5YVvN0qHFi
I68NqfYOZs9LMPD4eXWlnvbZKhH1E1oeqoIfe2XMnQ0kUAjFHtCQMyfqoelHW90a
qVSjPwrO+V8e+/Ke2+yu82Q5EdupHsRwvCq6p+vXGprJzwmCdXMzfo+ligm4bMju
WfLXVYdNmnW29chVJi3hW/ulhAJtM+4ueAwMfjxlnKltCcLeaSkbSFHqu4R8577I
PHAYbHYvL426iUshCPaLbHNWCIB2ypfGRtNxq0N8b00hWKHIlHmdZ5reLnurh7hh
Iarcovet9mYERCtnKLsXL4AjyRtW4gnA+n+/d7H1ad8WmG3ea2nZN3NG7pJFAhh7
KBarxMWAOg+BLN+xhKDOUesHVbmBxQY+B7vhUUQuxpcPt3DRMKghWwRV4qK1lr9/
TTugGpCY0L/jcAi+knBNSFwDQNWqLDOIFPsvOUySdQMuouv0L3U874XkWZAFg46p
JeQzBzWHom5eZCGqbjqS7gYSiZFEgfBUiIcBECVTXo4Xqw3C5G5ONQJ8yje82Bcq
levRNnjajspSJQd1SAXiLhLlm+5cun1D5/laoIAYGW0DOKL2Fhog+RISugumfY2R
OaPlcG1+U8tVRqP4RQPyIRNIxJP063DschYj1eaSCgYTjrutVzFrVG7J7CnR4VBb
tMshizfvaXzcvyKyjq1FikQQI3uQUYeUXQmsZQYVW7KxUo/lwhFhqU8ikg68Kaju
yfBxsjvSn9k3uFzP2yGsUvNKSJGZ1DDL5d6oC1TEetuRFuLvXfCQhJTB46KMMG+i
MOszsNBC7/gOGuSZxVR2QMnEkmU+JRmSFnrnih2k9JGmkl9a5nK+PLRsX6AnzL1/
yOZclh7hzlQyRVifTyAGoV7dGl6xvoAF5tpifTFEgYajE1uWcGorqI7l4KwXktlH
QMYZWsoT3wODsFZz9YzAyvX1GM5xTVyqtrfTDVdB9a9MH5kzRjjDIxDOQNw8Tj/G
ukXMrFcOsESkVmu2WN9JMbupwk3fo87GonsQMry2TjVZg9H8127OUoX42qo5scFP
Jg5WOlL9qnk1/ui9CvYyKVRDlfT1rVHCIdl4iYyRzLBN/6Cf7/GGmG+OCcMf6mFP
/afXyR9oxjFHQbZzHpRGy1lsm38p2ZS8jd8FvjC+a/osEAWPmDluAHhc6LhJWwsi
4kq/FwZOhD3uN0VwSI/sNbNqo82Rg1cnfMz3PA4mVJjijy8P4+3Bb+rVfv/FXktD
QC+TvaTsAdxIgs3IHPUdCM36k3t/DLOsQxEhwpr6Cp+u5zgVHxCpoDpIxOosN4e9
IcSmJnLe+7TOxDcwUCNq9NIuf+r5l3zntpJ2jj1XpxonF9EWGitAOE7LfCArq85E
DIfRw2R9zKxjcL9b+3UgcbagojCrWR+52Q48BKQvbGNlQBCOPp0c3L0s5ph4aD6r
ki58GwP+r5rcLmu2p6k4cpXO/pDro+r2cANDOBGpkKGULZS3wVHXvDWZi5TPRbV8
xKNANkQHdRT31z5S+nMW0R8HfZVsxTtAtxOtukZYsRPMDuZV/y6NcksIVPo68trU
Pfq7XHMJe3T0lo3nYkgauv4W8ufDEEcGuUYNHJfF7OiylDpih6t6/F+M2YQZ9KZZ
HYjCDOHmp8dwYNTm6dGn4+NmoMOjRoTAOQMdtrNdPpgbosmqj6xf4Gwnp8iES23X
vUdLK3MugLoBsLZgM/HRIS0NTsoTeZsKT3sOWCFnIOvkb8++Y56Nd7rsJVMHWjX8
yhlc75SVI78dnbM1rOfmzmgi8romOL2mRHZt04VxHsxdCMhFr88Oci8Bk7QuM6Au
+4QRNQuc1cPI+rSgyZOqNQCK9Wz1yXBZVVhotIJlbDaQh1rWWzpZMaRWNfVUc4J2
Ue7BZAy40z0whvDzkyxcPr8GrPNfM0fTI5dYRm2Wzb0EfKHO9wTrJHbi7jN82/3A
9LEKPboSLBJ0zkJia5oeeZjBfS5eOQtqSns8OMicJvhPU/vbunaKStJ+7tW25SeD
ztFlycp/AXtzMFazd8sIQpqTsfKezDDRUwP0pZDqQNMXpPAQizjF/I9p9ydKs/5d
c2hlZZEMyo4vLuQ4qxy60jVdNt1rBlclmsQ4C81RTzxSu+XiAlKVYoo+8Od2QvHU
MkfVgSRV/3G2DMUojRbcSWoJMoxjkWgWyBwlBBFFfnuVHUiehKJkjycvtrWUoZeL
6Q/nAMUmCll9AvzAwuuUdv+gB/Zi/i70ACT70HvXROJ8EJ47GdrWdWME9B2Somy2
1S1kEo5kQVQuTc0DDV4R3JfTeUUVre0aqNBzTRp2Jqx7uTH3U6UUAlP0K9ku9kcV
biTTlvON3OT//xZCHb2Su3lRHl3zTUniD67a04Q91Yw8v9HKqMzdLb+7pC4RWd60
B8EUB+rs3uX3IYYpGejLYT5ZwBzZmrDXYBov7u/KQWBhMJMmMXY6HXJ9pXa2eGIN
/PWWg43MfvKqORI4IEfjwOhv743U9O67ftgtIpD0e79cZvDCVS4CzjbBvlRk2mH2
sXoOfQNGmf1FlWK1SXFgMo74ifCiddtDjWFC32zZKjwWG8A6UWZlvNFf07yXTTZ3
VTrvJy54edvIKobluXZbSbXzGNrnZeuwuz5URfvNQWGKi/LFicOptMNcSXo6xS4A
qO/fv4Smr2tM+yBnVWw9fJSUK2xs12y5E2atnwOK0IXR1q9W++vB0UqdSA0XJAtz
gVTH6cmRSB571EMpSo3JBTV7bAGarUhN+4O10zmn2mp7zRUPVYmgVkJDPoOklUAq
UHPFrBUwC9PTbMhTvJshX6h7E92skqynctL6725DTOmpEndJ/JRhDt7DdeENZMuj
W4mANEucDpN5K9exveN3GVo89Ma4Mb4QOWGhRWAah6yv+bggDLS1Z02BjoBrzF4F
+jKgEt27KSiLEqV+HRRAlpXP+CQpeJjWgY6O2ZKI7skN6gWXAjMweA69FrTyZeAC
2LMfy87Q4bIKJVYKtsA4gkKncmACXzUPpA2cf65zVcC5GrvKZxYxcLNEeXxZk7LW
tmy6FLMTesGGPBSKypQQ8CzJLEWyCOgf69WVp7mqXIVVT6THhD23fpNXQPLYwOCU
AA2gNaRykuki1WP0pK0mPdJeAV6xG3YHQKC5F4adWoJ/0WMUfCktoyQcNKBA/q5X
atRYJsHWmlQi3+OaB/RHqby98OxPqRnfITyQHaf5Okyh/o3pWdWueLneheJvTlW4
pCaYHAv0LqMkZOMnzemfJ0W7tKPwrFpH8BrINES8vWypt5cKs8RX/ifw6bk2NJK2
eG5GaYlzh5RVH2M8iDNQvVj0RpO/AbsoBG54K6AYgspI2NZ++BBOtOM4Dn5HPRCs
PntptuOXp9nwGOQ1jxdnW3G+IPmqCT0Sl3oGQzhEtOy2B9p++HVot6BvpdwG7tcS
6/Vl0IsAm8blbHxCtRRlTCSWcFiqtpXEMAurEWwQuC/EdSY7Ae4GYw1de/0kGE/a
`pragma protect end_protected

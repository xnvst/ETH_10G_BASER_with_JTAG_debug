��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO���R��gɯ�Efn�L���\k�f� y��������i������	Y�'6�hMi�ꤳ��?!�mi@����Ur�/K[1�I���3�6:��L��И`+by���G�R42�`��:b,]���*�u7[0 ����"_
�YA���j}&�nH6��=�=����W�����
"~�{������ϊ�"aR<��^��9�L-bI?���¶�9(� �5_�q��5��Ӥ�W�'j|fk���P���D#3Xt/������(W���&x�e����}xY��aV�G�_�4�|?Q�.N�� �'L5��Ǭ4JA�P��P�6��n~!t6��>W�iD�`�Z�r�LX?c6���wH�iZ]���
t�5 �(�Q��$��9S@�#���HTpM� f#닸`ҏ�tA����d�SL>�	��`PSj<�	�j��6C ���r:Dc۳�t lY1�~����W�:dh�N4P�N��oz` ˩	��%��#�s:xެ���]\� lU�L��vdV�KB�`z���8�y���a^ �Tq3i��5<S�it���Ĥ��"o �I��@�D��BMSh��9LG-������1�zEH��������}��YEĜ]�FT�ˋ>ʥ	1�U��$�������v�W���<�%}q<���}l��M��t�1a�c��E��_��s۲I�*5�j2*F���gp4G�l��c�- ۵ ����En��N[��&Lan�O\���ܜb �(�8��]Ԋ.���!��1���ZX��mJJ�;��n�����ǅ�����^=����`�p�'�E��������������-�Zԯ�)uV�������'�x���ɨ�D�� aN4bB�1����v !TB}�Ց#`>�Uۉ��H����qw%��P��x^X^����Z9��[t��^����?��%��e��H�1����k�<"Ż4��2�V�tyo��0�H�ȴd�]�ݙ��M͊mŭ�^W���/�X��z�Bq��,w?��*�T���m'��鼦�q|�	E�{�N_��sK������@)���6�}{�+�@��'>�%-��FR�[��{X����^�͕���T�2�j	�1�L�L�0�*T��(=�RR
��)��t��m`ü��IU��]����ռ��e�RLH��te�+aeI�Z��44=�s_�ij��gp�x�շ��o�J�(�y���,��T=��q}��S�X.M =�+��5���	.�r�x��M�:��э��6����G>�#�D_?��#�����I�$F�V�i��=�j�Q�Y;s��E�E�Bn��;R�?�R\l��2�t�2Lذ�
�u�"b��c2�&v��a�yH��k��%��a�	㌋�֌��Ӭ��b_�Z�"�5��O�_0�\<��t�%�A��g��夁 �;����(���iПԛs���&�%���D��t��6�$g�7��,�Q�͍��WX����z�;��}��A�)����K6�o񒧘�����&���F��_��x����Ħ�����޹�0���Y������*�I��㣹���D�lt��E:����J}���Sq���SH�V��2.�@-��Q��y��:*�]��ߩ�Ԩ��$��q'�h�rȡ�jČ���͕_d 2�p�G������n
9��o@��i��,�E���~2*ҳՋ�';8ݡ������ �Dj��`N(���=/(.F̣�oWF��pG4�u�p}*C8���%SD�i5�y583�
\�Y�=�[�b4�o�wE7�L�ǀ���ⷛy�W��[�ʱ�u�pSĝ���A�Z����,�ߓ�'�T��IV6b��v�>6nݑ+5*ĬF�y�<�I�M�)�B��'A�A��H��7�ŭp2C<:
x����lg�$��9־s+�����O��_�vǊ@�uR5$0?��'L]P���f�k �/��&.��N}���/����1[����F�u�����%=�i�PLA'oW��Ro?Y����n�xJ���h�:�d����S��<[l/���A��'��a�9ۈ�Uј.#2�̵�ܘʆP�M�$�(��(!�*Q$�.B�CH�R�pt:m�&��D���o�4���M�)��86���d�s;q�n�=�E)�|��E��2N���B"#��I�[�E6�bo4�å32�Q9������D�ӢNq��j����k[A�ʼ��?��
��o�P�~���'�P�,/l,$��y@�r�#�!-[���a�gz�<���$�O=��@�;^��F���������_�g",�c)����9��F`[T�ҞŪ��k� j�wE8��2v[7[�+x�hDJ-�B���{G7q��խ*JH��CR%f~�Q	�P��Yƫ<���@P
��fs���1u�C!�[�w�ظs����j.0�0�r�5q�x�@C7Pf��Y��.<k�9���|܆�-]	~��J8ש5.�Mm�S�i����H9 +KE~�	 P��;�ğ^N%�̀nޞ��NPxb�e�.ƣ��j��#"=�_o���;0��O@BI��1q�}f&����8nO����0'Ǚ&f̲���J��ݡ�ސ�r��a�y�*P>~��9rH�e��v��{8�_jaj� �2/����|��2����Y4��c�6��v��  �4�-\�E}��V�>{*e?�o]�Q��A��eC<�Gd;�d�+b�XS:�x)b��i���<_g��o	m5��xW?�x���?�X��Z�uu�8K\Af+� ��C����祈d�C������U���]�����QW#ujM\�(b�X�n�m͚�V9����,e��G�4�$f����x�×���k&�#��	��W*��v�vV�J�Bn%v ��7f�L���\��h'3ܒ$�31)����)���2��HU����3%��\�o��㐃�>���3����cD�0+5t)
���S�����A:H��c����ξ�rƬ���r������@��}��c4{S����?��e6񷃡w7#O�*��ۍ����V�d�R��IY�-^ǧ��pV9K4�M�$W�,�h�]e�jus��4��M����91g��e$�;�� )[��@d����}}�lb%itM�d�Nu��jc�	x�`��R�d���Ά"_��`�qK^6��/I�BH����E���W���+��	����qD73�.
Z �fX��"D�e�I�Zf��)��"�&�H0YtI~۴W��Z�$_&��d�sX__�! �賠?i�� 0�܇�0Q���89�r�w^2,n29���J_T�2��3-�Z�,�LR�l:��73OX� ��&�( M��W��U��"��z�#�Oڊ�P�䘇����B�"7"����
// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:28 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MxPOo1TysV8ro3WCgr9w5Ebv4XDW983En/WICfzf9bNqt4fLs9UZvn/kjwJllHBO
ApYbOM0pBceXv8JLWe8FpmhH1n0vCkyNrbS/qrCLegk6xn/dSAaT6iFSLirqMTzs
fpT5SljwudYEu8l3ghBewcNX0zdC3uFUPHqlmma7dk8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 104832)
YjdRdd4rdKybfwD/0Fje5eUDcv+UtAn82nfEZT9WBW/3L8lSCO3g1Xnlnv+HWuDS
THEpt1dA/5BN10Za7DvWkz7zDGZoaXtJC+hOgBFxj5PA/A45tAbaU1Csx3u5s62Z
bUxTyq3fr0V+gFX+t4fKbWiwDo50hSC1GmsojuIUkXpuwOXU+CogKt6kBBM6eIpc
5Ur8qahr3vYX9vTl3c6kFtZpFvWDykbJLqjWLOJtRG6ZHIGm8gnbNDz/vdq+9VmR
8WwZs9DLbqSe8+fentHOGfasa0M22Jwy8uzq7GynWEfoJzrNBt7tBBkAzqy/t503
HxzkEHyQ3dP57lDm7ApaXB7r9IsSyYbyDv2IzU9pCkLXPtRcZcASNBTSuomj3v8q
xSPV0zAiZBHgI0/mB4BUbB9Lhf692k3W6VeTixNwUC88VR49hebT6l1Zxsp8JTih
KMmzlhlvniesCcMah4IO0NfiWPFFmjC52fH/G3h6QekDO3ce8lWZYFHCsH7c7Rey
pDxqFchzSo9NiiE9WtTqJsFIrPfpBvTf8SCbwt9aHz2wOCmVr1lWZu+VUwsFAydL
un5kjavOvGY9iMSIesGG+f0MnUhhCquNOnMc2G8O0RS/Yr7D4ZV9JuD+rH7wOiDr
9K0ksNwl9hkxEDFkoR347SVT98VCFlka/00jJXOpvMtcN7gEr4bJnKip6amrwTWz
T91m/dFzcgsazWhQNjOMhYSZlrwQWVoqNVAIBxXKUOdTCfxqyQ9+QvDd+ESo407E
RLh+JoHIxRC+3OP5hD3HlDj7r5AOvjpByMPMpEXiqV0aVaVfMcZxGlFhk5kWYgtO
AxlxzoMJ4Ei+iLIafRF5VdLPMo/KsvwwPc6qWQIhVs94OLiObl6ORKqx/wGVOUvl
b8A2RcSMKcseP4Ly4QeLfi3iNPrkDGSLq07xDxqnWgIZFNzvMV+owkxciY0WVv96
5uGVjZU0m2vRDfwwozSl8r6kPKMANl6Cp8n4mr1Vis4cBQbVJa7TiDTzsp1n9pFj
5hsqnwNGtpvzqSY5rMtI4D1q2504uJ9rxxqXEcWKlOU1vNIDDRgdHIfVcXRkLErh
T9rmcD9vUpDqGmjMD0+7NWUKivq05GszRdjuHrDVs8j/EusHscdeg5JmMFiTLnDn
CIK9SRo2oJjdfdxY0zKENwAuC3pxXcfbZp5CVXXtPh3zGrOmWyF3AFCt6seRIwwI
xcM1LKQy1A7XmOGRQ0OSTHtlYBIU3dCb2YSRMlq4iKURvxda281wXGjTfbAW6kzi
TzZT2UfzJBksJCKYr0PbxLKHFBcKn/mkc7yW72w/qKhTmNK/CnvIERzo3u4pDzDx
kG9/kjBBHHvntHoKleKywb7vB4vULrEsnP6HBDnc/TXYU+OnlqlgoCDRhYutNkv3
hSbKYBafJHsgaMK8f6e7pUAabm+w4tP0ugNxKmzY33bEJlqYq4PWwRLlkKCPSml8
/9mdY1hUE+WC/a7sqd7VSw3OlAjmCmh4TcoMDz6Pz/ABrimdX/O8mQwAL/Uk/rCj
BqQx1f2yvU3K6Cqm8CJtNM3LuqC5BEjlJh4pbHH0q1iHlSeP0Tfyw7cHZ+Qi8qLo
VGnvbU2B6F6H8ClsfLMDKzt+zXhET6n52bPTNxYA+HKZRms9X82OD0nS45JUtiGJ
slox8YBaNVZDkfHRHfowjgrTxVFO+AKoXWeGYN3ZSeRB6w9e/O14G+JbRdzyLtlV
HDLqfqz6i7pMByJ8T4KXf479brkI+SvUaRRMo/vvmsznkhTsHCXmSeu/7Wy2Vm/q
2nqg02C4KkXhNR3S5FZ/KSqi6g6qMYQrFQ2wQr7YUZhjn1ugGN0PXV9iP2tedpLy
1wjXK77ZXw9Pn+7xD61Kw0DZJqN4ZX7HvAqj3/VB6zT1bpn5cOdY96FZYkJ+brj9
MJeWT/e9A46FR3AqQONV+DBv2mZZGobl5yKfhC1Xa1eLA3YcLd7lufb89Qbfbhsy
zEfaTltKmD/Ga3KW7QBuLAzwEHTKcDRpBBC1gL0p6SbVeoHKbTuiDL3ljfXg+BZu
tQTXv6FW6dtCUnbPWx/hZ689guzDqkylQg2NfBcMTExv3ZTbxT+aOpo461GjGGrI
6n6IZwkc2WH91OQba6l++pZbG0qXuMVeglDPeiA95puwiHh96gvxjRrZ/l2/9Xjw
2yKaZADK3ydIbLUIFFkxo/CQ5e9Sd2Vi4QnMsh7yaXVLw8rLs+MARt5GkdfdK8Zn
Sdpvib3ev+ka9Up//iQzjpkBvmWcMvsfM98xbKEY7OrmiULEnczPE+hLsQKz27ts
iAu/vF8b+7Fw0FXWv8rlcF/3wwREiuIXmkLXN8PxmBf1jDe+iAOcxqSUvn8YSg32
KtIviuSKzG/3dVMXaCzX5honD0M/jmb6smIHBnGwA/qLsc9XBcy/3EzJ/Nc3d0zk
zmYreyKpD/jHOR/2WSGmtjAoj33iGB9MacIxROMykyUVX/FeznH1u3DTlD5vGN4w
VBCFoSLjyc44vesl5FDmwaQIgMqyML0ZX47yf8PevmX7IT2SERuBTYaMjsxzFGM8
HIccDxSY7kuHrILyPcH+OiBJQrQ9bj7VfCAPQbPRqN8VnAe2mWSm7hbuFOXi3QDr
s2AdceluaZ7jxIJpCRKTwQflf64eJBZGMCpA4a8n13e6FUylaCFaWRn1dnImgcRw
iItsQo/iyswH8EmJXBnw7TLuTZBr+QCYDdCivEWbelx2q4247Hv7WWtOcIHTJfGL
+UJkTU2axljjgF1deM7ZLQ8AmRT7CxZxfZdIsLnUS4s0PrNv4oxuQ5XdQDxGuxNE
Jx+SO+o51Dp7OpDYM9nR8VPNaP57jF7ao+DsbZEPm2Wxea5BOX3gZKNQUygApIiH
PLGgYAj1SLz9J1eQoPM+rSNkjSmN/xuq8ZABP8KZM0QnfEwYrHjwzxKm2DNxC3S7
oMhoqZ+eAsB0S/gNHxuNfp0GzhNtEyeg4MYGXC5jIYl3/8189d1eKW9YuBh0rm7d
4G0FUTpndCTR8I/tf/wpQVDc4vRWr5ajqQXO77gLJ2S8r4pO5na3b4eEeUFt2YUP
iUSm1Z29LOUXyWJMba7tw634NkRR6cCqYfySyPvrYuvRGNG7yIIHLnYy+vg3ZgY6
4lQBGnyA0YvoBHsOnYyKpZ0+x++h94yqh9XSMsAXiDW4RqfyJIdRICTJPl+dTCai
CArpmPjZQCIOuw7EN2tLbdtsmQUmXYzinPlZbWUyAl8+McQPdp7KP2mVpJE0WffL
RBaXMI7IuPMIE44cJVC22F1D6X+i1tD5fT5bxTUlNgQzIZsVq6kLhTG/yMvR1kNg
HAX1NEOjqgcmfm6mE7IbMYZ8985yazG+dRZio+r5eif1akYEdzwQxjXf95LQ/YpX
J9squbnuZkPlgdHBdIE/kMX7ED2GB4e75WCiMS8ErGhy4grgYV4QnWDpTDBT3WCP
mgN3kYuBw8l+6AVQ3ycu6RPlL+/GzidRG0+AqkN8qLopxG1cVQ4MgXdoeEPMKMfJ
Dv3DPGhLqrNSutHDxMFJ9Ui3Yrt1EYgpRdTuHSaXjhAcIaat4Zoth/oeXogpU23o
joLgp5GGp4XPeHqol12wRyHsmXqRF/afkugkv7t4WbsjIzf0zMJygkZgbbdMPrFD
PI12xlhaztKQZtmY0Qqa2nfBYb/TFqSyrN9DnTpbnP3VAVdT442uvdvNI1b6ueY7
8dR9R+D0TD+wcsS5OX9/rduelCEKilnKgZQZaSn8bZgYSmvsp/xXSSVvA344P8fh
WHX6bzQ+j/GGa4iq2I4hTXPpkK80bcdRCdxlcJ5JA0qYeCIb55vs7lMSFsZxtZtp
eaS9kQVstcrmj10xJzzETbUuQFk+lXpynzk5HVMQpVqtFXpdkuGyCZ04MKJ6S2QT
TLuoq2m+CifVq1Igidb8Tg82UwH0NG3Z0GVOJreCt1rsoOnBBzGNvNYnE0HmPIS1
rrlTvB/aEQESSLbVvw5/u2SkkjJ07HYryOp0JIvtreBmC3W2lJjdrD0AW23CK4rg
VL6dTKW6e4XkCLkEpORuLvHQPI1DGWqpqudrfH0h2Ca5vVJm5Md4vpFQzetPv7dl
IVO5py8TedlaEZevqBjWpMUPPJu1jxrLoyOWd13nZN0Iq1r43ZUsavJf7/W8EP/C
HGgkHy+mtH/VwrZmTe05GY+FYwkTG0r984/sEj94vFsfkoqe8aO6Rld9QnGxeomH
X/jQxsccAgCfn8nNCOC+bZOkwjQMrgyOI1gTEbNiyib6eFGGeOUoJKcV0YRKYtud
FLWKmNtcDfxjAPTIvM8zPPD35Ew0RGY1fp4fxSo8F664hnJ0/+uje09E+TWLvCri
lsCnZnh2Z6M70FOdJs3W3QOAK5ndijdfpocL3hU5PzXUx9E/+yLqKHudMPoJ21Lz
eJjU+Arz+TvdU2AltH9Coak74R4AZkRjWtzi6nVeQJehS7/Yk8xHneKPnmaRgnKE
+tyFpNSinD0HS1/SKc1NQnB9PTOfsApPzEOM9NeIjwfpBQBjCw9TZncZDRS68+Pk
zuQ0vGyc0RKmv9Ocp8x/eypuTZSkVm36Lgs1VihlgxgB8GGOArXkk50HCRpxgcmN
R6oJHcpMxcGqX6i6YQj4uEnBEVCadflH4AHgx2Pulx9I1A1HalS6vk+SBGODnVgT
jpJRSB/NIQbMfYIi7rIiTMqlN+L0Zd8KbPBMfztDsTP6tdMtcG9XI3atWQoyagQy
rLI6+tZ88p20DRdAv6FZxwyso9OMKwO6ZBA5itBBsHKxN1zpv1Yy1VRX1MQUvmc7
57QEgbTL+y2FCJepU8H1zJ6Q/Fn06MG7Eu0AJrET/ftEHccZYENYaYqzZBdbyPwB
tu4fCfOVR+tRjkZJlwDcrgE7hpxxfaB59Ry3qa+KKTyyZ6zqfs5xvNYYRbeMd6kS
VyDwfUFk1LDcHTkTbXHu2GANgKdOG1TimOeLQxVvJAmlyGPMPX2rG/1UqmzhLQe4
wV/jMvwLO/6dwSbfok0xebAkKrDjW3zBGhzCBFcHkNtvI15NFtqA1exbOUT855Bq
/oybC0Z1+WTGJo4OHSs356pp8V4AO9Wm1hsPwswE4Q3bCjvUQcnECwTryEFVfKF4
HP0s4jZxrVtnUGyaocy2fXHMnAAVW4mkae49ZC4wrOMuU9h8IvLdLcZYH0SFuYZC
bhelTwT4QNf/vEj6oYXAFIY7Z/3lgfwWxwsvYyQXNa5grQXwRjx5af9Ig6bjF059
mOtbb1bBfXfa3HrHP8YlpH5wW2D+qF/D6lKmkmEzLvE0f0CA+4u9gO8luFfTLFJE
e+IF0el2GEofD//uh43wYW+pOl+XW5kNiOVl8VBXCwtDX+rKgU60K0uDnh6a8D/0
yuZhoV+pwGN4bzm/v+ALAVDZh8YwW2xOup2/m+10d4vPwZBW12uzD6nnilr/kKzv
uUz2wOp/0d/xUJTBSffV55dqC95KV7fOu/MVYAmWUQdTFc5lg0+clPIknIg9VWLr
aBZCynVuKihnKIpk9qvi83Ns3w459xgtIwoZQB8Ab/XwVYZazz4EGeDScU8YOLmH
UHf2olnXPeI/145edNoQ8VR3TjL+f0sbAReAV2qK7H4j6P72cupplIGkPO8SQZtb
DXwAIusRhdfkoU9XaXfx+VhETdEownm4iZ8smfA/bhYKFaIOPJSmtjQ4Te5gy71K
gv2S2T/xzKmpEpH2JsmnZRmgzPHOg9bvIXfrB2hCmhbA63rVEYyfgjjy/idOcRdE
YtwI7YyB52fSu7s/axOmJlwHEshvLP8c+5ZubIWSbv+jqd0KBVFz1CiOXaRjnv/2
oBVvMENvLeHMgkdVOnFxvYglF1AZnlxsx7j1zPmKmTVzBlvcXeSHtBRVr/tQZX/h
bMW4pVyLVM4MWlz8V+hL8WA8w+DkQ+uY8pCmE3sZr6giNIHYytvoveoQvhlC2pVH
dYsJhQGuw0omb3nMlKdpbla9dGWZjNzWEhchpKqcNlJCKoRoboVT7Tx121pby9th
AyFCjYBy2tciNbaOCmXyJXhaKbzRJMxvOmw4nAxWdLRqVYfLlAfsl2FSyiGDK7nd
oIKL6gGVQbA/XT+QufXdZIoxpwb0bo9JGqDAnxjqsORlujKsqjTgrLSGDjkCGz8b
o42TtrXePF1nbxV7j0CcrGIJmwjrl7UzJmVCzBmQibf2PPa3x1oRQ+e2e4Axd5La
Q4j8u1nxctOjRwTKsDOeFGcky9GPUTSK/DoKBeH5C1qklxIPJl5djzNmw3lxqEeA
UTyM/YXofVSNajyJuN7XTfkVzlXJNQlYfcLjcYZoLogerV1SbmRRP/xl4MUNR2pd
vrJsugb16Y8iheUFCJDjlNL7JByjyvYdoay/nUVsckLtNL0pNaB9YVGQ+jknHzxh
7nz+aCvMANc6JC+dsx6k+0eWhOzmBjmKuWDdKp0+BuAA+69XAT3Qj5ED9o8ePRYT
D01OtAELMfEi6R9qAWIyEP0C4hTu7PXIDX6uYR9f1uxpzRGc8rv/WgVVmEkiVVs0
X9uG4xWr8bv37M0iUN4LAKmOxYQFUUK0ol6lyJqp5yJwkQnkvyLfEsRHnxpmyRRu
oX9gkTagzgF+Ox10D8+fJVk3OGBgWN1vLJphOMaQZbXSfOdtgWuWH6TyI5SMpegB
m5YCHDRxdNb9vu1732BBfDhR6Ny/gaZToh6QLpc6u4SvyBujwej/YU1yKmDuEveV
tGA/8HiAZfTk/mtQS3WCpuv0bIteDkpNedwwPDYHx/FVOCDerPH3XbvJuspo0rZq
kK4Z8ISzTsD6oSjt+osN3wdEGgfqCDEEvkadUWn1v1sFSpitFu/YhODXkTJWfzY/
zi4Y+iwJhA5I6GTEtcouoH+jCFQr9hW+1POewjOTdfSVtO1pO7cLbA6Vpoefj7w4
9DgEgO8EZ4SoaUOdANRs0Cz6qMxW64Q0SCg1u2RhteOFY/Df5E71LFyt9js6TaD/
V8mXalcePc7h1w5k8/3DItoOoptQPZ5tfw+rhPeycFkOrrs4YkPW+4I646Da5GjZ
PBnf9G+Pmat7Fj7hokE4fO8qQhtMPHtvcpxGgemz9s8q/4admmrwLOFmwRgg51K8
wm8/vNM3SkDHveY71pctaMPD7u/ZU63i4soHQr21rs0844qZ9Q89AdEsyQe35dl8
mOwfKamDAjuK2Gl2BnMnfomqVz4cty6YtiWgPKRSQri+h8M5AwbMw12w5d+BOSg2
mWtHEt69CscsUbaZOOE+Suj5sP2naKL4vS8Utk3Aj9YZF+T12neyftFgGWw5oUgv
28E9GymmZ50QHDb2/BSrr3mcVwxRiYZbCQVbwwOgTNyu7kkuy5M3th2ut9wi3ID1
NfAx1M6FhcEaxjix+uT6/7RweKu9jakBkMX1uRDvzCjlODqD0nhJZyYqKheevlLr
6Xlo2jwi+5fz5VMKBohosvGjosBPd8hVwsEA3NRCxilAq+ew+eB3a0kZDFEhHQeZ
Kqa86hamESBgPoIZj+SfHnftsNCfN0wFtkRXTbHz0c6cEGNt7x3k7fv2KrEtWIT7
uq0FZ/ymMPLT/gxErAD/WCEoBeegPx16pgF7RSgQ7NObbecrOAGt6dk5XhP4jbZn
Fww28QwsRghfEBOAGt/yj376dS07sKgFlggorHrJKC60QcEFz1POwL2oXcct/PO8
tWVOvuScLD4qy+QfcQqAplNldNWLCBvOGbxIyRuPOrjmKzbYk6mwUO2VdS+/1bFX
adhHRJbt6AV+3lDNl16c0J/qM7Q4lvK2abEL2FY+BD8RTXUZ3E2Ub2epBHzfbhEJ
ON5xs9YDKGPCCrw15bxSxwnhTg12d/BJAiYrvDKRqVv1phtsNrjz/k6nnZR08GGe
zDrXVYQBa+oi4n9yYbjZ9KzlNOZuwDYakvDvnOugV2Zz4CtmG+I40sm6P+qbyJIV
e7m/fbgHHQUCTlT1T0HSv1NAlmm8bWcMNSmj8nHI5CgBA+zpBtGYVhqIzenDTvYq
qp3Cr1HnIuAICnAW7ABAfSROWiP1CNnnmJ2k6IXbKRnUY0sxOyBakKG/60micjBn
zCDwuqFj0oifh2ZpU/ucqxpxPLW6j7MipM2GVAFxGP41GAd1XQsV9fwcsXS1unJS
dZVS1QvUXCayfKbhMFjzf0UDMfx4E5qrozrPQW24GfkOSXhK+25gRW+FfQVXvIBb
bh4KZqwOGYT51xXwtsys7e1bayAwW7eZrHVVQchBZi4YJs2UjUGqqwWPEGm/P4xB
qkZzP+mtb2aB9e8XZjKWrw5kS5he+u2q+2uazu4r34YJwbHaUse+O1nsU6EP/8OV
IDuZYDhGMVtac7NxEpToCO29ZbbRDTVPgci0yNLkGQs6s9AcxE01d6SO4L3m/K9D
nF6qQ0PwUcN06oc1yMlvPFZzbHnji/eEgkRezRJeTpHT5W3uk7Q9SQx9Z1DgU5yl
NM/I8e8iZSpwG48PbzYo/ts8iZWBj8sfmVM080tKEHKz61U9tIbutIOa4PzywA+i
WYW9/dTeNeGZQn2oe6YO0vUGNRWN6itM2VTMkObIoUHbunZEfBfrrMMI+DxVHgzG
qpEeDKb1SPhPK4SfzX3g/csmD1h5cif4UfkcgvFGvlZUiNeKNsFIu4PEEmWwNU+4
hphRgPtVELgAe1Yb4Q1RgTnQUUAqSWfkvCC6VBPGAKO7EpgFeBaxkX0/YftNpmi+
0zqBFZBaijjTvyHA5GB1ciTgQGU4PxqaW/PhCMBK1dTdTG7br9pHfyeBVlvnhBr7
sRZK6klnbpFo4F+GJj6nby8nmApK7jAxg5tt3OmOqNxKp6jZaQUEyroEAeUHVtPp
AoWpi2Q/uCW90zEWRg/ragNoOX8SmAHVOj8IxnqtTbYvEE/Jv0jnpnmsLqd2bqHN
Sqm/dlytqtGqZCF8FBhKhSIZ99jaUqONsBaqPWzo7ecp4wk3tZmVaZ/Xn/ZTTg9P
OKcdAN+EUj8bTpxVN6O7dtvdnRNxB8eF2wAvk6ZWTfZ4f4Btf6jqFXl8I8kb0nY2
RMwqnOOihrUtx76x7aP32lz27RN2Yy2ttuI6WkEYFePUQMdR1xDqK/jpai/ZAvJV
jkxaTb0LLyg6960dQ544ke6FMFSJudO1Pk9w9pBFxA55ZeqwBiYUhBNhMTIgEiSM
UIPJrCrBYqzvoFPqRwUP8sP5WTK0JhiTHxdnfq3F1YiAS2gUj8Hh8X0lEsjxBHa9
la2C1RtJAlWDUPKFZoD0ZCCUTnEwhwxhPY5UzdSl23MxtIVJE6jD0Rtgq08yTWel
ihHXyA1dAsDSXKooDdLZhjvbiE++e3XbNqPb2+UbPu4pscWwZqiB0in/vbuWoIJ9
YGdneys5ePRf6Na3hhgF+tRAE7SVGBdMyipfm2F77AOolqZ7FNEbybiHE3NwzTFD
BpEN7mp4NjwhPxM3GiiBBYl9GOVwere/0obuY6lU90asUHi6uEe4MQjZXKpozDaY
0wI2Sb8zuDL1pE5c1PWvaC4M6BXBFTyS8tg08JfHY6T2mpntquwiqLqFn1s4tG9x
k3VSKoJv/zl1d4kELIjjfg/0KOwwgxtrGCG8H7s6z7HP4qSjTZIAt3fw35Hu1cT+
HCJvceJtC55hg9LlYCLWms9aBeLQWjM8K9tPv8Xp0dcZOtdHmRGQUpMRdTIdbma3
49KZl/7zoS7UPSFjBjgawWicEhJb747RU/nwKTGUwRArtzXALplAVtzakATwUSGg
+2B9Vpy0PUF+NCt9himtpceBXyWey6hdd92is3Wh5A+bZnPlffiERq2FEefDkK6e
IPCuCb8XDoqI+6WNI+iJ8z2DyYWKY0W2ugQtc4N1bJkVLeQWB6vstWwc8TVn2qib
WTaSmU8Dlq48KVMXKxK9EEDDjUnRFox3G7DoDWt7j18Cez+vkz4nFwQv/bTNA5PY
xSFtcN0rzk3vn7T/9Yok/VBjk5XQxTdY9ljU/mNeR+wEloxDVblNjJ1lfGT7GJSQ
vv6fExp29jB5li3gRwoHoq1V//69nxQttdGeSeKTZz05ufqNlU8Y3eSyYbU3oAqw
4vA5e7N+PpzM1istaC7l0eYNK87HQ8g40FDOFNCV3/C8aqAHhq6ZF4HfS3Kb6kN+
VlICJ3OYWm6Jvufj0WQUGFCA4gMSyacnJa2cIjKEZaZmVxJHU5JmM8UrF9RiSbkM
dvYO5iXWfKjYXF3LXStEZOHFMtRQOnCNnx5PjKJ7rkdxRUHnsBbvleJqUNupMtza
VjBclOWgOX5vcXqyj61TSUpzW9HZpdCM55ouR0C2UlklpSEDqNenpRYhPVoVLYC5
weLVnQ+f1m49oBoR+H7h3jYfcsR9QKLu3/ZuKtinpaRDaahBOkeTSvuNbh92M9IK
RVWq2/B/rG+MySbZlv+gQ1iOiQywipmA+rbPy3fx/HEn7GIg477VZojfYaRJEGU5
53DRtMUYYX5lhSA3JtgkxsLHFgQZ0p4owWfXLfWm+0mM+4DZ8Hs2cPGS8E9ocxRC
jp2PrNNiSmZr2B0WzJBY+t029dLXTzZuTjc+VhIbHoS6hpDz1k49qHgVaIv/RPqg
Kzj0Mof1zfXi9Wo3S+x0ULUwxAxT/mbz5GhwvQjeW/5eAl/UY9wOszPf9mRLBhWm
hwLamzi8cjgNmAgRRMoF+t8xHAEWVIogKJX/hPtb1G9qCm+YXrunG+Ipg81FSnuv
A4qXEsPddmR0AUg9GO0Mr2gD9hFlMLxt/b4ui27j+2NX2xBSLs5Q/NwqVXol8gQ4
pLByNFi40uJkPpUvxCavdYc0Jpv2RHoKFPsAr1ZBShBi8nHRSp16dAAD+1bwcYs4
Z/FSdOVbAQMv2k8VRwh5xm/QbzGbKk9rLly4QCB/8S0PlXChNAb4mED35bL41o/+
2HrDhjzVGEKK95hgOk6ux/4WfW9IYuM2BWQLvdPagVrfCkehGEmo8GxMd2NhHSiu
DLIVs5L5HzLtVXpqEWOtj9b0Xa0oxBA1XlZLXS5U8ntHMZmm3Qxo1QcMN73zikE+
yNPoo+s3o+aNG6m0Jdj0NKvm460IossnU8E9Y5fv0zi1nCcSpnWCWXuMiYwHZN2H
dBXJJ5OSBclIs+76QyupduXE97QRZPf3o9e7E6ZCnL+0QfAzLWMWZdmTwMJm0rHL
/C5FkdCaaVEPR7Jge44MzIEqpsGnrupc2P/9HdI0mo8UEUz9CR3uRrFyHHvoMYEC
0p2vRtX89Azn84SmJprITTb0lSh8Jg5J05f0NShWfbYwwSRRe6iOUhS4KhsINOo1
Pm3u0gdeq8BK/quh+sHkBW7C1RISr0fOkDxxhLcQfXQHLYFpyy9fU1M5abcFPkVz
OrOPN7NO1eSxuml0gjXS8n8I7nNHXeyuHCURGcfmbRMbl3+h6h1Vx53yLTw8I5+B
DsA/J+SLIAkKpPFvPc9SC0C1V3qn8TV0FkYNX6sOpHiK3uBqq0hkLkOG22TUTZVf
K0uMJu8DNJFdjxs9OU3Br3Ghcu1qMLzafD9rxOPDSc4xKXnOJyGf4MuI4mKU9UBa
7cIGT3/778eAOhq7D4uUQD0PfrX25Tox3WVRrn2tYG3F/aqRkXHSQHvaaNz1GHbP
K5jdoBa46F8Oe0VxJhPZ9p3WuwaLUFuDlPCmFLcXQgD4i9SXya7RvTReXulxmNSP
CcaLenQhUlg7H7JyCmKKgNly04zFB4OSJsKiuC8sInzspvdkWtyLBRIM/L6YlxeH
D/nQL1XchV3tunxrpQaO2BPH8M4lmCIQP4g+fndJdRG09ZtV/noCEVciF9SdVWSr
YWJqzizMs2pn+U5u9g31l5neHkiCMA9lOm3qXd8CNYGsNcvtJZHFOgxOygOin9q6
UJw3PW3qVpO3tLKnd9ico627xa5bTKg1GZBZxMGqRBWOELDuzqx8AqaGz5bcctiM
GMx/kkzwLzRIX5UXPjRRh1w7yoEqsB0Ry0CTF8JlJPd5CU7tRgLD4ExZEzWHaIg/
qxlBxu8bFM+zPj2MPEQahefluIvvaxAXjidj9IiwO9lg+WiLw7aYSHdld2tQsBwP
vSU15UvwYRWGUeSFX86SjJF+Xp9ghMsuDu7ikTO3+He/2raKwK/djPUrNXBh1v7u
/TwkJVjH9gkUWaTQ1yyO5lAVP1qgJcrLEUI1E6/3wXiMjN4Dtnh2xR16jy5wbKVS
DnJ6WGBSE0R7EO2RLsv1Y4Lrt3qyyelnC79mfCSbmYUmaRhnGP9aDVOHereFJDUg
Ku9HCHg9cw2Om0RhpWdSHTQL2XI6SJEkXOmDFifOtZl2TCZY8Z7oqDbxGCnsoaUK
Rq7Y1cuxT3Gi35H+ghwrI1hveD5Qs9klL2Qa8LTiCzTVlbbhYKmEwiJmidwj/3/O
9KHPqHIihzFb1YJGB2pCAS/tG5eN/VmZvQ6LhFkx34O5gKtiqvQbfasRM1DpQ9uP
QU0KfuFcOJj199MCBYbRUPfmITMgZNKJ9/dBGx4b+xFFTd23JfPRqjgalqf4MLdc
/xo7O3IF8YUERR9FKJXEuYmbrOHbBuGYBRq7bqqTCRd00ofDA+ieNtBSgRr/r0N8
G4wYuD44FfFYmA6MpmaF5gRakEChNxSQmtHl6ZhAyBxdge3lOAfs91BW7YKPy9tv
BzfYfBZCXzp1QFeuga6/OQFQOrKgBvaU0mPlM2DjorvcadlgXVx1hvtQiwFgNK47
9+LUoI0jze0bnAJHAnjD0EPwln1bomXnDEzbLAfdVzutF8yPYda1bnXnPwFobZ8j
Uhy+olxqpqM333QVLXDAblBwIjUHU7saYtrMJv9cPdLkfQ9M2IpsQ6pwTzvcxk1J
b1+tsU3OTKma/9/ldWXzg4sHinJvTBmCSHRYmyVKm8DjuPWza4hGJDlmWu2KSNg4
fsZaB9RtyfHxpzposwqQIc2t9Cht1HPpgVjvbce2sxQuyJMMHLL7euZaHsW3fvc5
lJRiiOQuA1b75e3ciedNqEzffMPar7Xi5xWZdDZ8xYq2e/j9VztRf9fW4bEeileI
6IecalDNFrjjH8HbaVvjb1E03wKq4DQEZwGPm8Qlu04KgMMXu5z8tOrGY7FtKQk/
GkWGWK5I8qk1CKQ2tVtZeZVfrLLKhIUG9xkBFZbuRwC7e+drT8yjoYR1K/vVi5Yg
Xwp9FTkiFS8yrQFJM2qqjib/osQRmwFgHuYPjIF+Dao/hcJRo8e1yxU5B9jfwnrI
SWAXVMNj0gR1Ps3byNEteQo0ZFhZD588NSRqNJBs8BA5QCXLJJ/fQBSQ0NhcGTEp
o1270CBMjZvblCuEDTzdLqBIZStEvp4vSfs8HbpZKwIGEvuquEYnK6QFmy48A46f
nk6PBL5MC30vgxobzvSmqU2/klhbmXxPr7Iri7+NWscMBiDAfpm/YwlCJyZKK6zV
X/oVvVNcWuRPfdrqfrg4vg2nE6/oUojV4fl7UQKBeykVjXfQKPyUwPUaQm1DpVbf
JNyRJE7Z1vsbQT9VbLKZqOQ2OO0wqqPf7IK/TGtPtwA/3OXSTGadjtHqh0H2ARe6
REh0E3LQ2h2LHjX2c6YsnhfJCRxBXSRLoa6SQv+nI/n33bDr7vgpp9bAc30cOTD/
COj9umNFbMrsQTl6fHKzeQGS+3Enn+yNS44tPmf1GkOLKw+O2QYwDdUVbeE0mRRy
iiDMk5T1cYEJpzYAwAGFmy06wc0FDdN8neFxDywKEm54xiCWMSlPYQnvslOq4uz5
EvpDFU9rh6yctqXZvs3ezhu06AHpzxBiJSLNRiau6qKSsnkeDuLIC3oSUiWJsiSB
GUWNTtkEMwJ9WN1XabWcaMhgH8LASm5HU5fAQWQ7qXNFKs8yjeqq117ZU3TtIaXg
2Dfb0Gbdlw2r60lgXtHGJ5vuDNKETOVO3gV8FQAh+Rsu5CFnjxYdfWG/J+DOoULv
35nEHpuhM8SXS6BTUlQr1otpoELvfjDsEgzzrqwGpWzn1LL7A53N7pyrD1ASBCWd
k/T1dt66yuwPcwDRuBN7SC+J9J8jRhb9gjS4D8q418pwLlpiKujQgRQ6OiKpdtNt
RBARDPu7LDFhgC5TsmcnA0fy7R7+0pFallcC0jBixlvU4XaRLXQ9N2x6wl4rK/vb
zuIY6lH2ZQ2l6Ys6ZllN3zv4zjpV6m9QsdgcHFjzJe7oM8f/3HjaWUBEpkzDJlXD
UZhojVZHUjMITLKCsUiwNlIVim7rgW+GjJi4esBQmwqvaTJHspI+QA+XvqG8HvBQ
qKtY6PdQxS8ipu1dmhcEWVXhV1FOzOuQEvKIOVKYcIzhxLwEDGgBXl5wUc2ejvqV
9ZOXL+hgqtnxVRKQeFHTQrtEY2fG6w3o6fCboCZcORaJdVW9vkI76mX3A+OfZxem
nP7p8BsqQkD79lLLZwgwTkaNd8cB2+IlwTjdDiH8PKjJkKYAkY+pkzAE5lBMGsYV
xZenvxKBerXo9gwgblWCYvb9wTlv5LjxoBmanerTpwJmBGjIpyjTqOrz2OX23lmM
YfDzNP78pYLF3z+O5qqF9NifXTWE7AKYzSycp2t5GWhuqae0QtMRCEkDLr6KRP+O
hhYLRw2CEPA1DKTICauvw9WO4gwfn5E8lqBCZw5OQp+KIMkCDuT/tDHsRZ14vd4W
7XeB1T0UO1imGqGVfKiaJE+iLKxezJqtmWurX2HdiHAJPpaBt9I1A43zzBkZsy+J
btzO/e38Zhc9uwfYtuyZAP0r1wjXEOgNmHI2eXl4WcVRVVpwb22I8n27a+CHE8Hn
FvjT09LbQ96ZFw3KUjPTFy+p4T7iL+TGV3oa0Lzrem0hycxxN7K+HQUsDC2hk2lD
8PwFWBV0qvKzCLzR9iVVbmuM3qKsS59MKxcv42yzC1HVblYgm1d3nVo8COudpDAg
J/5UYRkb45uck1m9LOX7aP9ylxc9KBww21+TbLGqj6Dgr1LSPOrBYcxTQbQ+2U3j
D1J222ADQcFrIjM+t/Y4ySe8MfXEmQchVSC4sJhLl6jvYLCMkNAIccmCGCV8PR/p
qKLQIk24wKGAqkC+y54lpVj/NLVqV/CcxAzQU9Of+2w7C11ppGO9D73l7ht5vhQU
eV6sWxkGx7oBulH/p00UkJx6pZu5P6G6rSZn1udwpeTzhA2j8SRr0rk09LTJZEPi
uCprNU8HHM9XOCyeC0kR2WXlHzTkiYpL9g7HVB9OZ9nyM9zkd7EALplDqRWbgl04
DFxPPJnDYiZjoEZGHh81vysEw9Ea2gI8mNoi94t+nn+p1OdHergNly2hf5aKfTDz
vI5sf5d6IQbKhUwlJIumVs0Vz7dncm2BS4bEky0Xbx4icwveOC2igFxJ6ocIZlsj
MYqf3IKoZ6mj+c97P2alJmZsAAUWR38EDvTYB7PDUwV/FjRVpvB54VQVUmzxiLCh
qDrgZ4+jXSwD1cmodS02i9tGYpfu3v5D0cAgW3qfykh7a0fQWM7Ku7GCpW8Xr4MX
guObFeDQJJ4t+5Eht2oYiFvCdDqIMzWAzRO8XTYffgzqXTQajNwE0xuYJVSUnwvl
BUPiMkrUs2z1aQw4F4szbdo5zhkaLNbMsWIvCKcNdS3oJ1OJxXkP7eIDJ2dB9GAx
pC5IZFPp9mUZ77enfXu3i14Ouod+3J2MbFm0sztJ2BV1fyvic/nsTzQ+y+jZjmkq
Shjb6SbaVW9j/HzUxhK9M7NSZgfQJSz21GVDSCXc3ZPZSk/s4B/BrJfEQL4la88q
oOCgoIWtlV3muXfW5Epium1uORmD01AkMpEPpwH1SQQ/7U8lH4gTSMgE6dKJDoN5
ATYwN1xjlHOvRU7bUwmFmGhRbk0B/OvAMwzolXf+FFevk6mGGDPwGhfO6x4tBU8y
I6HK3hBwVvWcjVxCEPazc5mbj9rTcs5Mb6IkD80dt4MRIgIa27dkFPXSBExuy6D4
yD7TmTTIoyKMcvqi6m0Kt57aWpfTlN4KxTL7+jySZY3gmr1XkqUiNaVksK8gbL4Q
Qt9DNqCFzm+Dlim5/njBEH5kIxjQg1MBARgnSEl6LKTrrO1ubSNCwoQ5IOiSTmGx
ONSa9PmKFRppRH9/HZywiikItv+LHtJn9oOcTiMzqzNEro1glQZ3VIiJNy6nhk1S
J1walzVy8ACfCFyQA3xMZvyZNP7zhqe1MPRk+4YcVJzepTFwDOJpRlBxSudCMtSa
FbkaUA4OukWkcv6wx23mHHvGxUZW+sacBkywSUdzk9dmhFQ6dhtx7sqpPI1drt8s
V4PGivMgVuW8DCo8qN0XneDb+IehXVL8OdKMaZ0ViJsjRadfbjPjkNgJWSFWK/pJ
9JIw54q9+Se4nDHzj6+WGJyn0FMSBJfLNd7f+2YDVP9z585PdUBLdbVrdpteA6TH
KolyBfE9MWxBEHfc/fnN3R4QT+iHA7N9IEFpJ1vGJW9vsUq8AQ0eB39l5EAE+2wo
L0n0sTqAJe926SgZpXLzfAaogkr9TLal20SpHyB0+Wer6xGiS5i2M+ox6bS8Zi6H
uX3+fhdVZi8ghek1CwI3jjfidXnVv/MGZIpebNs83CleooWiZ2nQSf5LpHwZG8Ri
JMsiHJiFEJSc5VUxP9H5l0egodGpm7OlQNPzngT5abs8nlUiIubiMwOPLzyyFowk
dWHAEldbc3P1sbrBvyJbrd901RZcFimL8ygQAyrBd7OtkPYq8gnFVlKFRympa3be
GsVV2V9Iyaq9DdhPrJb3pSsA8iOi79ZOehjF4FJDPa1u5oSZlwkskv7JwSYPlVAJ
WzQmyjfveFv58dnMTUh5ekxzOK9wpde8Jfso9YXcCEg80mHsshenPrbqbBlGjZLT
SUcU2EAQHsRxU4rqAg/GoJP15L0m7bY4BoNsqM4+wcC2cis8aPKvebkYoYlDrBkH
P3uSa2vUehgHlv6icJ8UGLOztD7OkDpO5v2GZYuribdofX4AvfEa0PvnKry54VJO
5C+jfz1KmiDMPZoa4lWZaTBw9aCQaakjqlRSakhTuCOCU19U2s75PKM/IrMdeMHN
DFtOEi/E0HjDNZKgPgv24ut4bzHLv0BmDQdQye/YymQuVwU2iviITvboGk4L5qdD
rpGgMf7fVB+Gi+g7DBPZikx5Nc1uwD4CkWALp1ZHsb0A0pSeqx60/H3RVk4Y5fSM
QMSHiz9jBYEUjYFsbelDVzNN17yYsyuxUvEjfcak+MRWjHNx+yVT7svch8viFUD4
QZpwciDtVR2ukZmiFQmBt3vXvrnbZr3m8ifz6FurVtovom6teRvUj/TWfEpDS0Sk
5vXfFF+j9XelcxKpWpqopB/taYbCugTNRy1bUnHQp7VsIRvGyfsjzuw0gR2B06b6
ooQeBVgKHN//lY9DDJPHe5kE5bR4VVve4LojRHrPMkBOFBcQAFibC9QoZGVD4ESv
WKSjN5LRXi8UuArKSgTHTgX6SjCrmVC/QA++jl3kgesbZHh/uD2N9nIywrmPgunC
1fDsIrby+lTzhrLH9GOGr7TI5zpxr1ipBcwqSi3/b42YyQWH2ODQGQ5auKFQgJBT
P3o/H59mkM0LLyrwV2sHfQlDG5+J2fynBB3/hw96QJYDGBNMQnfop9qIH3yHQ0/p
TPmLUXHpfIDlD33kmSqX38B9XYJgPXBmlpvvEJk4aMEUfeWto6KXMNzfED6lHdkn
2X5GuXGRFsZ8ue7L3cWSO7+vqDeF04UH2dm4jiXyTbfnIvGEsIo2dJRG0MINe5iS
uGkeyNIl9Nj3YNR3OZc9UsQ4kMlg95bUC658GCrZYw6cAhNZxnAGfKyNB7s1qX/r
Zn9I/v/g6dEmMZ+B0ONYQlklkfeXGFEkVDV+fKioKvzWca6Fm/F20xVlcMQuIjDe
JuoQWbVw3QyVSAiDJz8owSDrUoVUWkdB5aYPNWmtXVsAYGohbaJsnbrdrWj8w/LE
ZDrXrFDLD+yhMIT5BQgxhejb/EgQT9L84ic3vJ4naE0Q7FBhlSQ+Km6+jNr7Q3i+
+Cy7ZsWbhkRMLmLH5/QysJebRsU1+145TqQ80IKr6Ddnut9SR9K9dSxg7vtPGYdO
RALjGBaK2NX8f3y1OeZVEtgkiKQdBcHO6M+PNU85iMmre4PIziAl9wUO/HZxg5a6
2kJr6++7+UFQZ58R0KZkQr2I/845z6HH4Jfizj/5+h0hhSgFgg19KSLvR9rTUyXJ
eGEZi4TzviyOuHNCf78aYHHkZq2myEQJsa/MfLsh5nsB8J1QypDVG1eLAJYlmZvQ
DMnMGzFYpuIHzCziK+REVDXHAi14RoOB2FmocbBLGbbrssyNKGRcppSCR5Kzy2O7
qTPH/07T45gA6y6wy8qF3h2A/gT0NZuvSaF1K0xItQFGUvgz/tkXATtPA6alNL3F
JTRCo/SZXheixqg0Ha+2TqitYYtvwWgQLT9KQHYI5spEapQ4eFxq49VoFbf/wNsT
ZHGpJz7qSv+O5lsiNhKItM71C31wwYJ6oD5i3byLN2lJfGscKpn1lx3AFG6zV2bi
H1LH21k74LXRrZQ9cKtrd+tWKXUNV/NhuK5eV4qOLcFt4iHM+NxgRcnS4SRQJAlY
AevQp9+ws5HYeR5Wbd7Pmbq4q0WrN3s2DoXoTqnB3oUoH09OQKu+HmwODajOAgb+
apzsJFHL0NQfId+VqrG2AJ5UHACHNPk1LoUC6pkAIxh2EDn7o7VsA9Sq4BqtxbVG
O3z98EeFMUPJZcztnEAseWGJRcdkygf1/tqHxwsfGut3o3I3XYdKhHsg3LdHDyH0
+RthfXMmMmJMdP44VnqKsIR/rN61PZoUi9aG1ALiOV4GoN8lB3+XnVrNUqb6Sd9N
lL9hiNTuoxWBBM8Z5/t8BF2sPujENVO8bAoWEs31ZmloDF6FuPWYPLycm/epgfmc
q975yXyF+F6JSSRa4e0pEajxIPkLMiVDwVwMaBEzXK30Aw+9EXs9gWGy+lMV8tLZ
sdSxT9Zs4bsGJWXIBSzTuTzJPkGnqznlFvJKl8FbEFgDbOT70ECsgDiSazI5hBLJ
EP7Fp6ZI/8kaXfcRC5naCUKb1Efs1hCKM3I0XA0C2HukKKDEkNC5RUIsLQwe1yfJ
tW0a0lmQAnCSBaDBEdqJD8nNpbgg7U3iwWBebQLyqEaMygHBRw13hH3EGJHf6ROJ
g7UfGex07QF79iRIAv6Pj7DEPseud9kW6jySJn4McCBWdrJJ2eSMShzip6ifx1Bi
AjhiDi4wUrEnAl8NebFV2MFvtM8irTYHivpYU8zrXIywemXxyLmJSwzTF0NGmHan
fVTQuh1VkD20IV5JmZejjvkVbxLqRpzBumnGL4PwG0rIk8oWhP0tePEIWTnrHY4p
KgAEsKhL+/VMR12/3KjRPcKe+6Llbugu7ADedToxMQFjh4++2jlOj8ehseQd4LG7
YWnJW9J9S1GGfDBLldkBGbh4w5k2XqABw5sH7SqUOB1A6dGg5eOGS91xiyPE8lfS
5b4I7je1ujfuWzE5muVu9pp3p24eh1UEdG3vODwJ5aZ4wKj9EqwwIl3+i0SYeMnC
v2LRvksv7bPUFBrCvAlZFzUkwBROWB+YqRkci5QoVZ67Bezs34EmDAUtzM0ASpkv
N4MCHP0XH7C9EBhrJaU8qSi/7KWAMBgkXD2+xQ2G64z4Nk7yuF5e863rlly6RE5+
b50/0a5wG/ISmJK+5FXFTYaVjIQuUxjXK+DRsPWOw9NFojG/mRys4sgAWR51kzYT
04azsoknnOKHOWYxeF/zEmKaEvN1rPPtY9DMrVMian0Y1ui7eqeU4WWWWjjT1ZKr
GtWIeDi21E8wzGe8PDSoqlN9+lhCY3GWUnnIvkO24KLij6upRYPVp6l2k7g/Mlon
hXosagCMs4UaczOZZcNlo/jRZpozRFEfRCL0rC1tatsq3cZTmACUBxleyJKUj8HX
MNtKVmc2WUpfuH6/T9VOm53QLu3WAjXO3aI99HWk277gS06yRfk/HmFZyOciwoDe
uO+8pZThULzyUWZM3ibseCT2OjgMXBzaNWDurrVhNHKDBkh67Noyp1lDqTCaefCA
VbWovHg2U+lrfnyufgNuGGF5ZuARMxinuoqY2ndExQOFlCg35S3xeUAjpCJyU2I8
D3LigL6bZdp9b+QLUGaBmDh88dIdpz0RHVqK6hItzmMOSAMsv7cvlaXeqsSoPZDo
Ysd2xqwnr7af9sBpotgBle+etKzrdhXP7gXhgGzi/3BtLKhU/Tkda/c/IU6Qm3bv
/uOIzUeOFy1EAvTpsOyQSp+t+mkabhozoEpxjofj3a5DAVctCXY6S7peQsv2BAwy
MsrIU2T1gTWut+V5zJjRRPq4vkTv81pio59qibpo3ieV4Mk0AsSAdIPtOSF2YNJM
J8CManHPAclYOe+ShGDsUMl+RuFtG0SSPd0ZaJeGy3dkKRw9RjVPHg/OXYTtZKI3
/sFH30GFdjpxq+I4bYVaRxdeuF12op/CCfVfVS4E/prlFVhjXWFhHvLW2Hvu76kc
VIOXe1KGAFylwux6XTMHktM+y7RrTAQPRetoCGIyBygsRkH7riMsQ2UFUvCMA0uK
jcxFwGvkXpO1r5KJmtdSMSnHMbLwGeWerZW/QzZJabxPn4MUeLuVxJypm2oZWS75
2fojF+pka57RMUOegKh31qnr1s2Lb+OgEW6ebubJZe6AgmYBCdCe4zcdPxdIukut
6tiZ6vl6q0WL+JigClzsZ4GPoP9zLfvgT3k+qS1qb2ZrT8oAaWmLFbA9E/nn03Hz
khbth77v+jXWceww+GbtVE9fUh8TthhDEU6yY8QFV1W4+2A/JvcKNcvc2T0zrAj6
/KeAxF+4Sjtot3TqHObeovucH48gXyzbYpkWPrty6VIYIEMwe+oKJ2cTa0n3rWXv
vUeV25Fiv9Dez2Ob+ID9OFMWMSJ3paQjYpwj8ZBSVclRO5mu+BefVR/m9Kd0P5kv
lpBrq3qJovvK0ZE9tdq6SHdSrovp7F1bAbDIoEci/o8m4zPo6lWgOW02bbplHVez
wujTqRbG43Tjw4lydAgu+cK/7m7a+dRbQu5djVC3pco+eQwlA7h/m8NW5ykx95tS
FDCPSCwJr/C+eMK/BNvdxl96yBzvQERgxv7F0STpncqQFV/u8z/+oPkioY6fPHBO
saoe7n1t4zoMia7cMBvrmh3NIYf/Aoy4X+YhOdzdj091sk2OtOWujQW2xqrU9AJ+
a62wkMWANykL3wxHgJnPvr3niu2F26N54bK/RRPi7ECLa5cnuAN+2II4L1S5RVJ5
Rbmx1fXXrjl5oR1fwFt481xIDTJRns658O36O7RT4jVAPCj40kNpO9IFkxP5pBDE
mfkipNOrW2w0fDR1Hl6jgYoaDcgi0TMdfacVsFp6DoA/BOZC+mKTPfHy9ZvpHxM7
nA6IXDZuWM9wooZQ4+rmW8ZMHLW+FCYWU7hm2NAevjHRDZwo03kvoJExXFi6kU1G
V/fk6WnOXy4mMHjrJF085ielBPaWq1mOfmT0zBmtSIBH3Pa1qaiGb+RrSje8J83G
xkikYkVPqyNTJLQwm4/Hw7r5t2SIQOngg2j3fqfzmlNmsdsD4U1gi7wJ2Et3Ag4U
d2uDv2Ok6wDVgw32zgQu9jV7oDYt8WjiU45W2IJVq3zquQvPEDQGMUjlurQo6f0J
NGtexeIq4EFwviSjeudQO6i6f+mWsUPWlj09JHOZMleU3tlgFLafq+yNriWxebeW
QicNKkVVeoAqc+CGDbgGwMgZJKxN91grGQDgr5w7d1BvSv6tw7JRjIhMUpGXbRw0
lAEuWSwQkfOKTgZip/E3lll+Kgn80hbmZ9SYsCuCyftC/IBMetY8seSR4tirnr99
juQGO0SlfCBYgFwmWU3VgLbZb4SDoGQG7A+fAR9uXNA28ISAFego8FzDS0zb20MC
8GaYSYjbTLC4T2Z+5d5zYp1ioEisJSun43lwjhaSGj+MhEcF88Um6mmswJAHue88
54ng87vJDHRTPypmWfIORNY1JGxyB4vGGTcT4TuFvKx/Z3lDkL6DiyJOaAKzN8k1
/zy+PoJyHjepqvbw56TtRV85T7/zFeH+v6zQwEcpFu+qR+UPJTICjsuMY4gojbsi
dz3B8dBN/WpGr8MXOEPDG9sw6F19Or+4HOUWgTTpAzYIGvxjTbd6XnBybXruedDb
Q0ZciBir/zGxBUYsSt4wSq82x9O+Uj9rGgSv79gsDYjuwE/maf14PwvoZUB2vRA1
l7J6GpMVzgjN6mRAjFP5XoyKYvG2yD4YBxJ2h79iLkl5p1FdVfxujU0NOTnVu5iv
WwKIC89d0agBrWyd+YGgRzZF/XyTqiXuzPta+z3NTsgrrdrENnBxKyZd7ujO0im7
PprZk3NZYTmA48n804TcuucV4igz1TSONtPq/lbH19ZGHs++z0vXMPHYyvjkX++G
oXunaIQMfdYp6xdPaLi7S6e5dnRdMbdbbe23FVqcORvJ8YS6C4qgEOfcXgXCJ5JP
NfXW1o6xhIFXiO6RAs0LJBFkRNSXvMhjIsW23dXZ4gsBPiTFw8yXU+K0DEIewcMe
dlPjMFz/+UEmgrESEZOVH1B3mDzBs40l5lKUScLQ2/M4LmlsGTt+Dfo1lJ0b1jGD
p3BklDRxhxuRFdoVpCasHpLDI5ZJZZQXk9sRCpRrrlyehguPJ7w4+vRj5NbYAfUs
b5WpzgVvZWJvvkLtWmodeWcb2qMkeS326eemf9thPlZ8bNnCdqWuYaMjo3zOmwiz
IfHxCYga1tPTUk7HP+8fODck0gN+dRFSq2vEj4BuIsaJltEwskuLxGu1AEeX0nXA
iJTD8pSpl+LUtRxyrdPaDnOMsiWqReDh/MmJUlhMokwthBDYN+/XP5amiHSVlcin
1V6z/WkHTJVl5J0CNX5L2hkSILs7qzZcbgz39+f5zgErjmDetrUhvQs7ugSoZ0HD
honHgSAcdXlDYWBAwSi4KJiUyfjkhGpukVVeR+YEjb64890HnKYJtoU9xXtMlmI/
Dz4S1n3p3na7YU7paDW1tNDbGlrKvKQdRUjKzy/eY2a2eINDHKUroh/pBQbRkKri
k9z06dgun134PGpYdG5C8pp0OVzPhb4XwCs8WASVxL55lzhN9MssrnLDvvKKBD3L
mNllVr6l8a/H3+bm1J3MYe8ixqd/Kzu60kFPC3gebQ73QTGmG2+4nvlH7QrfBETb
UI0Rjr1SGnJ4GOMOF9zYYmdPjQ66CTgR6mFFwYy9GYfvfj3EvGuF6UjVav9Au4or
AFvud4ZgoweGVRkox2k/DtQ0AUScSHcpGD/zFvCL8QTlYbH03uFFiFwMbQgIs2dh
N8PaHNizn73ISmAB6VFYMqycwnxH/MLN27iFVSjvQzxR3rX2ye2RNNruBWaZvgoz
MDL0Qpd4/AbnsEgEIRJLWcL6N/TBM5jJIYTFMbU9dBMxAJxBM3DfwjVNedYUt6/U
XjlSnwqyB9h1uaBIWauwQHQTddkiOU95ZlxDBHcIsKzTCbx+zpqcwtY/Rl+lku6N
wPxMWqZ61/eY1EMvdKf5MHvbNBRQNq4B3OVzmKMX4l0AhdzhyGWwUYX+SVtoXnO0
Va3Mftvzn96DNhaMkJZ3EGPWplPOLYvPOtvHN/+pKlb1Y27EXmvIEz38JkTUAklB
bOIrApv50YXFZAyB9Ipwg1YJqObFqfm6ZDK4Z2ZR4Z8oI0rO89IyuxXeKHt7tgXA
7xzrY9Q1vElYQmd5eGNfeBoHQhZF4X5it0hfPkJozN+lyR1X7Ih0/gBVzcJukTe6
Li2x8F2JJ8ARy9GAxIxwHxm+q3K4l46dPrOMVODDBwsiNeHmkYHiPy9Q4/JqdXZF
Dls2vl6WpY340F4PqiFMwtCybhAJYwZP8MIUnHZnITgpYjOOLgwGxtjVQA5etfXO
9UaPp3KhSN4SNcrh4NdBkL8xE9PyfmoRMwiqwjsNrPmnmOq5CsibaRCOjpQ00C2x
n2kiPWZkB3SDdwrjSlw0Z91DnajRz93hzlPA8UjOHjFu9PGGb+PMkBkaBraXtwMA
umoIufG2sOPWlHtBZO1pSpeZ5utMVUYhf0mDkBFX5WgSawV7GGBYUn9OXXfXys43
fcgZfN8tC+1ifdzjxgGjgHOPyBYJq+PZYz+/6SOVyqZwzB/SLUiGOeB/rMWjmQ5d
Kt2O+7LiBJ8JvxdlzC33o5zNKsUvPCICGxyB8CNDq3jU9EMFKcyWxIZcuazf6XwQ
uyLc8U78QOpPP9Mohk3+rMezBc6NcIg/JnHgMt/vNJfH4W1gVECtykz02Nwe/cxW
3ucQqISS7zxCbVUCVj2ALwd8+qRtTTG6QnmzSaoDCkXcP/xetjCVd+A3ddNE39md
eaCONqngoiSzwXoU9trrPPGqEqx4m9N0ZCMlY6ZH4L4uiqxwx5tJ7tq+LOQfM920
jnUyBXW72Zz0A49JpA48ynLvnsBT/hBwnFfOG/Uo4mi5FxlfBdUuTInrW5VMkoao
3jLSrRKFppbuWrQZG4+Y5Ed/xUqiaORPxwEhViKRDZ6s+csTE3YhXutqNqE2fKyE
f1cLGU7w8k5hKvIG1mdawrGdCRq4eKOHqqBX5EHatkpiNEja1NWJXE7UX/mFqd0P
grpmG23Y5YrcUzKAbRHChHv8oo8eUMI/nfS7P6Ql6RKPAjx78tZd9g1/RH4WPds/
2/Go/r1MNTA4pm2XeuKMIje8GO97Y0bXVUkps8kd3A2Zzd+P/qfzEYRaCb1KNBZU
Nsdq0QiaK6HqFckd13+VS4/X6sFpJxbJDjqscIZZSgg0hB8XswJMw1HjSzKnyWRa
zi+aox9363VKcBtUNmorb/s1WDgcPV/GrYsiHwlylT70VEMktJnKKmwZg+MQn//8
W4jYPv3I7vgq1w65TCCjOz//EaVfHVKGu3ho3n6Bftj9Gr5OHHPMl14fy/N0AgaH
sUwTCkox9E8/FGGRrShd4v9K/Z76lQrpVK3rgzJyjxP4JKaSw50g4TLrogRjivDZ
EMroipylVYO6WpQbzTDQleWL0UXOhIak0Sm03DZKIuQZgTgl6Rjb45gyJFnfXvxY
zLbz8cTX5fdkIsc/UbpZNQ6qkuDX242V2avPOELZ/BvbTRtzppTCqBxX33+TQBwp
W4rfwvqfaFjB2hoQJ91EL0ke4if/49TLrQUG8EplM7c7XF9nk0M3JCRKIU80181c
0uzF3Zh/pfan1hVek2BCaVBbfnDyxaTVqqsvk3cN1nxkhJeu9pIBoUQ6JflayMYC
OidUw94B15xrXRl5oAwvqqUdYBXJBk+2mC2/Fu2swCNpqWTg30mxt0HXWxyH/goA
mvhwqiSOQteqTL7bNYFkGpsdADlzLuo6VU3x9IyUhsUqeXoxRid1g9aFvq4Msb/C
LhlawzdpbDdWFiOAbiYR6ju3Diop2gJ34RF5l8X5glqw6LtkdXPjbfj2HSfC1qRx
aAMYEpjCZCD2vxywV8sxa5sZYmdEld7HorkS7aX+OR/421ZKPn/98TNB16FSDYW5
HKc9QSm6uwLnuhrnq/f6sGre/JyIfV3WneabpNi7I+2mfmE2ONRbW8QEon9DzP+I
xKCV9ENet25Rb2XDEeLQaz8+NlYKMmsA2krodiIgkOGar1ZaAA1nY+MXjFipBWPq
QPyaHNDtEzx+5fGkWBwstG2dzLgWwBiMIkat4c9s/C90UjaxyEQ2g96a8CCDHmSQ
TEJUD5k6BcTFi3O6ztX+Ytme6wV1ICl3IVb4PELNHeQl3W2YCj7aQMHweG3wrywL
w4pveWuSllUpWzhEjrV1d3n3GVcNJMFrw7I/FFdSvyJp071CLzftNBgcGdkcL9BM
bnuMZLU3t9nEcsaL3uxPklphcFwsiHCoMtZVQnG120Ypd6dxs5a35DC3qEMnfcqe
vQv5hSzkIs8tPuzCVKrXDyP84I+SIGGfObWo/1MeO3YtsPHCgubDe295yVKNaxEa
A224xo2nxo61KDHKf2527L2+TTabRysbB/oVt97HDNm/NnIEDONO+H9PWpsmpiw7
FRXgLXQ2NTlMN7QsxxMb0yCKIJtA3CnbEpP12zgV3qShGEzDCLtCUVA29EoR5mQ2
uVhh9ITuFnw515miU2IxkwB9jPvs+OdYKAjrhoiPvmNkIW5gOTOory4pY3q23hKa
y31a9jtSnZHFpustjGSP7b+6PiO9K29Iq0Fj9WiyD3nxEvLGDnRepaez7F+X9NDg
2QbB5gdrG/OPx2+mIh4hbbrlvXXI67NVXpBgD8pvNmPnbcUyMY2hAf/7U1pEOkt7
0tNG9o/60fJOskNA/1TN0BdvrAYOEDFU9gci2qEn65FYDgJTmmPJufv1bp0Na00R
U2qNXogkCD6+RUJEhj6hVaYb6t33/HRmKD+oB8FFlDjZtNaYYixRgl8CBFCltJ9X
6pFtO8fTvu/TvnEgFtI/vmUGsINjUmsR5eB+LnniTiJhGjKmHz3qX3hUJ83+V6Ok
WqFiC8docxy5Bp9U3gYKU3v7oxnXhSa3wey3FeKsEGSCQW7QdHc6zLgMfCKzUrCD
qxPFQrA4p8R2euXbPTZ75+08pY+FXpRY2IjTLR2OFJpqkiBYy2y0cE1COCYVLt6Q
h2aIaFnQz2Cy9gzmPQsIJk5MPQBgZtCRYxq+HQnuwH+5vaBS8phJjsmSEliCfSMU
fAJ25zdO44OcMeS7OhQeNdcp7KKLXs94Dn1IWk2v1nJukVYHCRpt23by42VMps/q
vPnwU4BoQEGVVJkAmSgYwcxSJY6ezlv+KIZyScM4zOdABsil1PS1JfX9GUOppGw7
aNpSS3zUALGG6zqcoJQKsuqenjYd85BWD/axn/MowJggYkWDrTIfK0cCD8yZbcBP
nPAGYU9/+Vjst7lAwf7nJkN8ki0egQmpfgLtaQC5w8uUcn26/J61v5BI9Wz6JPs3
sflmyJeqO2MzbcQSERRSMo1GJM4ZeSMzRXYx3N2zG3zn2fUz/c7RfzpRGFMBbSmk
aY00GB+1pJBfQBs9CYGDr5/pNQ8PhwK+/6E9xocHfCzsm5g17LLRMpocHLITjswG
BfkQDXF5ROHpDuMT6y/iBhd0oUecuzOtvvxljADLPS+AZ89FyRIaRFIfvrc/332H
NrPygkfHiG75GP/DWesrAOnPtHUHceKcf+YdgP5E1mfaEK+Is/y1qqJb1gy0jC4y
aHdrfXIJnYPKBe855rf+RZsit31VcfmZoP0XHV9t/DuF5bm4j2BMt95XPUkeGWM3
fPM2z+TXRatx3Rvt4B2oS0/bqOfJAFtujhCK0dr/KI2gz8fZbbGxUJfrUS6ltXPI
5T7n2e3kZbnG8g6yirhvYB0CFhQSBzk0oFfBS2kee1B/uFxTDhxaHd0PeSV7oo9c
uX34jFJkIQ5TS8Y5JOGDPz1/22VMqUtLtK2x9i/rTxIPnXtT2KDYCu8WQ5kgv6qz
GQYJo2BvTeqOQygSMQSzlnplaYb7tiUeAecdva2gqowTHgUBvA696z6iv4+zDMCc
yf5vojvwN356kH3ZNL4eczDerU4QJJsU1N1uKzqhUceev3RDj5MBDIDt8kZcjlmG
jmLWU3Ef4nIZF0pSbKZ/r9n9YcNz0XFLGVW48s3Hez30VvwsLPGOF2tNyM62YaCK
3HYnZ7Vv4gEdSGwxdQs8BvSSINGdvHZcSr38bmH95OS/lK9GvLvEzFHSe0Kpyekh
P6pFXdWoj7Lg0P9cx9Vln11pdvuKWkGuEx69ne16DPOGs/0H1FtrK7p8ysM1hjOs
6oRautMtN5l1JEhFAxCtYBZjijilv8KRfrt4S/ViWqiioqd6O8ToE5kXomBVsAiB
ajIX9cGIeN+OHTzonxh5xWRLMoDUYJE9mojfhzeVzRTz0tVL6OzjhyC66tNb5Fn8
g2WOdZhg7RqQpdLNal0h26W7IzJMLFPLeoCX2megpl6xiuRG9PiVjZTJKNaCZuAO
QH/Znmg3EXVg1RReG1I+DevacAWgmGdjcwz55qOKRQ6kbv8ApD55B/I7XnjUapdN
QNm1oSRrm36ULQ8m6kN8rpS8XrNXESbaQtpxDM+Toj5VIxXRxIhf/KpdZxsESpdx
XWFWJ923Z6BNmp6GjEHpS1X9ZFHunkB5ny6fazM+wpLTGqjPgYW71rhJ/tMUlbc+
F/zR0i3YcI+MSBcsYgUSLhGO9npP1S/f7Xqnm9kkLSF6BZnEtYgHnGIWwHjz4A2g
oabzO6GzYITX7v7gTNW/deBM7NrfuovEps3vx8eiQIHK0pD0lU/SDaH+eH7pu24A
gWahKUOpFpRnO15yY7Ib8xrc+srNV5UoEhxM75GV1IxC1LFHNtK3IEJPG809gb1k
60I3IlC5ZgxGAb59RBj8G/cZJ2Hc08fQL0g119DzSCb8LiGNRRWYZHrw//voz2wV
J+k6yFedi4NHSnlZn0zIuaMPVml8XFSBe79hTyatt7uCXFYE+1d4Ff5YWOQ7Oy+V
YxCHO0ToIhpaRzraXrQRY/e4424eRuULE5jYrpym7H2R60UKN94tZ08e3ypAWKqh
zmQ2FVdjyjZ0k9oi0wjeNv+mcZGDFJL6wx5YIAecaHN3r5WTDRJ4zRHL0Jes3ehr
RQMxHOGGi01tNrV+Z4foiG/bRIqVctmHrcODQ1uaodY5gs6smjQr2kVLGSNt9wb5
QJnmL/o/wPEsGcKirHD8WmCzxzhcsqogl+zieHuVehCCAaaSj8zHlM/GW99SCrOy
lTfOyxkZU5SBU5Bu1HiglUyMqWLSuo3p1GOp5aIOq0GKigtjW9rr8UGp5OA0SsLU
OGeag/kn1Bc3lOlCw9MPYN//fNvnkEmu60TuoYutRU8YHKMAQZAjBbIj6azTI0lh
PZodESzzHel8dYUby0OgIXZM5drJCudFeR48mvADzzgEACOp25Yq5oAorcPzCAOm
6TOspjX12o1TuNXaZLplAOtu4D75HFPgPTeouk3Btofe+dVYSRGzYHXAqzLv6mX6
XmoIcN5eFJXNa8UxH61uurHdi5vKUt9BxY2D59wJZcfRF298b8EZBLJlolHQKn/t
1JjR7Azt0iEG9fURDGsUO4ttinNQhj+UwAXG3XXvGbsBuZqAdYRe9maKJCrsz1O7
v/8wP872Yd1IPurMxG/dFjbfbK+l7t/q/bylotFmml1R99qq26yFwbt9Gslj6SLZ
a9KZxlvDMeRIU6lsaXc2BUBPn+6wLlYfAYimClzawQThp4BLL4rf94lIpHoikM8F
im3ZNK9kO2ZQ/BM5h/Dfj0vZgl0GEkKv28nW0DPuJnDW18jqn6F3NQvyV+Bh5BDg
SZLcKfd5YgQEH4t3SwmwGl75rPzLs9sIEuWbPjR2iqnHIe/460cvhOTguYHd0tBI
9Cd7gaVUgopLpc0bCqJPMEXQyNsMxTHuus/Erxe/ex36JryogZHxZoHT3jrdZh+A
AykI4+5llcbrP3BHg54JEFc2rBLauIN18lON+7HTH1t6MPo3J+hYqkF7WWcwXyQu
8++ig1GgpZxc6I4jvohlIe43HuJOnDgF6iEvPsGEck9hmcwaptVzvotYfV82YsQE
P+WG9+V+KOFD47Czy+birdybQnUoX8YgkgvGY60PwZoHWhgHzGEH+nXvg+oZzTWI
6tXmeWvo3QdY4el11sHNW3TyuW7fl9MeWejU1tk7FH/wTTj/EmYX47eHjkGiVUxS
9mjO3E+1RgdazQIhMSlLQJjOENma5+UsmDe+w78eL0AW8BqOxArHB7uZQVTzLnjP
X6e6GIAaWrZdLAvmwBMR3GYh59Yu8QBD8kEEsxd6TCLoFOMz+IDXBXnpgD4sbMEQ
N9mqoXH07/WE5C5pe7Lto1g2BxYpUn4dBklMn7oH55SHCyvO3LjPWcry93CJQ6AB
f5qPvIJQYAg4bNirMlxs9jCALasYL/kItObG9fDML2kqapsAtn+K3BgQfdV8ykKa
f/3OXbljJHJsXPvni7wbqrbaqCISr/pH/1ZZJZttHIyCGOh/jPuOKF+eZV5XxZzU
2CIpxMBlSHjyhQF9xjQRYJw5gKny+6ftlGhXLWvHE5mCb02HRlblAHFqyztGZByP
jxcJU3s6UOJRfD8IjZfeuyh+N1CeyUQSlLKzUz7nHNJle+wf4svSdYa7ez1rIJfW
/rHff+bQqFiqQ/fmn705BZArjI4yLfjo7I6Ka566yldhEjq/rlBT63BXF5x9x/ez
4EnNKdIhg4jixZ0qjg4Wu6gD3/V6fnRTsVpMhOEQ3eyHWFgPteVIRvArW3I2uput
89mTxRNoyEuQwyuKfrlGNUJDB55FBo/+He04DKwbN+OFIgB366Le4EVnFGa1LsXj
+83KXHab7/KugvY1osZ+KOvbHskIRq8mqvLA1R1TW5Cq2PGu66rj7DMZgN4C7QNE
YhjPLDC3ziXPeWM9He4xOsueLVReiRemxbD1j5c7mMcTw/9sIKI2y78C5SkTpcVA
jltncqGTGWieYqGIopbf9zaTAz5FMFu6CHGNBEBtsTI/UbLVfWwIKyxRhZzWdF21
QSSWajSyismN5NWu3agWBakwzw4ualoONXsQdZdRyXqYnYaz68JnEBPUQwX0UcfC
F6KLCEJP7fj62ZSixWR/9rqzP84fmkZ4UVePDLYoMOhJcrYTS6B4xG/Fe2mlpnht
X70RxLZuUIjJC23CDRxiMiGbqImghS63MUGPH7RHNCZYv4eCRUPJT+DAHaFtvL2T
mDxRYCAEuzSvTnZJhtMWrVyJGWr4LvQ9/7zJs6UDpnb65FQu/jh+TUdHbBOvZAkk
jM6icG7Vn8/B5GQXyHbYku4gob2lFg/rqsf9xT0RsCnNtnIy+NTzx6CGmwpzo5ZO
6tqzmcnH+E0Y1Te9qBEC+W6V8L+uqV6x8xgti63E9c2vyegT6J7uQFbjCmnKsj4f
l9vMRqzQCr+DVpZkUBGmLcCB5Jej/nXv3kMUihJTNb/C0B9mnN9/1zJkAVMXC9E8
nmJmopmicOY7EzfrqIEBCyyyZXaCIje5s+gyvIh9jSullF3X/Qg08jkr9L0fjbdN
IimiW5amGgDfIV/MW7xqKv+T0CkjSxNTAU4462qUJwThL3Wx6VqGa6OUZImCWqZD
sobuuw768lYhjaCkWH+xhGwyblfrSeIfQhCr1VGswr1MPxeWBbm9wlk+RKoklYz0
E+k/G+nQiREGZPKnbZsSDIG8m9EdvPWYNV1kSn4BYWQ5jg+xxpQ5NFAyATDY33RE
H1NWP97tzYZjwYc6pMl5YKeZTpPFfJQPMiuv5F6eVtimu2AnlfopNICSYfIwcs4c
xZDKB6568LQZaKGISnnlsO4pkW4tBU9l5pQRu2irBxTTmVv5z3NOBQbRqvC8vd6y
8H/RPn5W+1fDPATcJPy+DS2lE+G6B63TKZmH3r4QDw0SgdQjk/pO2x8CFqa+AXBG
yyWbdiTbCrWmRpDt03BJJjuSLDGIw6WdBdr+q+j5JCnEE7/5R6Okkx3WIR3dhiMg
O49wlh54LBUlAbtRXMLJ8JGdTU6ZKE/7xEfV2kh5xcQc8zt9EtlRoW5SDe2vjfbd
SRoCILaDTnLX320Y6BAJhW5hv6p9xjMzmb/2eGZcBjrYpCpVibJ1+7d8xrXQnWkv
DqjWIR2GYHNi2m91xc1+UBBvb55t4l3jcSN8bAiTeWDK1prIfGHp5dOfxKnbjSCv
VSD2odsGNjJYF0cCYzReplZ6C2oCMkr7AxW1dXAlC9zHqGapirWD+kNEUNGeOU/v
xLQiZpAJJ7XFPxKCFwPBdymwGl/9aMe/v9dGDtgxerwX4u6C3PsMypA7PmVIJ2oL
vKIn6N2tnERcKpZPoM3jAl008OBFiCuo22T20pIwTYXVCGET+XBLav4sKKUr03l4
wzyRKUav7hgzk65XwDs0ica3VbDX6oCsgffdkcqapEw9G/YWJ6j/kMKtLL+2Jngo
Yw1Q+qh5IidRy+TsBpOHVx9ecvjPdG+Na+cyVx18TQy3Qpl+2Q3p1ME4HkfSHNFA
U3E9AKUX5AicQsE2UgDWArc6ceP6ZDhZ3AmuDCMXGAO9Y+PJr9IepVuUMHXlNZy1
X8Bw0A7yPijQkGVPhqBauIC6eRl9kUJRJDv7x5Lb1NgOZ2ZukirBVsLyLMmgio6E
xGuHz+XQyMMsYArEBcSDmCvketIL9YrPpr6waS3UEtaQFLO4ma4GiUiCTtphXQF6
DVBptPO9rAY6WgiGzPpaNTm7gIiXqOSSAge6NFn10LxD6PebBGmC4/XUqQCDjJKO
7wDmFRJRiluTxUCNlKT0eOeamJ2oYvA4lFV3QMpTPughfuRa2TXOl0tesFQ2oreN
I2HWjMsCyQp44KprlXOgSBjmnrWeSYGBzyiZwxSGR4NE283jsWbv61HueYkJ4ek8
rKd+IGahHRcIGHXcfEfNH8XGsFxItNaQ6WuSiiGMEhDwPPR9IE6X4Abvux2wcStq
eddrLjn8kvsECFqx63yo53/u5CjHcdjnpXf/hTUi2+oHDglKAI3g5pwez2DBEJSy
4sJSVXqt/p+hV7hhSx0/zCWLz5S0amq2iILNK38uEliyHVVyJyREZAUnCJ2VzUz2
3nySkZ2jBi/jQd8awBK5LuTDWHwfE4BTTAmZwijuQBRoVfjvIPR4P4+cyuq0rxy2
rC4AgqVr6h9a1DeU/1ykyqnelA81iNvIRmWRa3lvU82Qd1KqNtAXpwb0lfeNgAiv
UfrRVOkSvRnRbwPHxOy/55BbjCfWeDaTCf9q080YhLvTaXx4oycd44D5XvP3kFlw
ZT4gLdGmqWFRAC7HFP72z9z0tRCN+QwmDWHuTwtU9MVTH2AG3kG9Iu+FH2UDgaec
aYt//WZusOUYmRUud4lDYGwlu3i+xj8Gl1QilcauwHiEaCWiZ8NGGCNNackWeCN/
Vy1107cAYoRH6SaU7uhAGHK00+E6clh8cBeiNe197We+FZAV1WHbtGz2FpjR8EAd
6r2XnSQ29ozi6hfYjUU4o1Cgkj/UPVkAjYo29Hgw0ksPgFbKEHzmEsHTVoasX00/
7L9E77VZqZiD/MBHKjCby+W7iiVDxjEwgVdS5ZgV2sBxDkobQp7bGCE40yTl8oRc
rkLm7ZLgzM5Iejcm+My+OG8rag5OJ1A15KwxTAPsjLvupPssORDgbTwKj92yca+3
OsaHhRcNh1V1bhaopB8Dr1L0neOBa6A3Ig8+EV71mhbjnQqi+iflDUPYizeCdL+Z
B2t7/PDUAQMtKjsWJqJ/ftXTe8fhBsJO/czLFoZiUWO1RhUBfIJTvDUbG5hzAlq6
laJLQixEGybtXUm5tT9cH80qKX4qoEuz7DP49cup67QkJsD2XhYVRMLQG+z9uG0l
hF2EnS4076RrWD3Uf8CYbqn1KqKe9YAOmVOFYvkWhKRzBkjK+MjnIki3JYHUpV8B
husZeWdCgX+Nn9J4Az+NVyPR/+N5bxl1r4Qf9k/kxmPOYQW5Vh4+eiZs9x43SekV
yfA5fp2p19MnJM9cOWT+4kJiTArCUTTjv/hF1bEbonaKdmgZ1iBaKjPRZAaZdLac
4MByII1YV4CF/gJ3UzQLd9/bmiMKuxWCqHJp5rC4OGS0uniFCfmFryNnbLNHok6x
vX/U91Spkzx61e5/t9XD/a6dRwKYtauyUCSWtFu8d0rOTS4MHjlibfe6yGY+CsaE
RInJXfT892QDxkheCg1GLEbS1g8B0D1h+O0LoPDEhRFYUedqNF/AFLCo6wJLU45f
G1dzr3iz0uEGItcOpNKJy6FmrD6t4rSRXZqm4MBlXfMdhzrW4+LEUDwsCdSeBDmC
7iX9YEodV9OuiPNS6jwlEjKD3QjZYYdzJ2xSk+GBFgjHw1Rqyx3BcadrerjXHStA
9hZJp8OhrbaSis+PKXLPEiFw9CbGjc3WQ2GvRIyCVzHfnFXqHmTh51Hd2sefdLWM
h6OzZFJGBn9rUk0cIYSUlGFJ6bhxfiDjSe8ypoCHrVpBpnGL+fyJ0CN1JehOGasZ
2sQ6CtuXKNa09oTfYXIWD6j/TIU6E1VD2WAXINuZBgqRIe9/IVk1P9/upJ7z//QE
8AMyFSXmQJ5cx8feKUfGrQu8DHRgu0I1EROTE9QudIFCN1AXfUcmNCGogXvEv8F9
DAXnGTqKfc12HwsGBRSrYnfUiNdpUuppt9bjwjBmSg71fydk7d8vFnTOeyipYO/Z
1MeOxSovMkAlVpgJELxmWRcLc3KfpxkOIKZ0sl6gaXl9OsL2acdHC/xO2335OXKd
ZK9DRcNXTGrZRnjheKqDN2hlSHjb6HV6ZFEiOEkWKh4tKGGrDSLkdCRqJvgspU8U
efDgSzVE7XvAwvTTNsrf2lt+5z6bdhwPi0KXwv4bdIPHD9jPx4znoCAI/d56qN+j
++T9PKl5POy6IgdV/lKyxOrZNzIoKCAP/m+jy2OOz4DBkiRVMr8Kyh9iyPGRKC/W
sRV2VV/eYVrZ0wY4iuI+fxxMqOqIzbvaEubxa6JSzNEpWhi051jGQzINupN46Zhd
Zpeg2ZVmg/kALUMCBTgcSLBFiAqJ7dU5ZIlu7RLCWNaqFUHvBoCuYxuD1iYR4q8o
tXnDgg4XAjld74MqKNvYuJJPcKvdaf0VfAt2clmceuHji55O0TEB2U3rxVpNziP/
riQoEmbTy19T9K0gWlZj9HTUe5Rvj45wliT3AjWR/fG6koWcWDy+lOZj1zuISWNe
qdMePn+gbL8NLgz6ZVprVlCESrUAuS2URTn1qyRMJwpT6RDTlxRN4XDS9EDV5s3m
5UHVIOUz5tKnw98qTQv6KRE+fz/+5Mnskpd6WfR8ii4xVAkFfDU8KSXicKuKJfSU
m4fqkqhNgJMMls02GRDy9igG3VzZlLABdJXOeFD/z+eUCM9O1IjrgTaC26Rs/v+n
bQLqX0HGYdMqcFG5KMU0GwWPKXQoUUgULDhYvyACQdZ66PhfzM+vLFK0GkhOlUVq
54nI0VTiFvzXiSjnXYSL51UthDAammiaGnapT6n0n3VWouCpzFxPWxO2Wj9XhotD
biZU1yuI9woeKkPtcLtdOZw/1eC6sCa9PGRqNe6EhuPX+snfqUfjVGo1LPZKyu7h
7TuxSLb590of2TBVUm//aa0qFUCch0LdtyFcLUS+RA0cOYsSTlP10V4P4feFIbOX
mQiuYASs3eWkvApZDePNP+/h/Y1mARu1S4pdi07XTKocXB+FV6kKbpixcDuCRhVN
Vj9XSdGwZELJ9e2MWs7WrZdfE2myi33OcJottsZApFeNnGoW0gGqblcJwciTJHJd
IFMvk8SnAcnDJX0AGq+Dmpi2UZG79YKPz220PyaZjE1T54IfxfvKXlr0+B3KWIlr
HtiBHmK98PQzmuSVlD+S8YobWqfm6i7Oj2IMvwFf3DA3lMJc10zV7Jt842V9v6x3
IqXtWs7d905szjackuyGVhaEEncea+F6FJuHjs86hbAQOteKIWDWU+kYxPSv1DZL
jRtcfahFIQF79ogxRkvoGb6Tksw0pAYNUPpuHLYZb05DTdNDo82u6qT9PluRTPce
TatwCpM0hlTL1c1yuaIwlqJ3WzODnEjFsRUWFEo/XFpaBJ3bXGiDu2OaOkVh1hKi
foujQBEsviEKDRN3CUE0qIpdlbDhXL3+uMTMNqlyw3m/zxtTdP6Y5g0nSK89dbHD
xnnP+W0x0cvXXQovoCdd0T1i0vfWUBAzfDLfOuqGFRfR4iM8bPkKir1C+1NCohux
35lGM14tIkEOZz1/X9kt4wcStrkVPX2bWa1dgKnRsmDB9rmbl18F+aYiRCIpqc9k
0DunVx58l5D+LUKV+jx2C0IF56C7+aRwFygzHgMtljjsaXHWB5eVPnVuw+eBBGVZ
CJdTgrGGUuwJmrp8d9m1N82c0PS89WBbY7kpyemyaB4EwwZjQ5ZycyzDiceQJZNO
ISMKj4jFihLZrvzdca2MxQgvcaGtKpYDmg6f1lq/NxcYW18OzsWfF4IuvmXg5gnN
9wbn1RjWNaBu59xORToxeLSgcld4nUEJit3RYFI8Z0F/IPQa+wnIuxt0TlzshhcE
nPHyoLEx6bDXUZT0JxpdEQBiVf0Zq1mJjXM/IX3+r0xE2i6rpN2jssjkiqZOKt3F
oWpypxPZmKCpHWLeCASoHgG2Jn4jYi339P8RvprL/tLHIMZRrEdypH7Vk9nXpj22
3hYg8YXULrPX0B8m8YlyQcU5+JFhgMqs3s8hXKfPsgHKpa+vbN6vf6MJHfz/gxwQ
TgPNaKPFkoACPn0TLsSW8Z5SwxbOMFFH6qqWzm5G6o87CTDBsJqm6E4jI1/LKix3
KtvCdzcSZOjxQbPpiZ9CGkuT0C77gUMaLyXeCUJ0iccaHQnZWO95+83/JIqNO+kd
6SiQb8UrJiyprOGX+c+MuRmSIBTQt7CV6TnpPClJg9VJjzSNNd1QMRftTUqXt/g/
Ge4s1mg4dBzC8ZbMITYDFSqxHaMGP0dypO9nJrLhJf5vsRFuFNL/1oWLI/xuH3L1
5QtOpHdKYVSjbsaRjCQittpuq63HawX8qyhx2JR4xlKydGsHf8DK/OwLNP/+1EZi
Rdxz45euXRUkI0OoGOZvYrN5z0l2TgbQKcWcA1pTt6erUkZmL3ivizPyVvqqvFSC
/GC9Fg8YyH1J0D7GYW5dMK5HqE7zBdyis9qI/v828QkFMauPkQwAGN+mfVJNNoaI
xSLz7IMfcXPtmp8MzbriDcBudsx5w8E4bzdhVdRDDB/gi+2vtRBd5olK40A/lgIt
HV21Xu8suiiNcfEeG/P6QYvaNLuUl6jJw52nAx0WrGr+MhuEfIkaDEoP/tN8G2b3
PO3WzhSfGmlgVPtIJNYq3lFWKXpcI2/BfaBWDW6Gcd2FQNn9lb+WJC52cxfHpmnA
gLFCJPHL7C7h+nFRpM9oDZMAIESOzuYSfzXoh/k9+stmrJ6DzU3XjMrUrQJ3FjZ5
UvnAhvwle2TUNipRvDWOxUXuv4ICCc4ncwLqVEZMekSvf5t7q/Y0xdnibqfVWTYA
SFZL0HuNEWLJYgp0Zg8pQWfWIZCgUACdBZj+Pra3HMpGEpbCiXiMsYtJ073R1nK/
Ahbdw5wpC0kkKhs4Y0S+a43H+bM1ks1pp12FaVkZ9sevtq+SZ0gxfvhMeExhWFrz
AhQQ2hXQx1nxhIfBDQph6ptPvmszt8Kyu8Auf0fmquCCXZgQ1APhHkErkW6lqh8Z
sJyxsdaUGm78hmcpDTROk4E4ZlXBwYJiI7kN3AghZSbwsE58Kj+2tj8caGsIL9Ro
VDfQMe0tEl962LEddDGUV4G4vURF6KtBX3NVFwQklGWHAVbVRfYgmzKXOUQoSGgX
9qO8j07h10/Ai+aDW+WjSeIm/qyQGPFniwG6DO3YPreTWFZNl4mO9dGZY9cPL+mI
DlQSlNTMSnB3+jJ8pWYQgPRXVHHuyRYV39OLnqL/a/cjPfCWedHSR5oOwPM/FT0Z
UOjUX5S1T8C8ItpCVneeMl7ErFf0Zx9Y6bBJ1jc6pmotqVi2UMKLu+BrakxebY78
OBIaqCcX/8sObk+DjCMYFVFXcOiMsMtUc3KF0aeLTcuJoau2pJk0ePYVS5GRESXx
lGpJuqms6hqUP19vR+rHutXDjjttN/mtTcag5HeYtwuPR45CNe6Jioe2rJQxB4YK
rW/w1AD9ePMzFmM3y0yIValD27r1QtbIrKCp4Fx/HApJd8rZIAeTduPz5iMogpfq
a1yzUiy3gadQG1++5nINne+McJoX9rBX/GMwtuZhJm0d7Fr9Jtn2jCaRW6fUUSx0
iJztj2peK8S9ln84qdKYVi6GeBFl0/8rMu8SivOSqmwhB4XFPOJW6bt7QWFrkHuW
xqpIVQDTxSd1gnGtBactF2/CeSgoW8+TIJP/gSqFk1HRgDahz6x3aiju938DRxoR
7yHVjl5Im1C+yKnmnlmJs3i/2iWFpAy3jIaya1OVga5kl6+/5YWaFdnNVWR7H01B
gP02JYJr3UTVFQI3HxhphhpOsZ3s7ovYo1XMqTBdGDTtUFervuHnDNa/XU++4e7W
PtWK8TZtoEZW23K0IVVKHC5PCZmY84nUSn80bEp6ml4jtnISJ/aZC2DPYV3KpaKT
hLUWc7toHPazDMBwNVzz94UwmZWKsaxb3NcGNN0ca1vhi15WShshsck/W+4XU0r6
oLLfnvUJbyB83/iOfO4DLiPnxIeuo8l94z/050/RWK+fYsxQb+NKhTs1JYSyazBp
ac2QKeaDbWDwbEaeoTJo2vYUkabUNJq7fYmp7EvTi8MkWUeU3E6x9DC06k0/khV1
Rkn6ig3+hkWnkDF0qveZKHDyxT61pghcmVSUNd5ulKeA1690bQrgt4W7tsb0QH27
sl4Ovj5/FuY5IxiQsphXBoHBuQykmdfDsg4Qcz0m3ShU8bk+V/swBi/5W+hsBdf7
F1aLf5qYNWx1BcitqZSTijfGhaqY7VVPqNJ3qqL5nQD9c4HA9Fv3nE/9dxQ0EJ10
CUZPxQp1unIak85sx8Dt2pqBgQtO5Kw14J/EdA6C91mQDC1tl9JFYx0bh7B0UE+G
MfbJvFIRTNsizyJPfoupWNUqH5LDHQcEBrKLUoF3TvhThG6z+vD6Ov0sN12bLuHI
eFexKlVSnqAnP2ru9fYiQBriYSzroIsSRnDU7jhYgDg2hVaeaaIO4oK9wRN6Upsa
ZzWB9hdOYoPXD84d4Q5nrmBj07PTtSJuP9kFVHlzh62LtBIFAgg42+/RZvohZV4i
f9o3Nd5q+iSW2+0AgWujxkXbK2J+K/KCbHCdJrEavSkdUI+9gjZM/9KeH1jqVAQY
6lfDirS0xDj+kCazAAKUPQ1fSnKnOP+TVgVPyzAii8cW7RmMj3xahP5kNrhnEdx6
aZ0moapC2T4jbdIOGccLowcG24TaL14nhhNbtEJqHCfYkZaP05rWWPxLHfUlok+E
kEVxPLHKqhGG7lMXHpw9xVU5S9dTPnPOn2uWzyD8u3UCHpjOgkKSwAmGbC7La25k
o/lD30hFWyFtswEICZw654qTL4uFQM6wNvA9F+mXV6gQOtsQTVNtOPoQ5UJ2IQWh
BpiwleFBM8nvwLacfLSbO3FlAlSolZqLY3gYcY/XCIliTlcHzYaRctOEeXr01wc2
3B9As6yz3S0SuhTAnqy4pppe4cMBxCsMRKhAxS8v5iOCpYvbMw8KQzNJTPoECEPe
3Xp+cAOq+9CyXFSFSJqEst7mgyWEqyJea3ixzaupfOyEndaLyn/0yohL+CbY6JXk
sgOF23QnNl0qs0if2HuJxsFujQbAD52nPx6kioVZc86iR3LZX0Jip6zQ6zZhBDtx
fEGizUEg/P+QFrv+K2lQfX5RxH6GGLk6hkRHTHG5ADTClXs75ky5Vc93U2mJB/RO
a7njpVlK90rPquEuXqShueX9R99xlHXo84+awieFiPR0D6fHW139atn7LPDg1XVM
UvXtwnl5U+XsrfYZujapgKUuoK303ygDd6F2NdMGudbf6jjs2IAiqZ/7xa1lbLae
AuOWEwNJZjgpsgmth1ClqRxR2t31heotbFrHgk/oVagwLc+YLuZnf1hMXvTK0Tdc
8MstNECCYPbu7vdNpQSW630naGTAn0OzNaquAT4AmAa6ab8AtJ2IDRsDGDIUsHcO
dGvnk4pgjT/jlJPAJs89fVBde5n4xt5S9fU8w/fbdVShE1AjN/ipxtXsKpGkxfiU
gXaijRllwLPkou5Go3JpFjX4bG3wq4iZRDgQWov0faTYF1Bjb41sjx2jCoq6DCBp
O08FwrNS8CbeLPT14If636n5HYNP+poZNCq2zpavMFm90NmfYb2UgGiApLEdF7uJ
LyPTnS2QLy5W3nRoUadoM+GTXUiFaIKSJo2vDtnSaJWjLf1p+mpfovi/0I2JtA4O
KMufopg6gv57VsHuavK6YXGGl1CF83GzSDFwrah0FQqmazcub63ua9hwnrYCQeo6
7QZaD+FF8Rn2EJb2DXRjQj1KBzgmL/eCxnjAqfrUNam3M3eDjswmpuicTemk7WyI
rXRhMTzAAFwdDpjYyMpvCsox1IGzDoTbsWPFukU5hYswfYEsSy6EbZx9kIahWKGk
cGpSZwkSFalvQyWYwIoDbE5DwLJ+Rq4//+AGvSlaWIeqnFP696WRobDZNsTV64mV
oiUIumpcfmFtNapHz8Yj5RH/1aiYxYSqenvKDN4MjeEKmmjsnJrLbyM63FS2U96S
zuNsdphVF7UQZtAFfJQWXnL0yqaT9NoxVvcpJC+0DtzSSx+IsTsSO4rJMGE7zckv
qmJuc09bwarYbsU3SAfeFprmLeStiQ0cW0whmLOIjJtasA6RAx+ek4gKkjKVEzKT
5ogoAOpDYn5NDgU1+SN4qeYu8WOk49y7vxR3cod/yo7te3oYPcG13QTxhJHPWLzl
iCebKYTM1uhXBUFmVGi+aN6Vp78awATbhmxw8AlsbfEvEeEcpu8gsu5fE62A6nMh
UjVSCvjL+eIQ72uk0IXArnPP16AY8HOQ7kfDngfupewqSJNmH2xAMV4TcxdzuB5o
rFNMG7nEVNQhMAk2XHuI7mvd5UHlW/6q8HUjWf8r3K4vdG7sx0v35SFSVjBodHJn
6CrwbU2NmHrXRwjsxEMiDV4zGP+RfrLgqmp5tZ8uLbC0B0TnLS43k6fKTRDOrKcA
8F16XLafsFBma5eEHpkSgbooUgWO+tSM61wl89BKWps/owmEjrQXhvnkhKiXtApn
ZiOGBFmsRt7rOSbsDqOO+YIlamZt3GHGy0VzYvMtu+9tvIIHGvR/WcuFKZXht0sj
ewZClUoY9OURJzeQ4N+JLF5ExtCDtT1n4TTgcHT3U8eXWDJzHx0YlqF4OSc/E7vn
EXfIzag6dyIiH12lJVwie/qmR0Hy254L6W4OmZq58pz3UwcpAZVuzKzkOc2RECSz
QYZ7RR2f6lTOGfv2ewIGimsJbJL6726O88zqG0HJJ1Z6v1G2pH+RbOYuTUUUu0L3
piUyHNEfoslsXTsMK/BWrkSQeAOxf7q0SepXz8uwhM/PLbMG3bqGm1oR07UiGOsc
fLCTCb9loDSEctroROTD8GGt9J7CrP/ZVQYZf7ynPuXW33XG40vExRddN5XQCrWH
mnv9/XJ6YqMjQX1n4M9OfPQ36nZWsvixpTzkRr31zMx8pHMRZ3ITYLytfi1Rws9A
3Hmi0EBdtM7qp24hg4Q95vQTErs3dQU0ptCk5mjkpTvbRjI6omkoyNTFqbd8ylw8
PnoRluAokQQzagehgklzq/GhZELfYYGaXStYI8Gl4PNr0rIkdu1T5E29ozkFjD4U
l3JPj8GegqZpIdY88A/h5uwQkdxJKoqE6fmKCkB8R0kcmE/rJhV5ixJi4K/b3rpt
hVuKtpqP7TsycdAF9SQnntNFT2LbIcemkPL4JLSW0IKsI8ewGR2cCHOLfVQST15I
HMQZ3iwOQ9wRqqNi9WgYKpFY8yGjr14nqoh55Zwg0TvcH5QQ7qmP79mHn1gXTfaU
m9fl91RhuOOArriRSHVF9c/1ZBhWnj7TBV+NOaotOy2+1Xz0UdK7OZh9zfJWA4Z0
mMePaLzecsbTzn4j7S7KlzzOytHXMUH1XC1wQ0/rrdUCcARhRhP6nhcb7qM1a3a2
jdeVPeCQ5xGb7GmBG/iXpJkcVXVnMdBbQjxurJAYp2vvhkQY1QgpXuG4qK0JgMI/
jBLg6z99HUXNqSngrimpiaI/POOmEbPtLm4771zFtTtS/yJKcBR+X2f4acBWO2il
aMMJDIRS/qVa11sdldaQg3G9KnRP3Lp2Mnsv+uRkU81jbvFzUQxNuIPwK5nVVoK9
yzCkTmedd7fF+BF0LNEvVXb3QOsS/priUBMvCMJIlz2Bq6Q8nLL3k05yvcOmF/hi
e1We6Z0H5POUbageIiq6JJyliB+ub8oHih3+B4elbuAdl0DVv94ftX03gZ95VgwL
XHrL+UtHAoeGO3K1e5Y0q18EE3LwQW8iSJfK2R6LQ/k4nuL4qwUIpEn6BuHm0Gjd
r+DO92JRE8J7BOxTrvQElT/jvFAvnE92NfiGgwrfcBjDH93+R7m3yfG2tue10iC8
OP6T8v6sQ8IPWkV3vj7oGDkdMXRyT5vVbskCAlRuqlxToUWkBcdilKFDGvoRcpfc
uLdfPZN6D0OGSEohtH/S74e41VtezbkyTisvOY+T1PrnE9gJloG8V4oEjA4xbEyJ
hGg+6e/vxvk9YlYm2ja3Ohf5FK9wm4uH04tZjUh3IfAs2sT5EkLD6O0IS2kdTwbg
/FDt23WU9oZnJS9ur5RUhWlP4/PNJl6Rg36+B9XQW1zDnk7aEkpFk85ecQJq9jOB
DmfyozcxAjjSpGj8XD+uLXZxkxtSuSdYzacIjIZDeX7uhGVwzIkT0h1UK5+DokEF
I7BrIBXdpR3PtFS1w4Q3G/Uzd7GnlpgQXeT6uj+iYX/qxTHW6UXVxPcW0/6GtEHt
m7RS9Y5E+5g/c2ecbRJtr7xH3HRRNhPHQwplSKN/EOr+Cn1VB8tG46cV46uqjEDQ
xtL+jrkx+jhVdz3yHYzn3xCuc8VY8TUKXjkUM+eocesHCawI5v0CujtrURgfqmyK
CaM1syNHPKAYrm4qKFDyYFFYv5LPfY+2R7uXPxlqBdIuBoxeWeyZq0Rs2QChvTA4
+HdpCMIqaO9b4hKHoPKMp3ZxJcNl7K8iyYa/ZwlvKwtbCH0pOXzTW0F6xfKLqw5H
FfQTPK1aVC7GC47brAobpCU3KKp0Y6Si/w0jlF6tUY78tL7Fl7CDcfbY333dcYwq
W5Ryh7H7cCHyrPriWo3OI//DnOxRkwc3xY7BoPTANHY0OO3JcBt6vUXRcSgc6IFc
gsrBQmO7dJsGVqx2CT/Ty/6zXUUKZNVPb8XIsNx3VzzcMpADLvLukwh09wi2o73u
nl14smPW/v9dn53VAoBwjLp/QvB4Fg2P4boIu780YDT640hDUYsdHAuBnO1cfNxE
+v6HT8Yj4SBQKrApKywQEezB2bymbmffR65S2QohbwF7aiH45iSRYsg171wHE+wQ
eqJxOYNmpcABeKMeb+DqgbxqXT+SrpURWTBZUyzg995LO6gNKIhEArzC3/amg9x4
5OMbtMIsZm2jZlP5Wo7z1YsueLOpKSuwwjpnD1qFh/bXcfXip62t2P+qheK53A+K
07HWx9+dKbgsbnLWSQ/yhHe1VVcnM4ewwN8LiCHv5krwM5sxcUuIhb5p277lZL6v
WEJ4frDWYzJBwljOmF5hXcgb7ZSR2MlBnlXBi2d5it+Cs9tKv/itG+RMbTx/ln47
xVJyurFImQNitb10R/eGc1xPCemEoOi3N/6wr0OXxVmJOoU29Sw1/mvQwJGnvDMF
3SAqvuEkAiKKkXZLVXEoaH0oabY62UkYUtSzdJ0xUJ+5Ho3bFYltVdP2EKFYi1gw
ZnIJvmIZ3UV8q/pW5BtJM+KuGtZ6kS1w+QjC1EmZiNRquU3hM2SGe8NJY7r4G++P
W/NJIBlU6JTcpcmPwBnBwl6FiAMbUt0rn+o6I+4K75UYuNw5vpeQbdO8fzaJwb6l
YH7RgDJwkF5EclDljBWTqKZodH3FjvwzO0Wc0l8CvdTe/crvNMlYlREfXZPfoYk0
mV90X2zkGH0HKfwUXFTeEhbQW0YXXpa3QoZb9qlDMD/Iyly7n2oMXKpS0WEdE9qx
qXL+99QJdK26vKhGiBwwpuYfYNLhK78yFVNTaNue0TIjXw3ydx77Pzyt+BqtZ4XN
Y/jrWjuyKXPQYTna9T4nxqwrsOvGvRUHJD+thIvn/f3HFouWsph66gH98CwMg7Ac
F7PX+9zLEfzwon0vG+1AxGLXN5CBFxzovgFefy8USgsxI8IlC1z3HsXytU4XeKf9
Q+XcgHJPajjnvZKaid4SB1ucYZnU1T5nTt0FoU3ZTdB2JvHmonu3xi6vOYgo7cqW
is92GLzaOI4cRBIhORFUj1Ryqw2tenJJwqjdqXnFNCJ1zz7rJV0Frhi/eb+5uxT0
971gTY82F/AEm5eTWrste1R2ln0FDkzi+xY9LE7GV+lQk4J4jNSzthOFpAa0P0Wa
SFykbq1QKpOkgBtCE1hgh97Q4czwzttniuHydWEJts/3VE6xrWU2pneVKp/Wf9yw
2EYPZ7/ZSFAWpWyUSZCy6gbhFIW5VmbGgl752Omyf1DWQk7x+3ggxtdjH6WS9Jw8
ploRq2cLC7/ImJ1wsqbgBNu40u9GrDJe+SuWDUw+5ucWT8SpaWOJ02bjvZUNWdMI
wk3lCkZrXcuGtM4tlxl3Yc7SdX1vbQLC4mfQPgBKetXxhq6/aJeyv1C7kwglQ9Jv
KPeUztCF/gMBnUk+XuAiz/B4870oVOFpZKy/2+VEHOXUHK3VI3kVGpMkb2Q5C/fC
IipYXwn/6u5OjwRH0GHN3KhSaDnR2PKWoLYW+0qUWTVc+aDYFhZhu1uC2vRuWcHh
a/InqWB1fZD8QM4TkzOI9HszNfhx/DGHig8vyCjFuJRIJ6oq2WpVWP7I9WNZ4IH+
k2DSgQ9rt/Sc/aCoKaakeQTzeXs5PqzS8YwB1t16rwL1cDkXF/Mm9SpwGM83Ee9G
lDM/YJPUWzJaCu7vXivp2lEWySNGY0QgZKhPCNY/FbITmSPSAaHfRrII3TWw81Di
KnvXbj4ccgb8z2x1HQ4xHMkPwPwI7ByRzdmybwx04ao0Q+HCAnWw3HAx8kRvAOJ+
vGR3K7727DnCILsg51GKuvlUWZ1daFXe+ZohJ1novyxZlLNRZw1uRH690Dnixpcb
MTpnb0DOgIKYcaT2A9tCpeil/OziYdYxpsUBRdLWAp2H+JENBAeV0HJZvpRiHTYW
WzmsHB5Nm2JhXtili+kcfGLZ8HVmuSSGWWFYcMWBPVqXMmckN9vEWzWTiceOhYq9
NCbhi0XZsMq7QYOSxJoUnUAUpTEM/lukhGSKDDrivZO2+h8nRlfHW9QbCT/J7v7c
aPmi71gUQ3hfNEFDN/LV57G3P8sTM2yfrQi4105fQdxiAbc8Ximj3FmIYODx7yG4
l1uGRACUL2pN8YSxRTYJUL+vJupklK+Y/B8PwHRwYa6oEfl8Xj8Y4XaXS7A3R5I5
QVfUReIVGePxflggcLyFhR5/0WdauE3QHC76ousCz/vJyj+NX2FwTfn3dTNax5N8
BEWOpzvg9FR0I3/82wbacUAbv+TPaXNvXYZBiRvxyjKinfwF9VZtPneICAm/qcZ6
aAZeXoissr+V7qeQNuMXwwiGIMKuM+gFB6muwVR1TEOCnhH/9nDeD0ByYb+a1y3H
Eq3aZ1VyoNX8/Ojynlu5fk03hTdlK9J1OdNYMQo0h3RpHjAQ4Qw1tLMnUfgn6G5X
r837LmuQrBPyWWhcnImRQJp7yNj0+dUJsAu/EEM9iEqBHJ7smhZ3dErxIurgb+U3
WWDGwEJLkrkDTd/0qSJ5nmWT+iTKIMpjghaUWRYCXTxJ6ju7zWu0aIXKo6266rPz
DvhHSLQLeokF+6QBH5iymIA61cXWPH91jOv+uyCdXBcixOXLYhbQwaaZfJv4QywY
mmFUJ2QuPHGZjJpeK8eaRD5eLef4gSppJTna8eoxvZ6KjxNeM/K1uWDil9VG89QD
+RiNW7zvsoHEG9ZLhGp+mZvcyURm1hTL5YWt1WzjbairS5f0r1zwgUiQOv1eQJ+D
p7xT6/Fc/gs6Vlm7GPqmQEpBSGWzkgV2gfcanxxgE10gWlGHp+hrC+EULQgjn7r/
lVhIL0soUfhoQG7VBJFI/aUXigS7J78igAp3wPXRCBfP7dgzUzsmf+6LIi//6HnM
cEjYlV31SY7CaAHq7djVqpXFKqqYQ9nRWkKOp+m+QfPoOZbD6r22r5kxKYRiyxR5
DdHbJHbetTCQzSZ95HEjS2t6enUefGJ7cl7vOM/qnMIl/YUFzOGcFR1ahpeEKNJ8
wmVy+04uSR0hFQg2cHpiiGM0O7xm9Ke9U9bchJd2EmJk1bC6c4ckKOnJI7/s99Hn
jbcc2GLdHpjeFGkPOLwBF/I2Yp9uWdVKQoqxX6Zt5sYX/LR8Z3FGvU/C9CWuPK+q
qw40bb3p8iyLiNB3DEM5Py+Fzyocq+SHTmbsKihDb++2m4VFb+ZRFMlLmD0v8fgR
fr6bKGtS+0UTLivgiT1n+1tn5ZFrRx1Asga3QbMST3fYwiBSukaL1ZTUaBHk/RTT
fUYlLhB9enzl2OReORWzVM+fKOsrXpTZ4CuXFiOqb5BSV7SD7w8XO1JskPNPYlOH
oE5qUytMWShHlnA3VDNhur6zF3jijo8aSZHP4DR+zpZGrcXvlT/CRyVbtkSR7IMV
He39w+NhbB0/TN3mk9qe5xpLMsr2zHwrJN4ht8hu5Ymz9D21b9Q5YypQk/H1lazd
EK9NwXUen9xTXCJ8VVOESQO2XpDNDX/iZ8KuOUv/cqTPV7yJSjfl1HSAtXM5Zje1
KWft+cZS2IH8GfioaTSQAzSM9/ymmsUKEmB6w6/rMTWEAY8Urid5Tbo9WxHQFpbM
mGVEpHNOY3Q1MknWgoLmIRyPNuKzaO20tzVMq7uGoo39z8B7seuou39aqfY/GCR3
jRj662Pp65Vsx2RRuF3oYd1ebQaKL1WrKnQVCYDwDf1F2/76vgPY5nIKBC1Gk54k
flYg4uFvRIUbrAPKQSJ7NoDwbsnTZqpzbKzVG4tDuqTHtN9clKcPBZZubnSPkfUP
/uyTbIaovZyDJGvgO7j+tw2RM6U1emGaohrwPBODkJDIX0OfGEYJxtAIq9DAoi0q
r7h+ZteUmd/Bc99DGxNi6lwP9GDxf8J5gg9bqwI7cfPWEI1JNmcElp37frYu2rgP
K67D0LKyxtkIX6JnmdrpykDkxtLRL5k+Xu088XVuOECUflLZCwAaX2wkiLX05Oaw
7pEoaQ/zJRPalVeL5eV7bWr43kFPuZTzWsicPHC8TW27peTM2G8F00MN9OOq/CMn
4dED2DAsbC4O3KjxXAFknHAnl9jwuiIkUMuY+XiN4hl2W2t/NY43MBgs+CUjGCpb
RzqYJGFKM+HPnvUbsXPk7ShqwgdmCzB2uSaeq67+RwvWB1r5p+esnTK6rNg6Gua4
/k9unKgXpMv1SzGbCzkdQWFFhNRpu94h2Vlt+GnMNk58PsreILo3Ujv+CoXqWHuO
k520mSPQoLHG+7aVP0PG2rEG3pvFe5mTYOCMXS65jiGDMKehuWCAhIOXO3Vdfr2E
Dd5pJcQjrx40x8VlE3ZNwZW9FexYFQ6OvUHQ73jNkmg516vARayH+b6ovDoscZh8
0oH2ZEsfzVJs966Q+TKETgGcxXx1sFi7A2bPiY6W3e2PmRy2EqEx6qukxaR1VK/j
M1uGyGJR8YRplO1tHRxuT/Jl6uZt/obSL8lpo4+mbPIsVKM3/sdZiLv+1jEHFkHq
4W9LnDf6Zu9BZpTW4tWc+Cu/Mr6RWzfIWZhIsVXvlQk/FXpiTOYJClyS+vPUDqBW
//BEAZVy963RSz7aQGcBWrw6uRBK6zozJ61z/3JI7FFROz/ImnK2Md3N3joUdq3Q
FzQoSTJ/U2ffgCBFRtuIYE2QV+vGxAX89E9w26+6WR0juN6YGGM1+1mXxqE6aTiX
RDQrKcT0g6QSmnzQIw2fJzhpP4DPepMEXluTUVqBtjIPr039Nn2/lhI7iXdnC3Th
FOfY1VFlmEFPag1DUUFrKPNm78oBsWYz2UTrhQ98ZjtDd8++JYMV4gwuTjjwnLol
YjjbEZSiCN7J1MCVskx/jPqSiDaF2OfNOEVLRr6MYrAiGf9lCZgIWLVS8kNg4lk8
EH5ML/j5arK2rlWmIYgwxdeH8w4Z2ScG6GytuOcz5s07fWhRCNnYeJtBAgottnU2
8hj+jzYvZTZZ4bgHH8PVFbev+T99LN9lpV6ddlolpS5qMzzmONqDxWfleo9O3UZp
k+fL4un/JDwweLfImh6WsO9Gi9fmKeboJdy8QeNjdmuo6RERdJpOc8DuVjtfykk1
fhYe2GuNXt5gNofGid835sJ73yxhkW4eTxQtUTfb9hhkUc7Z3wuANHivcPj/Bf0a
VBkIU/mFlJH+06q7TtK5euR2QPY34rvJJ5H3tQMOL7JAGw27cRuSawthYZUg/8Hm
hLoFIvet+y3KHxbT8qnfIVjD73+Vid/zLJ3CUKPj1toFP6UUygOzeM7+wwdJghCM
jMODgFWbLaZhNZkuMtD+1OI6XpAqHjaGBd/sLniVYUoQOJCnS+tt7Vz8p85CzdBg
tSDvxSDEMLePjRUbWaG9qGm3Kwzgmnme8kFfxx/yo4MFFyuctwC2W183JfuBnP7a
XhDPqwhNOQ7oWgKjthEHC5QPfFk8NAolXGVL35hRz24Pi7pAZJjEOoFO1KDGrQmN
SRUNTCyACT8Ev8CL64hfFm6qrvPv0AeKRJoeJptHeT9pDlt5Cve6YXIR+oo+Fs05
eeAz+G4EV2WFaCAx5qXh/gRijs/jqXDBlgO3eHW3O2hbmnMQPQzCTwIBE7REzxfI
skwqZs0T2SwO3MgaEXd0Nv09K54gz4fAV6pymEY7Re18X/F2b6EESqKFdBXZhDo1
9+b3GoWt7l4GrnyZDM9TYe3NcYAHcZ1UZ5OF928PwEnSxWZpOHnykWb0X7dAUgN6
5j1YQwkFZuj7fQ4VXZAWC2JpHnM9HQ+CCMPF4golyxbgaDUEh0+iQIRcQY2KXQMq
UUMO9uSa5Xr6hOmf4dRXXfv8V7c6YMFQJqx2QT8XiiW4r75Orldffrw1AEKHFT32
l5lmY84M7qCsgz1wUrsfPKLnaVapNTK+dw20729eJaTYW1kECM42QcuRsoqa0eCg
AFwwkmb0JHXK5NBvSSdBgu8+2zlc88FY7fvw/rEzeuMj+mnjcwNqYqjQpOXBR2zC
prXSthHjVOJtLtwx+SlxzZXyVz91MIxpPHzUwUjqjDPalSVFl0zF0l8ACbxkRAqX
z5HDnc08qPFThWbq/lmXwpH2m6rSG30stxiou1vwOOpU6KMO0hxOeiAoc7B/Zbsd
giLYSc7wu/2ThNIUM5zQcvqljekNlpas4Bys3kpVfhEUIGI9kqVzt86vDYggW183
LAYfIB26xUCB1BsQoLHt0RyZ+LfcXQZw+AkGT+BE154m6uWBeV/v8rlmIVV5REJj
Yy6phaRDB2qOP3Ol4KZjQMZ8Wa1gOdaWkJGtkXjfT3TAMjGskzojMzY8pTxlQO57
JQR5BT4ZV1rIzgPk/FyzG6kOrd/jJ0anfizthpszo484ftLNFMe0izR59G1UGx6j
XFA2oH2dWPsXuBdLde8baaRZQ7Y+FUUmKXNI6wRlR3n4GDHDdmvrRSdBdyFUH2ys
hB5JmGrroXcjBK8hqbMwGwpLfli0a5ug3eZH1q7aJ0lSCxWb9S1wR5d+z/f8dA0J
yUTqI4OhGQsp7459PjeiGqYJ34llnUbgB3ycFur1Ec6Q02IK6dVwBuUgLCyFGcwy
2iTt5ucX1AurwxXmyXVXNDUDPgqSbii4D/HZ+bB5M9XIHHYXwy/n8hmxbRQGMktC
BqaDYpK+nB1dMT4IiZdJ6reT9OEOfA0LO4CL3HjhsmgI1Li6Xs92lwf04eJOT+L3
42JVnVkdqCXH1MHsklNF/rrvqCKGHgVHiyVnHgyHwGWPDSZSK0PXaunbdvwM5Ef5
uP3CdNkgjS6VScJ5ZYiUAktSGY5STZp9V/Xu1fbg0/CXLUoOB8DSOUi3nVlYkSqO
QOmw+pHBrLTAC9ng/u7GFHFrr9Dfn+WtOyt4mFeGRq1AMh1y8vK0yZEnQ1PlkNVJ
wsZ2JaTCZNikWfPwt/mYR/3p9/mVDMKsngGeZGJ2DWHUQN5ut540Wl4I+VNHr4A/
Nn6V4sfATk1IzSjkeEOTm4EmSKKZhbEwGwlMqFVDQ06PLtWEzktokZY/0ajxu8vX
CrPz2w+QggminKYqyVq07RbU4TwVaJye8dACkCno7196h3AMv+m+NCxJAtPIO20o
aVm0+DKt+Q/Hl+O9phpeDGBvx521TC17TbAXC3mNFd2XlawbQgecSi5Is7QAau6o
opsxqJhYeU7gTIm6/l+WGe3MKMe5/G7KbSkRRRdUXwStBZelNxiVwh+2+4QPgqkC
BU5HRQNnrvj8Tt0xkISRp5xkZKOqKsdOkNlaaHvGcpNp5hf8OkGEMnAE++OEcJK1
Za16tnwkq9GtKf28itGzb9+gmT9JxUXfTs4b5ZQVSJ8llTkWonD0s6w8Zst9YSHY
n2wFFAyCX427rOLPxLjYTcNC1Ee+sWuRoiZogRXkR48fLRIIspej4B+y5+tqFmv5
HcH6EW5+JZzc/kYdy0duLxBLoRoK+al796gEyhq7KIb2Dq1xD/HtEX8jEC6Y1NIc
40lbd0i6B+HEICsNgwPiRby/wqgicJmn8MVBj9EKnxVYqxWTnu+cZNC+13nbRm92
KUr3cagZRnWuX+k+0j3hsJffuXt4DQxWqGWJrcPbmLs0/8UNu4R9CBDurHE/iOfw
GfVKLz2pjFExHa9wR7mf/B5KMMEfk1WKbv+KPk2gbKqrptfIDCLG2r+VM6c6bQ5y
kp3JZZbkVhhj2dlTrtkrDI7C8GUv20QDbkuWpDqApvMYN8p8MSmViG7mzJ7aYeJG
oIQ/CvqD1e3GvST/XxlsX8gGis6bA0Qy+BWbCBoW7buuUCxY0HMjMwF8l+7/aJZQ
q35fX8cwy94NqXkf1IynnYpOzdFUQyemJ2pTpVLDMBrztw4on6L6jiuyXpE3VIM+
rXNr/EkNFauex7Qtx/DMGvAH6mwzXux/51vQEpJu8uMeF1lj207bNuv4BNOOUV2g
W5xRqeSVpmuN1X4uWYYkjUDp1KzCLz0gCDpb/uqw6ZO1e6Or1fIayd+1S3fzKGXL
dk6EI8to5KTXK9NNCcJUqAouh29UvjAzeCMlQ3ICs9dBBiL6a3zrhZQm7paip9gk
wSoWE7jQ28z0063azLuPt3goR6BrYqWZ8fywF++2THXchr5JufutiCA0z1VV3sbQ
uE24u0TXO3mOr1g6koh6zgAeU70mUAJH5SEjbNArgbBCZDO5hjUCh23fy9W5GUSC
6VsFBo2bPVXYDsv8zEcBOmOSyr1SLHo/CVUCszOOmwF8NS+edjStXhNiVxOB/Ynf
e3ua96X2jjyjVfLNMvWQeh5YYgi3bhCyUhqtsaHYVWuD2vkYf95SFIABbiU2F7ro
DYjn2cnNvD43W06/mmCGMXcUCPNA/s/vG6qWE+9f0UPQS2Rse4IuvVGsMP1yLBig
bnXyWj/tyyDznuqDD9zQyECE6AU5QwElhKuh+3hFPN7Ne58GveX0De09exKc4D7X
YNldpHY/47+5YFVfVFChOf0n1Zlw/4cmh7uVl95HgsX/nrxU6kFJyMew910oDRJg
2fuEXKe2XIVmhRy8oANgwpYTdHYY2Ah7b9BZ+4evtRbrn3clCFD/C98DnEtCcwIO
PTefSo/VGgxAa9jChVuxPnp56/gzvPaY9RdDJDKpyUlF9ox/tqLPcIc8uJD+JvfN
aNTO8RMMkJs+ZoXSs0tMMOGUs6KfJQIoJ7CChre0DsG8Zb9zsTj+PyQpbCxISyK+
EsTQyPo9oZEfic2MRllruARJ8Qt+8NOhy5OVibb3hAuP3Q1DeUrxJ5R1WG5m2EtE
1AhQxsADvj3SanGN7CV8I0u8vFlZ+k89GUeCdJkOcVuD72fJSm6EMVrgf9OBuJpv
lUYddj20AE7v3oYCV04Hx3qjcAk48wvGH/3bn+ZXF7b5U4s97uM+HRvCyTMva1re
rkDzIWMaNF8CP1DS2Cck9tssGmGQebsy6nuHIYeRrU8NsZyR4B21isl1BiZxYIvL
SUahf6LqKeWAPDzlwh1vRcKLWTAY0F2vQazVMF1KKDdBOIzGtVgK8GJxUeG0V6nd
qZR/rj+Dm03QZogHG4pKfDzb7nV+UG8Lb5RUeMYwcVlHiRF7f1f0UigDV56somf0
O7FeGJgu+HUYh1qKHjpLHjpez1bR1Buvd65xuqFEAtsDjS8v3mbCUO62fPzbptlW
LC/zQcaEExCZ6OBnCz5fIZFObTCAhhY78gB2uThPgNulCWCw5fYUP/BQFBWUx9lo
qf1dRO9LIgGqACVXBoFf033iMY3NfmezX/Ts+zie1k9xhIyDt5gaV0hG57+eEA6O
Vz7Du7tKHwzUlseweQjx1gicyXLRvOZu/HS/4ErdsrTtESuQTjN1W5uLgofB3oS3
G4OijhD/Iy+SEhZb1T5bcjvwrPCXPwcNkKYZvyAUBLQZoqtq6Evd2wnkdl4wsViS
AYYmknBnRjQ8xKZcoZ2kEaNeyyu/EX6ZJPY5xFKxZEa3RrpUUWyDjMeDvZJ3EAqv
oQ7ut71jbHS+zKOAkke1b9zRDh+TorXNzE3GuzNTjsVwO34Ch9PWYkbleje7byhn
qVoonVz2eLdni3VVCgKoUKKrXNv8crjbjFBr/l+6qOTE88VTM7YWQmNos5zT++Gp
sqyfivPehJhOYaW4d0NCNuo69EIICn+9yQMiouOp7On1UiXN1T61ASAoHC3QUyok
mqPoI+bhMr6ENK0etsW2ESAz/UEPt7hhebHg/fG2Z7hw05/by69Za6ft7z2NpQ2D
KBla5fCsn7uxiSWUJy+B+w63blMRa45Vl3tWlzqCLzJscsaz57KJDtZCwot9wT+G
CggWXgjnxgNq7u4YPoHzcO82qWKhYwfYeGCf5SZGR2zGCS+/lZawCWtZMHeHCJAO
wQQ9BtkConAl5T2nNB3PTywKPvtcWs0fJ9F9msspExLfYH8bF+qOwmgFWtKJo3lq
GmOFw50H7ewq4gPhnsJ6zM1cc2bjgHilDeIM1QKfqQFOLN8uV006feptTRkHaiio
i/Ka75aP07EKSYqnECMTaMRuUk+6FmcEagJBI1X29C4eQ+9p7eAtcFiYITAFLRQ5
qaod0vfylm52NvNS7xAJ3d4gY4B4P4hYYL7PP+MfK0mposYkXELpPM4QfrUUo2Sn
+i1A0U+/f3u1Qo3wl/fOFejmkLGV8kThoFCBRWwZ6IvhvivI/l4awgcwYyQS7CTe
/HUJmnx0maPxOxjVu9gUKJVSlgr+ThF9yW89XkGTM07ld0XgADuYWGQ5FczxkgVR
SJ5qPDlqd6PrBRfUR5prfXmjnVGzp7Hk9YhUWZ1sJ/N7azJo0Ou8hEvEH+A9pijX
o8mEW9H5DwCEDFEDWqIliFaG9zdkNzJyAMVv5c27J+ZSisU2RaFar5FulzmamxNu
Dysjc9YxkOIauvW4SZfp6TW3utF6rTkCZnNJ2jDUMQla/zz3NMWXK/4vkdDUrCNT
hIzByvwTPyoRXdWvE2gZVImRvqFpKy+NX2Q9RpNy0eLhqCjhh7i8Vg3fHEHb4k1H
eMD5djWTXoH2ShBSJvX9xTH0KvfY4wGfY3X/cruaKLCriEiPmj6yllI1xbrlMwCH
LDcgxKOqYB0ZxZLQJZIwM3nkl7DP5hGm+SzRuUbBps6VTB1asS3T5ideplrwW6Vs
TuyDDMhLhF/gYaYa72Wu2kqtRoI0CsHubp04uBP21znwcSuDzV9CmEC47mNZ668L
3mvh+pqt5TT9MlodCopADtZcgXiEB3D8WeQpZaOyhc29OlYe4azjZ1CEYgA4ttJj
a/ZoD5j2V36tsjG3lnclDWWBO8YsY1Yf99DC8ctfZZnyPvAmb2tIIhzmjRZ7U6tw
ncor54lGTh3Q5wSHjZ6VWw8x9KYOsycDF16CVGqugo9rbo9gM/hci5Inm7jYT/aX
5+AxctYAfF397a1Vxg1z45BXf4QEKRYxZXV+NkmSp/hCXweERNexdkQ6mNxVM7Kt
SUxsBRL0l2MNtxJcyEJxGWf4/Q8gX/j0Jnhn+sb/kOoegSHItD5wC8jMN/HzWamE
lCiyHGKKm9wgQmSEnrVjznxpIGtdUBYy/AmhLpVUkAd2vxeuCpxg/p+DxBOJ0ANP
j8g95weB8C2bnE3OphEH1Ub+S9VAUje58zjjeXZvJblYwh8qLlb41LJ2Hpfaz+dI
KnU24b/S6WGgJqwiW+088o1Dxrbf1C0Wlyx1EumCTFV00Am/rlP2rAPFYBKO4Cvf
3SVOWl06IVRu8NnTzLe2CLuFe31mMUK7gysFcR5mNj7CxCojCg5kksCE5K//7IVY
/RUYoSB+xrCBG+jNxqtLIZ2bWfo69J99t56UneQXUYrhEPy0brxlxWv6zC0rA7x8
/2+oZRqvt8O8amoVL12XFaILSarCkB64/qIbM/pQ3y6b0qpa8y84hranjAsp+CSW
Fs56rehZZdv8LXhxomTBneUpBeBAYcLzc6/QQ9d6TVmq8bgH4E7Qb3lGyiPm1+j2
WU7tj9N2L75TbRp+OFUdGArxU0Io16m55JbojL3/6PXYgvY0M2q51R4/gzThDas+
Gprd3cYuMs9P6ohGIzZgYo8CtG5fslXhSX62PpIOYEAMkLFrX+7VUcKlY0iNdFPR
PJXUpjKo7f3wDzf7ETpTG1Cn7sK3fpUldEiJSeaPz1+NyoYGY1vhnEEIZHMqwUA9
K1sMm1EXbGNfpnYiKIEegh+W6UJRcJhbBLMj/FSTb7oNgNrQ5T5y4Z9l9cWtUjHd
ImvgC7La2vj82PheOM/HyDIOP2U9XoVWAVwC+sGWxsPso3mAxY3xHrvdtK0VjRX8
ub8k8t/OQPCABjBGz4z3Jhtr5kCWY6yIRkfYfA6MBdguFjgKRVpzObsEW427357E
bz82cjKm6baxlpy5vLAtteQCOwjnwFS6UdAlXw5yhDU6CSXJr2NNC4ZSVQWi3mpH
m/x023G+14qTbylzBUG8xZVmVbEuoU1YkvfYzNEg927pnQGlr84vaF5j80Qk5Fbz
y1mstb7VsuS89G7IsQwEZ+SGQ6PsKJheqNtB1cghkNofWELLR++9fpq6dnnEKvxF
gsh7VU7aNEB4pmpQaVdtCMwixB8h1oVYIECCFMOdSjUa+hTc3pmdOn8AuIH8nGq6
67TGdE7kefvS4FCVTmT0cD189tOPTaPAmE49PV5DdEzeXJmwx/q7tkV/q9zZD6yF
CLCTTRJXaXD/U7pVTLLO/QHbpX8TSnfMn+ZrbDzVuxs4JdpwAX+csztKQ1SPqoaD
ask+Ofgob6GewWprwrfsW7NyUup0y7ly4uFVIMJa0yLCmFjUnxU01M7qWUG5tRML
GMWefLe4dMWwJrtdVJTNUbB2rOSake27puPFU3qrMhnpQV3u7Og2Ppi0baV3MtO9
+eSG9QTOkCh1WGnE5Z4H4sqW+VOoa0Yt/0p1tAiBXu2CJidiSnEm92m0T5ZFCY1F
lmxcKYD3I1z4TWndW1polwukbo65DWT+OX9SNyeRbodcKvEYrup2iEriz+7KH9A0
tB22gEStWXuysKZUKGVba/ucNTxNFlx8ZuhkTLzSbqePPrddJE+6mva2Ymoy6dyN
g7cEQAglbW3miwCShhZZrqXBGvqZ3V0ejTuGLdRocXWlPQYp/bvMDM3SPlwA0kpg
DVCTlFb7vSg0xEcyP4P6pncWduWwSYHChb5ZmLQwitljqC6BEFE1S85z/u5u1Niv
waQo8HT/ZfIVmSyS+BH2fQju5NpbnnbgwWkJ6P0ohKqan4+n6JZk8kf3pB54He0+
DUesoxYwWO3c+fGSs6i3R5RIPlj0I3QCQa4i7f/m9XaKOXditbg0/l94LXJtkdFV
ZTCLJyzhq8u8L5SXdG8JkLiIA8aSjOpAWfXoZEv+PA8MZ2tHZkttPOanlILkgz0H
58zz8sO461jEYqeF7RqqW/pkRRVQoVM1a6e9emtthYdPHMSvhjlSeVUQifrD5y3a
a7UF1zmZZrcXsrJofPFMLTqefMvgSO5plhz+fL9jczu4dS9JuH8VTQxXRjQ6xgcm
OiFJKFrVndXXd0QSSQXcOR8i89KYfgh4BiZlJtKXmiXTCjF1q7vOc9JF/muFRw1Q
P/eK6iPVI+/TfwmFaM9HxL6EFZhbYbrcuFFTkmI8yE7I/aSIvI7ayBQkTNEFWVnA
wbnnDWgSt0G+O1r9SE/beMmCEJl53CCzlqUZI7VeyNonZg8SWECA8hYhZxrYZh7R
yxJ3Eh2gmwhbUNllMtosHKs96GPWUO1VbU2MBxefsFlrohpsnymFtVilZuAbleM8
LcBapamcww0gSX9SpztHl/RHD5K5CHH4sgMCyGI3nNoI0o3wGGQMDJwOhaOXsCYM
yA+nlI36u2tIc0BRL8iGiztNtMpZQneyT1fOuZBVDJxyKJahAhMISsg6eWk+XqNd
8KXxTftUIMz6ypb+59Jp+5Pk/lSJumVGDSpMoaJbaRItaILOicH5TyWNVN35qOKm
57ydSyNpl8SBonvZbLYHzr98GEAUwVHiizG7w5PQnVx+Uf4uZl6DpVTfBfYRPyuV
rCHlXiY/z37d0hALQz1MdeURWGGu0OQPqhG5tCG0ngjwGqHr31oQ67dtwKoMA1tl
M8E+fU9AO99lllQhmLsVvCVTTVMug0hDMsQtaI6xAMKkSD9ulhIIFisKYk/u0G+m
HL/07onw/svMOh8hvbG6kaKRVxR9ZiBDDMvce8KwqjD/h2wCXRHrWOZACJA9+FTz
9CCRBztxQzUBubOxXwFk+HXJicwEloBC+ks3h9CjAxo2SAwisoABsvLSolSWfGON
n+YtKYh4ASe03X7rikMPKfo5A5oeMgL4vlBWVTryP6qNpvfBbT4LM18Q8PFU2DkF
oxTAB3Zk0gjOEipiPEVu5EHr00sIu88eHTOyaU57aAwai3IH5IzddyKsSEBItJgu
6IcwQpMhUsdNiy6tUBRKG5uOZpLZ2cmh130PTo0jIYzebtT+VEua0Nl/gETuVIHC
AqfKJF/aQ5te/HsuH9NIjCh/TCTGGjMDQcW4+qM8d7R9NI5pndAospR0va6yx/Vr
jLtYtpMZ2BIKvG68Z6S26mPz3QcRDsu0sTDxQ8eOjN5BxpZ5fH3pTtOSpcMxtS+5
qRBIxfH8iWsUhmqgRb2HNKn4+hYO72iHxB59RDAkq+qwwfpr3V9+nZOtmfulP9Mb
LMW5PLjohC613N2fxGLkKJ7ntzcjzS8HKqoxcjNfGxXmNJt/kTc76kJqJn6t71BA
F90f6Ce+gG6T46qWOFOksj8blErpQzaoHg0jYSobvJDoWqGL5A8amKinL0pjYg+O
ZzgF9ISYoKBMA16flNbFuldCmvyZpMbwEhWLhcTjAmYG2t9DNg+8oEOSZMxWGuPp
lMVSBz1tXyPa91lgLIsdNplEACrldtVi2PWHdGy4FfD+HwLcYyy+kRzvXG3AORv3
QPBREJWqd0vRwkiqeTUP3o+NYrPu43PkvLClYFA+Tglby9CcPwuIl9yb2WbMeFDD
BTG/klnmNSOpKSDUJo1zRTkA+3TB6vxdAIYLd/FIL8LzMLwR/goy+TqD8c9UmVCy
TY6dvik1IomA4Z+5MR6Rg1uyKWShrD6T+CiWFkD5BtYTBlM2pBPNX8gUu8uvnKKa
b5fYHr6FyDaXgYN4WWKnTemHQLizNC7nTFOTyVa3zfRPL20TzFlNHe6apwpiqHYQ
fD7wwPW06WFHjvP60B9tpIC9P7j25qxEDKNHa2TYXBJFY+297hed6j9d6n4Yoe9+
lBdy45evGOXAikb9HYfGV5QQyiMoYd0xHwZpzFtVy65bTa72VyYN3irAbfYKbTRi
V9CxKmkehA4+bI5Dif8yT4e/iJ0BV9lCjEaSlsFLfvKduax1fpewRVKaMwAI454X
bpx5at4Uid2ftnJVKMqNluzcEMqW32l0Q9Ed7OBk52dM+n6rYHEPP0VmYNttcMHa
CXyLODbZ5eF3NP+qqDKb5VF0A8szePHdoZDGkV6L1xO/KkiEL3nLvBEAUDPnNy1O
1vIzV2mMj7ItR9Pq94OVG4VQ7kMzFzlGsdJLdtFlZDzwE7CHpd8qjPeXejsCb7zi
KUPRtwR/HFfqlz6MHqDlnZMT+JfeSYFlZoi5h5xNvd7rH6jK9Mi+92wAYPSK3W5G
bc7h6OKiMq4asOKr5rFU1N0uZGfOkz9DagdGpeGUwfaH2VflYKW2AfIlduLyQJij
e1TB0rVbdTd9+wiVbcuvPtRyEH7ypyXc2WGEVWblgHTE01zw030FOE+hZTZ7eh4H
lGLjufkLEWK2GVuCPRztRr8G3E2dn05h4TYJvlvCs7Iwr3BsK3pnfgz21tOTBPlR
BzIY/6i83fZS2+YkRTqvgsZ1IEvH0+1H3Dh2ExtImCyD9G0yf/1aEBnS99uwrFN1
kVqz+PHn9VtAoSTqbH+XCKMBEekmi+PHDBipVGzaWIQEGqly66a3h1cqEuyyL0QY
cGUFeKiC+L322+23aaQNLIKviGDALqbKF3SHtIJbjSyIulZSK/2fZ/DBSzKfMxyW
g3ePDdsKLjxw2CgSl9MoGhpX4WCOHdkgUNx5AVanIYAB9LS1tGgl0LhpkIFEQ+lb
0k+GSIz9Zm6D3wuuVBFkiHzs+7zA3HF+05BmjDcJABKHgtOomNFi02i8aDa0eDlt
QjcKwDwpU4ingDGZggiEN5jyTradID3TZ0HwR3a08sJXZF1AfJS9FUvSf96BPgO+
yreL6jEs7Z4bM0j8lPcdnY8m8YokbeJGQWnntIbAF6O3cHPC5mQvLDQMs4gi2QOI
h+nPzYS09DiCcQ7/jGuo1Cg8EckN/o4jB2AIF9KiJ21/cxlUaLcOckgxgDItQz4l
hYJDk9fetgenvC8T9RzTXf0m92A6wokNJgBCfQurzuUnFBvQcc7IAXnbUm07Rf01
n+qZPkVXMBTV1LXKt8Qq1gzhUUXfEm8gDllbb/pIlLGLvHpmGieS3ODEyH+DNfAx
Ec6ACMZ+OzzILtm7A+CltrwqDIkCwvkLJ5I5pjtV5APYaNlfMDFPx9jfb4ipFIA7
eX4TlXRdiKe4pL8WHkemdUUfgSL8EIzka8P/pwrk73+6Gac62JtmSLV0vGHZAEba
pLWZIBU6XQgP+0/WTksmMYeRLYquwOciea+MOkEXBUCbp8/C3z00FS+ba91hNzne
ww5U8BkFK9ceCJVxW6LSA+/ykHw/FhU2qZnN/aIJZ8KcwZcTLZCY1+7wkFFfv2Sl
okAuOVwXX3sNiV67oZ1S55j+lNr+0ilNumCop2zrl0MGFUBS/Z0SyDwCfchia6LE
IhPIbb8wimLG5I1lirDWZpoiWFHUzjsEvl1rrcuc/0aEkSdchY2k6re43uFMSvAM
D0FTiLvWeOqGf31FMq9GH6wk7++i6jyaxzElgpThccNiQip2rhOIM6GZqWM5Lc2w
Ym/6XKCyW4+IN7T+aoMSw/hEWTRT/OQCJIuRP5hUWtRZY1iuAYpHCpGdPhuQ03hO
0e3IEUTHgh2JGYV91ssWqUn0dFAhH6zbW2C9DasCCbeYULIPJtJgft9HNEMbMG41
kbOJjttP79e4iCqvm+ATEmbENAKfoQrULA5QGRb/0esCSRdovzJaHjSn1VmBmucS
+wlyscKtvDm2l96tw7RqmINL5X7tdcpYwa90FL0oXTzI59T3mIvembBRCuqgRvAL
9FMFCjijVRaGRKj4nuPdCyligteXxQT9NSZIFWWLzvu4npINsCaQ/4aztpyeT8CZ
Oqw9jCOjVme9njvifCRaNqS3Nye3bzAz4BFFgKBQOgzQDTpjas6TAl2K6lZR314O
f+jZlsXjuVllWb72/k+Zdib6yn2r25r7vfDRC5nemahgxxfv2OmmFIYnzpkkGwrW
KM+DDrQ4zhvmoyoocNcH9jtlVlrJd6dxTf0d54ZCSaJ0rseuI42qQaUHpMCAO7AQ
+VlYBqpYocbH6d9Th2NczslylsS9Mt9NGWOZOd8excpaob3UL4MKCXyH0vbdBKbo
ziYHNAmokaI1++/LmpGcos44X/1PF9+JFcX9LB9NKrsFPz2Xp+RsyfE7PxrYs3Bv
zAhOyIJpq+1+PUAGzpz+dFR2wrCzovi4MKNsuFeA+j99/rAHuxwqRfAeydnBzV4U
pRfAAsl2lRKvbTf+aId5DLk4ctg999pzGtGaB8xQB1ztCCh6C0o6fEhho+h5KaJ8
PAi54k00QEFtjAl3YsgUegJtCTpzA8TnollBwKJz5YPtKEAadnM/7vz64eXInf1d
fw8xK7JCRRKh/Sag1TcbD7oxqngFnvfECPrJcEFYU4vvnMpGjfF/gqo0jHCouE62
bL0FqmDPReKrDI7Rdtsqep5orma/8gFBV7GEuu9J1kPLUZ1H7VjYdvTxTO05/PdK
48rIe7Kx4g+CZXzStu9AmltrS0hNcZ8sMKg5TUXTz6eDDrX6qXgoSa4YaHEQJZ2E
K5wzIZNUxT+xqY8v/SuYeRH84qY1hJoeQmCIOkeV0aKp2oB3Od3cPVywSs8bYNQi
k29t2AeCacMkTWW5yoiAa7kVvB8f9VbPRzBB7YdYO0cIjAwW0JHoT/RGaukAemHv
1ErliJkKSdiPy30k8bYkLNcMj3SA4nImCBDXDT8lU0bNelC3I1DC9Ruj0hjv1Rcx
r7lqGafOzsac5DZmuGyfzsG1dEP+clsSsIOdRa/j1gUlPXADXz6WRZi0dLfiywok
Pt7K1msFLSfpQ1s+Jkpfo17+3FMJgU0ZMrV94/OuB6K/tLJnjFAl7GSlqRU86XfI
MUjB/EFhdvLiVhvTT2GDzHR11j8KP7UJdwbWd/4Xz1/hPPGxXDWMDHIiLiiAWKjU
65j1BrB7Zx4DWZLs1rsoxKofMpPbM9wE+q3wDDE5qYAFRyNaDjT52rkR/8Z/tRSf
1ewxK09JLF6hDGPI5gkYCIuV1DHMNQkFRrrSFv7xJeEHGjqJC/izm0pWAoYuHXPm
JF80Xk023J4tNSBFm9diMkQgH2WZxyVEv3o9joeKRCoAsj7dufzsevVtYgNAsz2S
BuOp0HYbWJCnptSbWBK/jVjHvywJXYareyi8tWmAuHgWaZ1ePyPe5QpF57/+cZ7w
mIN7gVM5qP2Y7TbBPBSqX0523oWsbjtsdq2NPDYn0Dvbs53fjyWCRMppsR04lRv9
tBXBNeb7OMdjumFU0K6QtmLUBWGz9h8kAbGqQvSHbsQvad7PUPJLkBc+M3VN5l14
8alP29+Nwoskddvx4WosKg8ubDSllVL4K351r5VgSlMtiXeGtiVsXkzJfmHwLU7t
h1HRX8lTmc4haBe89ZHYo4UpwFiZUnlN5hJqpih+UxGJyoc8fA/4LBVpZEg1iPzk
11TCrspLC2tJkZnlpFpEvGrEL/9ZgPY1oljdfXSZHzTNmV2Thfd22vLNzGnnHjAX
k5qZGuRDEy/lcWEKtI+VbESPa2u9Q/yiKA0EFJRgWit+wFlBWL/iuAG2/n1d5w17
29tvA2uAJy8CtSFLMLPwjOX570+qGbjopeaeSshzHPDrExTxEGeB05kzAhOup32t
lA4UGpVMhs2dxRtp5ueto+loIKZuwpkgLy2PIo/eXy/EDn01b6JfvgUo/pW6aG7F
jRvgz5w0HxmDiAeOdkcNd6S+Zm5fTxXBSqjslhVy0sf7bmTIL61lwtaivyw7NNtK
cNy8ID7Jf5HkY+z5bbpQSVk4sd5/eyzcp+B6zT4M62URF1RA/CdXsghz4Bs6C2GV
DqgeHo77oJOXj1BMSYQ2UzCl19Ux3RjLt0B8znMd7pZEbI1iGVFR57jKtT5s26XD
TH9xIYRSrGE1idayCs9bk7EhfLF7ggz5n7KVMP4w5nmDxnoPOYZ/u2kpDQv2dHis
GiXkZumx+POAwjt1zwaociox19LGKO8a8lClXieJAdHUyk0nCJYfHOyIE8AUIhhz
OM/NmhhJhyGzmW0w4UPsxbK1PDfchW/QOyGd9pHhbGfMr47tq6bMg5rMirnqWj/l
OAV8sSfFpf2MWduydrlxMl7DIp9pZ5x4iU+Lx0gLQ6jLkKBDqNPqJiVFvJ6Qsd0S
Ae4t1GUIYw7M4lxZPuXighq+Qe8mvjhAaU44whdIDMX/9IB301xwyqUlnwhgIyaL
KtnQzbDMgPszFPFG24cSY6/4RH3+nINiSk56KEnfNdjaep+xJiXzn6dn5sCgJeWJ
voqzWLEGLGnOEm3tfminIquSLPYQ+LiW5uYhR/9/P4xcbQ1QqTNybcfgUnlLOkmo
ycsNk+bOXDUrGMZ6iqbZqNVl2mRfV5FRZnpjBrmwbatAvlTYIoCbz/rrST778oW9
oWe+idQpmuK7QbsNSJ87RU8EiJyOP2zvEz6oRQ17q7a0Lq9AMR1qKIFrnnAwEO96
WFFD8/Rp05YW9VPtmo4jLrtCAh9iEFoR4XKp1H7UJU6cNTOmus1W1tEUerXnMH8I
wmd9p6bTp4EY9N8vg2zuhOxWMzKyyxmGkFSQb0qh1UKY63mesnw3eC4dLQ+Ni7fE
zkF9dGH2d6kccXfS4AWVZi/jYCEjkh4BaejyZToY8BD7EWY9KdP2zpNheLSD8YQ5
+akkcwrBIxawfWqXukZZxfiaxfjbjGFTnWKRKS4u+WgCCsHM7KIbbRk/9KQmKzHt
naDX4Ob74pA4Xp3fzf38vMcObCu1nflYqircRjrjr1lTJ6pcvA4J1Fw3IeVJm4FA
G2FIkNMhvUz/gkmmeTLBJtyY3CY7Lx4YKxoPNZV1w3vRZPecDnfD8eK0l83SWlXQ
r06kAfceX01twmSPcXfC8WAEo3MrhlcSLammFHIgJSzBJfJ6zir42itjHJLCu+p7
Og+DIxPjCh/6/num1Of3xU4xD5ZZrsVQMoXJ7TqeoOO64RspF+1ThCpwLtWayvMs
A+78FBbkLjc9niSaXJ56XL5DwRECRhvnOaD06NsEukhgvMb3f8V6LwcpY3oyI5Vf
D8LNv58jdnrmE8aZEbMO+gyRC/JquMUl81ePpjLJeHVNumjI6dOQnNuDTRROlUTd
j1+N/SFL9muHuyds5t+0ox+P/K7Um/Ngjm4JJtY/JgjUj4mO770z+0FRDKUVF6hN
/wOtpdyeIzeh6F4zm+692wLKTsptCPW3AKdt8PrQHGHId69GAfuizc41Y19ceMit
sgVpGpf43ksTtRjbHtp3SHW5lcHyBbp4PFHmA5qvX9rOLN1v0qfhAjlZM89Jp8QA
iQHKjFuZq8IlKXUOpgZ7PT3jHRK5/1TsH47xPHu7Olxd0mc/r2IuXFmhx+h0R/4R
8Yk8aKePLTIykFaGymV/rCjxzzSBq/xyLjojl1rBcoaXy3cr9n6PEBtGAeEmwzCr
eooYoEu9d3tscKbWsbgkFwpP53DlVIttEmBurI0n9Sxe1EedBH6sHUQ7kYnbPwMT
c/3EGlOyfG8y65GfLe9VAymr81wmHp5ejJYvY7hNo6vvAmNW+SmFuc5Xe2BOUXEU
nsDJEbVORyfa5kHpWuy4SQSbnVkO8iYrUUOIXk4T9vcx7hB3+cVLFyBhp2gXiyD0
7VMZmfEvdKQtnJTqb7IXf6UmlD8jNVJjSI1Li9gJBnJUsmHB873R+DxjqJm0aL+N
/PSrKXuolkRBz+31Y7sWq2uUhTXZdSzI5728rxtVwuF25mcIXiLbDfbozyK9hW/f
/P+RXgWokZIUAia63bEmuRsIcjaz5tKamF+PXiD5mFWSRurMDAGFjcLme4jugKZn
hPeW7ZiLgWolf+NY1ONBoIIvFHER1wxIoJ7zCvqzpr+XuHKEDz8yO4RS2mJUm4yt
+jTB3eUlQuh6vgw0NpM5OlLH5HFuA0YWi8ijMIkiF6xufkN32tkxfmkBGhdwKx7y
9fTTXTuqWQkBqQZRTHUt5T1lXQzyvkUny6Jav7jRngEbtAMHoMOq1rJvZpXxmAig
4zZtGr+jXJ3yxuasj9IETANPHZPUb7ouK5jqDtJaY05YvfVsZ9Z+KCidWANLY49T
tw+YmtWAfrKtSNE+q6XECabI5ELtd6TJRT70Rh+9knZtnSBWieP++bHbewgARyBw
lctvXZAiuYxRmkyy3/LdBqHxivyeRYhgXlNl53MjoalKWzIwGY6/7ojam02tABms
B2mPHQY6imVG3vw5OPtTt5ONOjXdC1YL8JaTId7PZiXGrKDADxmhHsSfTDaBALWh
DHHIXgSsjJ5em+1ys3qaKDAi/h+ugkjE50buQcjvfEJZTCVNHD7SvGcOMJycJoB0
Mlf3/STJ3UQ2H2fRZ2Gs3iu5WCT5Xea4GUq6zNjBTAL+f/rk177hUE2cXieA0elQ
DkXNNTVWL/2u8c/T7tpDiEWBmYLd6s3OF5onOL9llKQKJCA2p2rJtZ5ZGX83Tlnt
svqx3mquLibAma201MZ3ecV5PKB+eeciwn9ycI8PCWAEmD+x3kqgZ2oL7jl77eXM
l2UZfM/CyqkR/KK2SWZz9xT+JQ7NxApcqcWu/2iPfrzPzZ4/pnaCigOckdVxXc6C
tT8zXBcW4UbsH7Tkh449hYNdxm8k1oAac09rgIIxkhEzS85LqcpEBczdw2g6gTNp
lzy0QmHCK/5EU5OODuBNpKZ4R6ZwUrUOGbNv43/Lp6Z/NZoZ8+i+v+HOQaF12cZ0
sLTLiWUiId6iXH2ZmBf1v7lgmD1EhVu8igLa/5ydSh/4gNAqZwFb43AWLl/JcdrP
Kx3n/P6BIbrOOGbsclPOmOk8Ze1FO3dhAqmILcGLumr9QUikMwBBak0Efrb1UNMh
g2+ZOJWn/hBBL2U450JrT+nripA3wn10Xyg25VfyutG6Gbw8ZgkC5/mFuHSvzkZQ
LmCTkbKT6lk5A7yARDHsluSt40MnDI5LiXAwYRD/GaVdzunWdW9xtrRwNuFe1ct0
k2WZ4Sn1CPXrFX8fT9ePPBtEtiVOICeq1HV0k8iq4GqJJgcX+WulBQ9iB2yllnyM
I1kL65rMt4SK0XPq0lX+ggfEhq+okIMpDsH/xjzKF1VK9vZOpM0lEM6w4dnvvDnc
FsB1Lod++j6m+2dwXzldPYerQPh2ZdDPwnnbZ3WLBZaWGhIfLdO7nfYDdo/jMJRA
NsCJyD6Uru3KZjvNB+JJ7Sutko5Fs8Yn+6K34PKdSqyY6/tyz1Ej9JB3ZHOhWvy/
/HoWOF6JYFhFWSsObdQCuHM+jk3Eac7qyiQsWTJ6rv5FnwinfrsvEr/vx7wy5M77
5JhDsl+10pHuQzLxIJavmnFR+DL5DiK+M+aaoZYvXCyVfoQh5r8Sz3Nqk2xFznD9
WT5OJPY1uXd6oCUCg/4kAx7MNNa8wuhJTurimzJg1bHrYg5kMPA6QpnJAtPK/Xhe
Z3SV/FESSa3OzCIhPwG7PQbQMHE3OjsqfxKyO0ZJ8ugbXKa3vJytB00mq/evIDVB
mVEFAM6C4Wq9RTz0PRjm+7XWatImPuuNNPGFd1gVZjXS0Qbyt8t1UyACBLETFgI8
L+9oUpcCnPbpmZGNHn5QDFG+Th+baFWwJN4hcS/QRb2zG0QOugbolB+sgVaFS8JS
V1NPRgopHyqqKd6G7PvxXU0m8sBECsnQqzBBJeFnJWmd2H3Rz73v7eykuLGhS4V5
I7M1rKZdoOtpwrQJGtGi22vGFJvSJ8JTwqN3VzrpaEtsWl/KXiYqLC9XaIEsoW8Z
eiXli871Wj8oXsrgxVSIGTDUrng/4cSeLRqkekXs33M54akQ2khN4VAzR4/iibhi
LVf48tLd/Wtz2u6t92ve6PnH2NZ5PAKbgZRrqTB7tDs1+bcCgW0t7aHvlbvbWEPP
ZrAE2hOolVlgZIiH3j+Ze1ET2GH5RnqjS/mbcgJw+nPp3BU07+cvAqDR7A8XoFZO
6agZus5hL/9k9iHIynwQzMeGwEk922SAynLRlSA4vw9gcLWrRShLCw61SqY+Kj6s
xFUEpmZDwyfTMChG18Cbo/5kLrpGUAF4weKCSwoaql+V2bRxy1kdW+4J+WDYyITm
uGpIYw9xCW8S0RxwH8zTqEZmMEZRrNN5BX0Ph5t2LIshdBQ203egzzaEqXPB5e1v
Y3KV2nWSDqzIpXNpi95x1UHcm7/wL2eM38Hw52Sk8Bgg3rZnKUK8rv6otoFz7IJM
IXg9JfAZSH61WnZL2xXIcGe5IdOyrDi+tip36JYO8OHfRzEahY8bnEzRXNK/O1t8
66qA1+7LpvIFkB/JHG5x/IG/F5pq/8+hXNz0GlMoesb6AeckF1cj0yk+rvuHP3vF
6jA0oRo/skqVVs5X1u0gNByJfQAhsyO5MzYYXLJOka3wH7VQH3a/0r6nEyhBCtL5
jSbaEPbwDN2ovhSBqkJlpX76XFHxXN03c6qE7PP1J0oYzcatDRXfPn9TkIa8tPpa
SG13uGVRDngFFsJ2iMh5LIp60niYzx/0+Ty/7oUSF6oJj88i302ye6v3F3mgcvko
km6LUbuP0Wzdnj/R7VOkrX0dx1nncq6k8dRRpbtDJJ3vl8MaklCBHt3zRLE6skEg
6vXgzhbSkVSTCEZuAVV42j+5u29igXzjLWBZaPzjCEwWH+q0+URvkLFD984K1kHC
H+z7dDE17YvRX1cMD85i38IfeuphiPILGtLsSSFFlqBF7fWAjQ74RMF+dFI+P+pY
AisNQvIgmowtsZd0IqcGhxdFHYSE6kAFyJ4n/Kunss5U2vTVMKWXv0FMWr8ZWlPA
NR0O3VXP0R4P4/L5nO7SB8SJawjzcqloF0z3qs9akjR2ezTCMr+TaM7Cvt3JCj2Y
l+OQN7hm1tLHmQg+xZuPJDB+13FRSFUe5vAwu2XNVUOnMyyagVA0wvH/5cctji5M
rAazLIDiuT+lkKnoN78skF0RTzG6MSz2Wnn7X9WwqhFdol70rEXrB0Pofv18x9Qj
0sdiHRF+70NyYLXLSyD9oWMxKh4abhwiUk1pWctLNvQGQF3pcbjA5XE2n0w8z9c/
5luP1MMMMvxl0R2+A4IFPTweimGVFuI2kW2YaOD6RkKJyzR5d1XeeEGbUJNW6BJJ
cvdlTjZ0gP2DKbgE0YdqCBIiDTKIUQ7Wbto+QaEu+zLIdGFlgGIXrqBAKLexvATb
GeS2tKJUYaIeRInN/finvqf2A9G4ykH5/sgPL6t03K4SmJC80dVOGUdcTvWABHOW
nGtwrUd8lJJqybpYD2h6CDgs5UhAudlfIHG1DHOYNITuDmja6ep7vHMLvilQCgnc
sjQkUngS9sOyCKORrXuxq0rAyMY81rGG8vwRS9e2loYr8cO4PObn0OcMmaAAfzzY
Wjgme2HIIEbRENfuv2iyO7VGD0/WpT0xoZkw01ZqlVUcf/bVSjc0MKONQQbkbgW+
F19OcB4gvjypBNggkoCjTbM160rdrGmUIeKBB1w8pPlwIG8DCMDs70HUf9uobEMD
TXXkRfXMDED98MvEyFpkocpKEy6S1JjZf3BhnHs8P5H/LHjIekPGctoKYPbpqfHT
6bsUrZKwRlsonkPmraoNMzUiRgjDRj+xa7sS/E9Klet0h4ClyDh+ZIHOsx8aDw4v
SHRoGeV5/9VZOMcezD/HPDDAW/m5ae71LPHn3A6tV7CVF0bnRgB011C/H5CXv0pF
yRpbyfaYlU/fRIOC2s3WqdAR79UwjcVp3LAIHnyFLUAO7UnZOY9S1K460V4rBJkj
ezaMmI+zR5R1pDcDFCsOFc2tBJXTZTRd61zR+S4TTfk22+hX17EQ8nNvFAlIKIIi
TcH8gsW+ieswn1tmqcad+CzvG/CNo6I1pda6cWVkfaFRWGwOtquy07rPDlBLnJt0
kHkaSLup61Zx81oqutNVsWI/AKx1AoHXAJ1pfYETr90/ZBSaOSxvjeDar35VP2pw
AhWlCRZFQYCQEUXRfaLNVYqIg8ouQa2dvxwd7hTmEv7WWJrmN196nN8k82FvAwRQ
K1t4dsyyZ5zeVRuLHBRbTebxzKQW37xWw5BSWnYfc4T8i1JX/uPDuM9ELqSKkMDg
B5DtJnHMNlrSnSjL/4EVM1vo1s8ftl4uxImZZl0IH6Es5WOHWZBLCr1W4f6DNK8R
M/NemWTn7mRroHcELZsKi9Ce10uUTXdYogW2OzIojWcu/6qrjJYmfzzyh1AHV4yk
1O28b2huKDIld46oDLW7hmbAHh7hYmpTECdruaKZwDKKXwAYByuwpHXS4cmWRifG
UVSWiGGf6Rn/jUHvR9+j+H+wAdXkR/ochGLqaj62EqvaoKfhzzv3v6SvgJrSC92S
0F04aeWpTRQ9GZX0Mdk94kVqFpUsCQ/yklC26t0omPx2U7VSeHBKiSsCTIbb/AWg
eKAy4KyRnIqL+3NXlMw/H/UOwWAzFF5DLUT289P3LMmYqsOoeKkK6KMFDp05B/2U
6DWHTk0rmB6y3cvQQ1VFkYj3TrC2Z86qWUqr7DQH2TJLNan/gOXNP0jbeGRDBpzg
ZmAm2F8Az4UDxkox+uG5LB6HoxoYXBURo6jWLD59cvSZtM0iCeIibQJhWpyuMnoN
wjKaLgrMfYom5SMDTju5j4xoyffTzTTKGAXUJvyi62hYkUkvRnq585s3qf0Tg519
FRRb0INgjBuZXW9y8EKfQzosUG8qYsFOLmInna/2ARGY/Hifb3NnT7GAwzfclc85
8SJztESosS41FttbVAqdRxM4PImfUHUyP3xFCIWXvCBdO59y3bizxVDYjZpGAuFk
MaDekVckIrPbBBWn5iOlH2YCpCT8i43f5Rv6w/1esVzQeUHr5M42ZH5K8b7cbKlQ
tQtlJ6pQjUo3Bv2LIvP3v096LkyKPhMWAyALyLPsNneL4Y1G1GfGkvBQptgaqJpj
YIsAKwtmnuz5cfyOEzsba0A84C3jSiBtXKmjSTKXqIET8wUDFqTSSUVZ8sNnJXBK
n7lnc4da5lyfZTDOIOQhYaMUPBW6Eg/Ekl6qsw1j08Mlp9JfED9+1wpnML+RZWMy
KhGn87+Lzhrk1x95L+0CC8AUgxQHuaFE7uLyu2R1dmYN5VC4+Y9dBT8AqzbovxnU
a/56pHy9fYJISp6tGdoZ/2NscpM0Esl/sxAFN7bal8heydSp0GMfKiJYY6yCDHSC
wIp+xPZTi/OUx+yjARnQz6q8vaYNm5Cw53VVSETYjMfJn95Xh/MdAy3NSTBCMNF7
P/fbFMhyuQ/kwz7o1LqyYfpYb+oKT2BtdtLQST/qd+IdagDpxwEHv2AJRO9scAnZ
pMlid5PssaX8XRn75udVIc3bEw5+jIEmsv2JkT4iIevqmf957q6tZYcjUQsoK0Lo
QVxqF/uw5yOwWCsaTHFmKqu6y5gwTrUiJDH4xr6PtT7vOCuWJMI7mUCbamhN1ULU
8C5k+7PcKNcwamy2P9WcT3aWjf5pykaA5TFP/IPNGPvN3zytDkzumbzRSUTt76XZ
SKxOXMJEIDL7W58LWXWsU6aRPgtm1YBqMm+eBf19ljjxkfAFQAjz4aI33Wsi8Ggw
XrznXbL4migUh7trCZMp0na+OsK6C2mgYWVEiATURyXKoph77qdOrrqjjdpJIgVj
qYupwwvsoM20xiijkQEZZhjjxTebudLTRUsPLMFfB+4uSxEBNcFjDtnxrLfXsvlL
Cah0W+/WaIMeQSkEFxpouNNMqBSKqPsQhc0nHxwO+wvlJ2EiifAFn7sXzXenLf/N
Q2wtzOUNE90RTLMICOeUU4/bmRmFy+wTQeCVvQtLb6f64qShKmpb3bmtfhZreuuy
CsQXeUm55mCscdP/KZV43VEKyJijsBAAHWuXAMkiowfBKUoDlF6VXRPlvTfjHHU9
jMuNgQ8nToLMPFmaTGPFR9IEoPw7sg2mWMqrcCV2Pba2Ys93pNa8ezS1jUAvNmtv
clxGoFWUSK43/rhWfC6ZJ2FXcsORVJJvZ2iInHzskkN6tO++r8vtjOH2dfs6jH0i
uR5whHhccyJRn1njB/NbJsjg3cObkkuhAaPDegVJUJvOnoBJHAcLsTlt1iwIYK1+
nEZQRjs/Z4hiOqZx7yfc8cEpUCVcG2/lhfBpCh0crMduF2gby3r5WpKITKKszGUz
tNyTvtWUd5PZn6d4YZxx3JHRAZtk6kfb/gZ19q76t8FRdpf9fM9MVQOtbkqippBy
Az98hUBQKU4Q5jgp7vr0eTAwti1NZ/FRLwdYEg/yGVl3z0INtmpmPcwyeleGpeq7
CyFdaiAd9KkLyqd0VqAjWptCO3IIwwE8sk91bGgDjdkZka0xAGXbrksIx9OdLLjN
9YABnHJs51xrbUgkOsACANBRJJAzwdJTxit/1h2NNnFxB9wAuFOdWw718VR3G8X5
JndZ6bUZchLAacaQMmjWTlIRtLGtL3FGBrBBzPHwdSyQITNuLeSDOZcQMvdCqjpk
U4HDErz/nD0z52ICKF+2NGkrlhSWvYDtrb4sD57kigqOc6EMIdqUCZ0rXX70pY5o
NGCHmfzAjlMNQ02zvH2MSSzPvg54HMSrbasS56XqzOUi6nbhQJVP5h0VQLMmk4jJ
Y9gA+SH3NF5Yk0LT7Plkab4khPvc9Hxd6YKG1zDUgggY8cdrVPzmnK4JHS20KMM0
L1snQ3cxHpWV4G754CTURnWRa99FgZcrpKgviaiPDov26X0ZBuVCSbMlAoqLb+45
KapK+ZTg3KTv8yD4nLUuOzI5lb4CLAb71tofJEJhsiCJrp9B2L+w4x23IufXkJPe
uz/ngOjbpDFDmxrSxbrLVk3V0miRLQkVnfksTRlHQHGLeR4BqhYxnanTY5k/NW/e
o4v7rWO85ynV4YFAeJR5sbFJILkG3URNndbzPnoQNiztNxJgIkSyp+8z/c3RXLKk
DzQlfMDHaQLBEWBE3txM21rgBvcMDjS7qxGrYoBjzynw9jsw2TWBq0k+yxL/dGdG
jhPPWbDe0MZrjwHHQJGIZoC0jQJ5nBi+lPITpd7sfrZNRpEGNGXj0k7M5cTnmtnQ
9BzmnTQe5dhSLMCxKEbL5iQvxmrGujgtm4PdxOStDwEIgPDcVcDXzzC2RcESF8rw
UEqqAyQhzrMl///joMkfC9LIhJ78UaWQa1dQ+OcpK/cKKaA5HGoskeUE6VrqT9n1
fPjxpV/oAkn7A2/N8oFBzMWwBbnIbxjPyU57aaXtP0zct7n0O8H+Ym3BF/fQ1j4I
JchrgqcKF2Zmitt7sHj//OJfFGG0EQkqGdP8YY+gymgTsYnju0p5ZLnS+QbWVtwt
WrI0UgFN5WZknlvVLpEfvZNBge/PCWzbU/W+uS3dX3vM4QpiEbyDwxe99bcD2AOM
u9huMfKjEMXHCetIJ1A3QkCbo9JY3hytZZSfLgaeg+VWAUNY5ERNV/G/9wcoXoft
AQJhm9KgtCRqcEuGbLjA3B5zT0DKo7KdHq3GSIJgwzveL+XqmUMzcRS8HFykwsvM
VmMczW/J5iIxRqCkvCTIhqP8tzDoJu5PAAfpYWHe4Jact3BNB+Kpzp9aOuvWwGWq
MZcvx9bxZqxUJ7yBCwj/L4lGkrdkOHPVNzhi/6PhEf8IIXEt6ip00EQWSULz1K7D
laCmcgsn/gUfMkmzFoImYBvrn2GmQFAe/EdDjIaZlJzAX4K4gIjFSDv3s0icCAMX
YYNcWhuGshd/FHGaAM/6qxAs/kA9i9e9yXuOmAryMScUY4ru9YFfuDeLDQtEQXtd
zd+eCFkEYWnlOx1uiGp7v9VeJx7DWzoiAT8veCC0nk1uJ7TXGNcyfm5ZlZEpvxyF
jMEpzDBzl+4VN2iYEvooFx1QuwwO0BUI8ZxVlmG0+udkGLzyD8ZiDMYKN8GXlcfb
g74E6GZf94euVaTJQljW+K1Kye+GUPDqrm4KbY9iZonqB94QbIDb1jv+93hibw8o
855Sq4nsJ7OIJy7rFbW8TypL7TCwg9eeiCA90VtMWdY0OwE7m3kcgBPcvvJ97IpA
oLlQz8qjbLJdkLZPPOt3w/hqIWy2q9+lRZ02Tu35ZFyWnY6Yslaib3yUSN3oyj7F
msSCOEpi8D7scBGfLvfNlhN2NZCbuWZGBc2pUAtsHX7IAWmqMuAmJc4W+2qtjndM
2xvlNFkkbS0E5OOGFSGX8oQQZ2W/HH74c9FJhSnjNaiZCL1yIj1sAs5Jb/qhNRId
s2YrRWNjNE3N2wW+AvIeaNHsdBRrdU3hxqxdc06uVPYFJePAAehodLovFneuuDcP
tbDt329Uj5hmBF2Ct2n/p6kI0JmDh6OWEaPn6CTlUF9AmoFRAF0ButQ4j7u3+z83
JitpkaZhxb8rGqbz2dodifS9zWNiLFxr1bAKcSmeuV9TlEOHKqIhq5i3FpDMo2n4
bW9QLjPFpXDXHkZ4SbBk4s7SBR2wC2JS/LhbjX8SOYXmFezk7L37bAr1gPA312d4
h2QjbtqeDwtLhq+dMcy4Jneh/S1pIKjlmvZDLuaoiHLwalL2mpoy9j0Jcfa0aaCN
WmYWMGGT6gOyq76GQ+NUMEuJcf9ltDpm2tz1QsWhQzYZAthuc76NzxXNXIG/jJlk
b1SSQosf0uQqoS6UwNjtyYv0Q8ORAvRTTwdNnMOfhBI/ffLs9CpgEBrtaaoqDsfb
AWbRfI8OWSkfN/gFPsxG3UPYtyHGQSIxyqSY4SMFsw/eFGz/mBzTqYRDWcuyjNhJ
uPkHdFhNTQe3v9iLnQoZAaZO/pDim7SEKCkilJ4mDsWDNjypUPh2F3ubFraM+Vh/
vF0FR326NPJ/gTZVGLoVJv7NVgTi963fdfUgCvRZCxGdXv5Ye6N/o+kjKprFb4PP
VqacF3D1O8QF//14/GQlBar+M2PU1fEi0hlUaK/5oXLjuIHCBHsiNfbZS7Qc0h7W
P5dpHIGYSGCG58ckTkLa7XXy8EsWR/MDqz3yM6P0ImLGvUNi7QL/wMs8NPvMxjRA
iLI1Rn5mI0DjINgKAtvjMtQyz+aBnVhq0V2hbrXmWd9z6Br01XZN7BLBmtKALmLu
t7oNMDAOuJHRRP0xzycMoqRzqoJ47bTYK2jF7w/bvFpQQR2SiyS0j7kxwxGQSBz1
0MdkmXeygJ6yFB3qC/Esy7gF1WnNFz0B7y1rb5pwUrly02FAhghXFRaY/VVbLTVo
cTkVDN2wSTz4fhYZsUGRqNqha2TW5CzfOb0jOUMCEgb9PmwtV3CKZmWK0SfYjxzG
mLuA9Fi16WR43FuLjUDBK9sl5WUSD3j2xq+V4muEUp8yG8brRk5jVYJ2avLWcKGo
FZgYxGUyLYIMR8SesuOFOkUlnWYCzb7fj1JCAAzfO8vD/JwTyWg4QSmyy8TQfq7y
b3m2samRhDLZwMSwRnoF3ppkfTWgi5Y85p4xUDo4BVqHSLAttTgLushRiuRtdgmP
mXPfF8uH13Qu/adiflTpH35oWOyk1c6avx6mk8EDTS7bLnr8F7WIqDrFAhH51Edy
ZieIkilXz3plXE4OPwtPf0d+DCIoNj2GRFD7pozDnK8NNOo4/tw3e5rS8rBzbxcc
65tGZeba1e82ADmjZncLMmi/T83lnyZXYv8F40FacBFGtlTCdQsFfCJg2hPMxSm8
PZbp4KADZMirrX8lBB2mdeZQbQADN5eXa4GHkN4pQBQOZ5Lu0LtVLSNaF+aEEoao
GhV7/YcrzgYojL/mXNvC1riOUOWdVXn7ipK9RIAkFGsoCa1ZHbwXpizDnEZlUNGb
RZydRGWp9CZyVth/F4n4x+JsieMAiSRdAsegGPV9BqV89j0k+gmirXGoSy1Rwp2O
seN0Xg6vsGGyJEOsQWOW726Ps4tQyB4PpqVgsGuXd+TwOmtpNATQCEqCi+1AjLQj
soZHPq/naIumRDTNHevaxlQ+745hnmsiFEkU55MoaUGiL0KgfTwCK3wnnNSWR2AB
bv4XKhafpjx2lZQREDliOnZhsfBZWICyyLcVtUV/wYSEzZ9eSmcKyWN3MvuGSJgi
Sx6JJUQ2lr2dlwV72vSq79QYwB1UqM5g+5Bl2aUlUUxyJGz85Uv005inCIjXlbRI
DtsvuP1xL/yOMpGwfKiq7TIyeIVJAfKFh7gRcY7yp7/AxiuIdJtjmMD5JFVqo4rZ
O2SZ74s9dUMe9b/Oa3xrxkrNm0ewxy/7RSVKGC1BbMeWfAdeQwKvJ7KwLiDhXEC8
AbE2HC+aRZG0Tc+VsOG+tXV0IA+mAsJ+u3S1+S+3cdmoKAcHt65INj9YKzfFLJgR
4j7LeUREkoG/tdZxdvafDubjjoDzm8qDA0Jtf2FHSQp4/NYJDN+SYKVJHKc5xgcp
dcYjGHSCvJaz24ynxFlFQqMA2uh80bxA5Xg8sX9jzFNAAtadHggne5FaDPugamnT
pkH699QLwE9EcZBN2YCLr8lYI3yphod5K5ePrqeLwH043OyALUjPOagddyl6PHeZ
1p3dxHDhmc2GQoP1m0LNqKAfSt8cQtARinKaytHV24y7zcLbfr8pGa1BUEG4JF/+
QyWNm39F/7qNq2zsu8bt8m8Jm6XWzpxZnn3XzBcCZwdpTyVbrrgOcZrnc8/SpwZO
b45KbTS8IUw9LqenwDeMEklKqgomhfA/RHA6zL7/c6X4vjuTffaPXe4rv8kswQui
Of4n2qKxYULEaHPMw9YoCJ/UaXJGMUmJWv3TldgD26Kkz6zc6nTb5qMLe84Z6UTO
ZTa6BWceSJrrgMSRPA2NvSNqoOkJ57mXAKCmbEnbHfJvC7p/6vH83GpXXme7BHBS
2V6twGRf0/CwEXpibnzN6KaZLWetgVtfmA/2U16mxjfTovNa+fPtDXWGDZoEEn5I
qHLKqstOInnu3WwilrrRfYlP91InBjqmWidpgOyfWtshErWI+99DmoC8QByR6S3m
FEpz8lqI9eaaLjgG//bAwLEUITV9J+ValFmFBs1w6NqVj02PX6tqWi7apbnqbSbe
cM4SDpKfM9yVeHJYYc4t6UiYl1ccqH/SMLw4gYEmTHkUAfbePCratmX7xG9qvQof
BQbW8oczk9GM9mdJF+fKJF7hFFtLqLKFiwoMkeMhysUVGjbmnUVy10YX+VkWN7c+
rcZZhDkhYMHqLoM3MO3UKzQ98KAMV2T04d3pqi6y4eNCXiBZwLm1Cb6hFgv/usDj
zkYzVb7jP+Fzqv8GY+FIlawW1o5lqnd0MTUj0ftlPGJ/WZ4EW3WiiHwexP7Tpv/a
xZZfaOqfjHaT+SoxDMRYmdUd9q3fFPiUQTyxKoSF4JGHnKUAM6/hDaBpTce4t5Ox
ll3G2mec/3BFrQHUQ7Zq0pcTMPULRWF5C68Qf1yCnHO0X+xYtP0aJ8DXj35xeDvl
3u0T6LXbUZGEBP2cu6QaTZ3YKeGcrb4rxJINtFMI39FMwzWlGsmWGb3HCetaybvc
low8GfTe0xzZBdEhxpjKm7ggNF4UKqoxTeq+KkqW7m/W9VFjupxyQDcXoiJqsRpJ
1I5v+qE81joix2EW2kRuiL0haSqxrmxx3cOai5GFENXD/MbvKUWHXKXTeR55zHSO
d+ehdPqhLg67EW66n2Z32/KBlpW0uieiHc6pljdzwVb5zNYo9r51g5I5blHq0Vns
YAIzZ5TkV+PBJf/yM+j0KAFXbtvZzXdSU8vJVLfz4WCWarHs/yZhx/5a9bQH5/oX
yzxR6Rmq9FTw5inFGjsk1U3+yehdskGSYTtMXXcPr+zh32MKRvXyS6sp6k2xWEIm
sfQ2ynH8D3xqy64Bc4wB9sXfpcGR3LKKF5+HdK1YBRGZ7JB+WLkqdsIl11QrxAVf
11STw+14nSIuubwzwpuQpO+3QqNt08oE1hYaKG89vP8brs44AaWRJX81DIYRWNgc
zPRoUSjjN8j1XtXjX3cQ3U0vt7RSplk4iHisJF8HIAXBI2qtWx9cu/zzFEFwKaYJ
0YA5Xr3xHH7PSnvqxb0cpfiyhYcAgqynsGZTQooXvFHp3oIob5p7nCaWPn3Vf6Ax
bVCUUL31eVLmdXHgYpo4l50kdqlbuJOjCHwyBr+kJxUC6wuFzfRuJpX4eShAzE6b
Fug51QdDnUzFksOy2ZkAqsR6ssdlDi1GMksfLYD/b0e23/mY7gDP6rRSkc/9xfNa
j5yTyQBiR3wmV+gs+OXr+N5jcz+aSegdc9dfvztregRXb/yEFJ3xSCtnlUXoYaFG
gsKRdkEZL9I6Mvk50krOuZDshujELfAIjYy29jG7MapWE6TrzJ8K67Lv31/XzwWo
DE+Ugp/tMc5luscCkhTZDxmT8hnFhlwwBug8RW807n24lExtjqogJCfZdVuQozdC
st6CJHXFUxKI+kE9JY8El8bn6bix1dzM4ktpz+ihB91DLTro4JGp+CZhnXupxgnY
8aHdm19FtHFnzuSQe3b0RZHuvysSVcs0JzQsFvNM3VDGiOamSfLXdTAtgQ8khb3w
DkFOCXMh/4alT/1Yv5R0qdzyGJRH2IIsKU245RySS/gZALcU1cWM19+QwniDI3FC
bk9GGRz7T0NqgacemNG6i7gNVWafskVhByUSi8+AhnsPuFZ1ZfDFSxC7B+nNCSjy
uJmoTr/BkYCxdcMUeievx1fkVlLUHAHLgEjMKLhwWO0JfioOKK5T0MbcC5km3gK6
qyCBz6rjHU5Owv5P3o7I8yiCxWJaRzOjAnGajfx//b2iF6/i1yt0HUpKSEgX5xSL
OlhJdneKVtbg0GmZsMDbGGMDbVya6qNd5F0Zx4xqjqTRb/T1Jjlj+0aVIS2joIyL
YCoVo6F/6umCLzQr6G9qbFJJAfKOg823cX2+SYUeRITRe6AtBx4JymilwdHvsq7X
obnYRt9SCNGhX0YyNxGs0l9HUogQC2s9ftMlI7v2Wq+ZjWbZyaqbRSSt4KUpDkfL
dXQngJA+xUEP7g+bWoZWOEB/oCtpAeLv9n6r2AIpas0oc6DRbvcMO++WvFjW71+M
uGRdToe3witafoP4E8Ubb4JI0rp3+xtJsEih/80nfZ4UJ/06jFZ28ifZJETSm5N+
ZpOgFMGCVIcHP6Y/Z8+gvzI+GmvIXzH4HsQzuifaGEXGODb/lR+oCo9/Heistyel
O/LLtr4np3BsV8SO/RLHDb/+qwvKbGppiFP67wbGUQLHouWyx+eI6x1WxlRY54qC
8wG/PSdJBAy7upd5R6+4t6Qhcdwei9fG1LLKOr3dXqYh5W62Ub0O1Mw0qlbm64tb
fuT6gRR3Gco5PBK2DmZURnk3HbOvUshKTHTnBkJFi6pGe6Zym0IVnl12kKjDZb5V
r4P+Tsh4UuJTEFjxLp9nl8QmJr9O8gBVpJpvRbNrPNnBu8VUqyyCIQLtbrYh1Q/7
0leiULfg3nJhK7LTLcPwqGjYJTzGeJeJr3x1H8VsCjX9XVh37jbmAed3N8RnfqJS
7fk3zflfze+M2oJAC/sLgCX9BtUup7v5Bbp0Uuka2NwLqijmd4SiNEVaU32uCAm5
IxoztGv0ZL9Jqsymywxf9ZVol6qtXMeLl1ypYenPFloYc2MM5y+LMvpUjD32wiyZ
/XGFcfMOXg8eKLJ100DbRxEpH1esJ+d0qVvho4hVm5VHtlcQU5VsbtDKyl262Lev
ssFpeqyk9/yy5ClGAV4t1f9j0uyZq3wNsgIVFoTLsxa9FAHkLwQIZVfZnqa8OsSs
BFPK1Q8Uwnj17bVbTPPY8wZScjjhzQAOpqTKd+auya9QwNwtLS6oMz0qxWgc4kqA
HuU8k6AMhWl1qljbJXO4G1kju8zm6zG5SvxL6QuvkIZ9q3NlcuxavsnH2uTBI8/B
WoMDAwLFZgnMLPrxQxOghVqFx0Nj+Wl2Xx5H8q5Sqr2o1iX32/n42m9B7vdL2PLa
ltpBxT7shbQR+POt//gVvXgeMJM320zQ2d/+jL7Q9sC1AG5N+mcja65kcWamaugH
ni+kJqtWjHUTB7WUKMB3+tCAtikRGdj7io6Stz2UIt5LmwvM9ZYONJaXEfAHIFt0
mgOyXaMb1315h/EaxPDROWruexa62aJpBpOxg0QOtzpiSLNP21YnGmOuan4FFQgi
EwTmoxXuAGA/Ipwf7dEQ1W9zAAeetE04XZWgDBIVyCM2ASGiP261yA1fCeZ8xda2
ltVgHknGhW1bAlemV2dmzMXi9tu7ugIVoVCmvZt82yNYmUCD28GItY0HA/pNukDr
GJMEfYtysm1nZXNbkdsNa9DZ1qiGctQHr0jzjUfxu3gOolZErGV/FQqcCzoCwPAQ
pj3zA2QdE3tSPEfpFL8ojOGu6+XJMZ/lNB/hs653B1V5kU3GWe7JsptgoTZP2kBq
wTOd9oHFi3O/EG4ruo9MEKeZGZx+cexBrmFaWKCMxHhZ1OkBcB40CtBOAHz8ndsy
53UCWG/wUNFbXzzE/kQh6c7+6V/W9Ul7fs4Gi7iLS3MyOpl1asr9PO5sGw4k8AUB
Q8vN9muwPuoaySRv+QO3Z7ilGZIehuxwDzQpcmL+eawazvycDvZ8tros0nTL1Gqn
VxDy94kXFGQp36FFVnK1AOx1Bi39NvRLjD3eQsBK0kjK3nKCzhL1ir+Mcpt14ZQg
rDv4g6Bpp5pJlkqvVWHZmgLm4iAOqY9GQ8cnd516PJ0+grTleY3PL+n0WAklmcrA
g8ubhOxixR1Q+XovZgT/G5QtrMAAksO9w47PR0EKwt0VQ1O8QSisVn0/fDKdV6Ot
aCg8Mr3eyHWQwF52tNaq4BAYyV4sy7+Axywxaz4kwtwAf9Tm2vxqp+zXBOpt+0mc
yPs8AfFjsMP+XqldzubBSdMKD7IriYMvJCA4AplmpvchlSB2r1gP757qQkGjLwoV
cTTt2bb8+WYnk9DGfzZg/hmATKE9UsLfICb66vqqQEBZr0g3dFm7U+tYcMVu3Fr4
mjvXqECyPc+EeB7/wYBHWFA1HFtbxtLrUX2bqJqFqUZdPQX45roLmH05RXGZbydP
qPVy3wqXZPYEiRWPEWQRrIGowAo2pPA2fjkmw1x12FnojB85+l53jR/mBe+ITcGm
DREEi5dGktw4rxS4EojaLw8LY3ouEwsNlWyl9Zk7bRszgw8juBEUvhPVtYUrOogn
gXVYkTpvDebNedUbk5rHM/3FNlY2cFv/jDp4i+9VzoCWLivnNuU5ih00tVrfWG+p
SQt0L4VA3sKxK/CTN/yv8OkcQ1nOjdYWAHZSHpCxnfH5vHKcXOrwHfqiYAm+0fW/
im8a3r9KA9EYdBGTt0FulFyHYXZXU7gq1x7A1uSLWc51C8yqSK3peesD7MXcbtpg
tI9oALF7heL1Pbl6jd0p+rUHk7hDvt7hE5u/7itjDSmu+xYSSMsGhowSLHCt8TA+
Z0RQsKSkhb9LivGTs43dU4KlZwGKgRISBTV7VnXG4kfTqIle+yGpvDE1zEd/hUAL
PeofenvWON+YhMz+TpVG8hLEEDT+yXuOx7yWOdnmkqvz6fX8qsVTqvHKOEiSMTpS
P9ZpgIE/4XvhLySOI5ulRKMCjo4RJwX4fkEfOyy0VI50fl0O4Ru5aVf4IFyq4pZm
yRQ4s8Dr+LfQtwbdioyoVY9QHSl5pRCompdprzccmLwzHWiGei/ky+IVEIgcjeNu
Bl8B0pA5fIH58RHqUKCQmOBBtJaib/NCNfJNxxZHZSBYxoWw8V5ZI/0aRageBEHZ
uW1kKRKuJyBc+SdUrI8zInO+M2Pf0mMVG89guLfVC62lvyqUqRTKWnnrjIhU3nlF
CpvqqHISVaNKmtIlrjYST6x7w/MdF0u0FrSCes9QYVOjYAMaR3aBJq0Uo+ldW6Y+
9g1fQmuVUtikwFhIoFE9SuLK8QkOKR3o5g3KA4Wa24fn+zhtBdI3k4ZMXR5Z8Wt2
KAF51OHXK0lnLnfIorrqSFgUNYXE8d8S6NqzK6EGP2RT1wb8VIA5HD0yWC3N6rZf
roSaymy6QGk/ZBPlTdhZsFyq084dkGTxclVGVbIb8JcGed73IQfyB8F6CUCyTIiX
iDQo/f66Q/543mhX3QKREZwQRtQ4jekPviBBvIZ22XTbeh16sWkdoK2Zd9WwCaEj
JPwcR0fbONBanKzhJXUTCJJdVShSy0fmIsNszg+czXeuAagRpHrEzhSM60cKqfBC
HYvtnlF0q62eiSeP+UlQZbWD21xFU2UBJnseAzdsNMr0a2gn3Jaafvgh//LErtjt
zhs9VmnDZG/XdLDKFrOSt2DdRwmn4I4mveC2ut0Ppgv3Rg6xKL7euWDMbWq6mv2Q
8qU9xBhqhLI+hi/l10QvvPKkcTav5zGp2EZ1eYO6FMweFjYN4K2POFHWxyP3yODL
RADUQpVwbD1sUuLHUxxsNINXFiX9Rg25rVmO9hHDI+oDVq5NCHl50446EYVP+cg4
An/u/9a4NVY8pfILGgh8oJB4zkhzTEUQ+WH5fczzh1qAdB2wNa2Hx5XJiwElSdYV
Av3mpZjwYlTvjin09FS680pZFIGjNlsFK6uyxfnDCwTN2GVK4mJ0ePJcAz9NcdhF
0Gx/jfTQYwcbghXapQwxR+4S8xK82nNW08dVpvrMUnF2DbW+IgwBNIOzGU1pol3r
0YlK1vj+YOnkqP5A49AdBzRE4FYI3mXbjkhUYveTXMRY8xVZlLmdIzmVj5oqdmJH
i+kQbdOAx7DEaK1ibzjUxmcNNGZa+ZCcT25Znng6SCPoi/s2Lpsz+CP54tECxUee
8PpkQv3jP5H6gMzXjRlVDimaDP1hrY6ABKNtJ0hXRL+Y25/B0hiX9IIM3WpVMHpd
fkgF2qn6Wxb6rx+BlKDcN3MlvNGiM/v1xoBYxYS5E4tmwLlatwnz1/m8oqgBTdFO
LNtv5dsqumA1iwYSfINKF4K1onjZegqICiMnpzf8CU6O0EUOFTWZEPlMlin/lGKl
U6nIQl7m0oPuaGnR0PUjBOMaOKRoIlNI2GfH3De7sFi7PZREElMcROWyn90J4diZ
D7xptVCma6HOEYvnwC2Q/hWcRjWKEjVHVIJArukyaty3Ef9l+I64onHmPlVqBDe6
T6RklCl8TyAWB9INSaPdWdrf4uahTajAtvoIHGXgsHWKGz/17CxQ0IypciuAwKJ3
Z/hrlGf4Do6B6Z1dlfeahSMNKRh96xUlKb7aYeO66TE+oCEfk6XQXRDgDU9LnB7G
5O+o4MjlQCUSW6KqbUvj0kec5tJmgc76DD3dBWhv0WxVA8DzgWiOAnbt8cxBMQck
oWAV6cCBEG+6SG4QwltW4dN4CpTH+kADvpi7cfPzrJwKrlutpja7ynh5a9lkJUf2
s5z+Bp+elh7OHwx7h7a0HSTUxhMSty34svJbjMBvaeoaWo7PSZyguBVjHkCYcLGF
BjCowDujl+gVe7u3tFPE16HHhHFw38lC4Ll9XtrQWtbyfhYcbv3Vj7ZOJpmnBpPX
wfOux5BNwwqSqOxJ4iLY9YKT8hY0XKC97aUZxyzoH/zv2OXNwZhrGdDVXRFODLf7
1Qz8g1nGOFWNpZVsoF4aMMVn2Grb/bsB70wecBpmE5rcquC+hRdw/rj5isDWYWp0
q7IeqX452Qh7FwXggv+U1AHSJgaVAq8RRk+9tsJWmNNWB6gFbzeiOm0bEgCt9TyA
XI7k2D4FCeAuajqDc47P8/17PNm1Jg9d1TlOjZUdbre9qSjqafFYpRrjAcGqkwGB
YFlrT0n3jHxXG3DxKtloGn5z9HZwrRS7BaIAypzdl1eQxYvdfBw6DSkRTcQRPLDZ
xTTrNqwOv4hTb+LRvV86yx6DHPv6xH3UThGNn5wMqqeJOikBzJZsJXRB5A8HdJIT
/24GmIFWlBrgIZsoYWYdrS4vGn86qHSyeJil2xGE+ak5iFK7OFU5LxKEuDkAGQoJ
4CPc9y3nQedEPqfQMu/fPavYdtmDI3QsT54KGFulbV7XRX+0u6cewrI5o3GJhv8y
3VADIlur+wygXxrnCkB75C9sXE2GxjVVcIM9gVPgKEt54mGSE5zOrFLN+vLJStMH
C9GZkM8zbDsVLNIgwyukMdUj6xz1k0cUaciHaKCMLN6egM2lfvqMTWDB9/HYUL7J
3kvY+Qv1Peujt3VqoPISX48iKEFYpBCEL/6HByxMfzdHh94Ba0BGVj+DNmaIPhIj
DDwrlfYJbIppDtF5vrxvSkTOM2FT2RiO9F3zg6Kc+VNn/1IPojAFNRg/0n7T4jo0
bzgRVZzhb2bpjvV+GzW3yUTjXYXDyaaucOsc4bUYvHRM/Zx10lRL/B4l7DV/LXtP
LDEV2WxSmG+wcqq3OveV6pORXRVz4WSAarf32jJncpVFS3V33xkE3VxEPwlMIq0T
jjp9wFo5sF0WPKzVsr9PJpJJzsiyVlEwG9Y4a/xj6BevqtPHZY9GK4dBkMfZ7C1r
VqmDDRPbJc8R+Ok6X6PZ84o0flslV15In/FYCcFjF+nBmEtNUJxTbvsB2jkXsnkn
9chrYjMr0ghnmqtprIzfJaMV0GfWYibsb0MM/NTN+JzRj2mBmJiAsPTcvNWBCSkq
R3gjSi3oeNnjccyy/4zOhkrPp1f2WVfM4ZGNgI0vMLaH12RTrOXK3rGPvszpN31o
44uuHaQ+IVOhL3Qlfpbiyzx7a2ydP/fFpZjkgJDP13Jw0zipKp8KfFj3sDVjcU7k
NhXSaVZX6CQbGTsqcne0o6NiZ9ePVUtqKp1Hf8J5J8Ez4IBcC059UjYFgO1nP8Qw
7fA7LmTO2qcfufQqXfRb2n+U9oT7Y1jRiFTpNoitEQa6Ze3EmGKiPRBiMFRns6+F
Ocpr8ehOyNhak9sQI9Wgti1FLcuUf2dJYm73mQz4nCVbP+wHLkvRFryD4mwkGLbD
CTISfcf0T781zQbAg/tnNWWnxvJ2/jhsh79AhvXthe3jnK+XwjgqDnsgywud/nj3
u2pWZfCBpP1xo4ssopsBFpDB2xbWTmSvL43BalS0DMXEtfja+2g0pqc3jvtpso1q
ml0x8MYQzr0bmQPOkOJk7Sq7DEhXLLSUULdXDqbTI0VpeK8flfoDYdCQImIYPfDq
bXFvmGqqqcRGjxg4YB7OUY7bv7C3ad2lyFlDN699rPfH6oA/ZxPzccUCvBu6D6eA
ax6dtM9ZWkGhGXVR4TZJyiFe/kMIpDOrs++1/uWqSn7W0WOywzhfAsCIoMsBVlxu
BQlb7iv6Oc6F2Yy6qq7MXebm8sX8fPzJNVfxvePQAR7LUD5Tp8cz7EF8SVJMjrab
u1LVfXiTYaMZT3EiPUCEksyUfSVZKUC+wKs16assTqHFd0oevMiMLL1urhk5n1iN
egMUTwrunoC0txxeRKN6w5HeN7LGDMapm/47MQBf2x8CGIkL55d8YPe4anOv5vhs
OvxwlkAEuCMAlUvhQIQKQgISMwH3doBqYdTmoCV5yiRqMU6hEuT6/otFZ8AE34xS
uqTdqs9WQrkFXK/OMihj9k6MnK1sugL8y0GbUNwpLrMTzBRGrnWpNDifRr3Docyj
+zoa0IYPRPc02w3fwyCMDDr71yPSfRnUoidtRpjhSGROcqKTh4noAwMgFrfOY8yr
OpwkAe/4l27w3nGC/gmXKALSinnioYx5h1VXmVhAPh+K6aoptGjLhB9Rpk5FZIny
G9Az0uG/iujfZ2AvdHFgJDduQZGmkPFnUb/MXxAbBWhhacE6uccTDrapvWueGTqx
rJM6/Q+p9kq8tCJU+wYshVaCUIVlTVivckdWsK2+36nxuBh+8fEA24Cai2jfcMgq
OTvOZf443VN+qzC7JXsJ0gEtkEauQI1XzF3+/RT8AyocLl2L7jL+fd0GJqvNjqNz
PL/CN7U2iGzeMVcOf86X4jXn6026xkwK/0xnPYAaxCMopq7oaAmm3BdrJ/thnxKZ
Roa1feBELaJJ3u5Xqk7+Dbq2FEuKNZnhFG84rICOfTC4SslIpaNWJSJkjzs4DusA
rjaAialH/6UuEzfsgVTsS4NZ5n3Da5VCIsfGTYisx3FPm17DmCC7RnI+i5Y4gJnW
PPksOhJDfqmkArJeoQAOFVPiNporVwOfNhgRITCkIg7C/x9WJaTOBphEdRDc6gXK
eBMxxuVcwqNYOKen5WyFm1n0jg4hTGdbl3OdQPSL9dmqfX9QJNQpeCJ6MJIb3sZ2
9YdcTgj5cjc5bUWWOirF+lwmgNo3XUqrCZ2/gjLTAOZZ050qqXPxlb/EqYI2vx4s
o65BnTPy8NHED9FUhTMO94UG0jC1n/V6osE8zstgGkzJcym4pM3xirIZXdt0uyof
+MAWDHZ5rSjFBLPisIK4gZmDfeFHu9Mici+Z+Zbybv6IeYiQD7SIotO+nRRpko3L
DVrbMVEXLkt8Y0vASsS9PWXpAYngm/PfT+hW8KQFoiGAqnxcYD7oiGlItTLJm3DY
zlXNQlhQbsSkYuHk+nWpQuo6ktYZQepQWtjmVGbu3V5MfPuNJ52ouRR9hUR3htK6
NeYvfsQk7V46ZZDw8KQrokpHcIRp0Z8YHdg91XkWpYpRHDbes/F+42WxxRw0zLX6
IWAQAVbnCX5S7r8Esoo4JpfisG7OkiufIiHytoak1JOgCXoLDSDn2S5MIASVuc/W
MEJ+j9CvfpzYXS/XRQaUhF5P7UG+URFLu0zHzEPE9hPwJpUqfAN5Dlb0mD4m+iCi
eG8zbarALg1VrepmRz0UuexxF8Xo9kc1kWg9way9J2qmzI7VlC9OpOzUrH7clj7f
5t5bRc6YfmxHk1oOimIsXkMUVKJbsQvZE76HdNpYtWzM3nUH8vnL07V4/0nzG7Mw
j8jxzdneVkK4jdH0VSv3Hyjnx9/FzQX6t/KRzxGSKjCvBq0Y0jAGT7ewdcOyqdVp
iAAklW53KhzWIjYoxsi8D0wgErsBsJmy7DE1rVPxDvo2hxPSxmSCI5mIyAlJ5U/L
y5zivxvGMzA+kn09BIYjeBwPOPSmEVO7XYHk5vhFLnEZuij+qMNQMBjSTz0dy/cY
vO0zRWwJrHl0OUKc+AI8n8dgBOmzeIG1A/yHsT3x/sj3kLurYHmh+91/T823pSj4
phMnPXHn6U+xHNuZVybo5x7nDkOHXdZOW4HTD5b65/zSGZ4Jt1COZk3x4UpBD+9p
Y2WZPiGcAaZKn6HNdq3/jzMqjmdLfLkMAwAD9EEExxxdl3PlKL7H+EvtV/3jiYuX
aj7srVqf7R+i2ePLOVLNnIhRnfHQbA7REj19yaCDcLjba+tn+dQiXLMpIiLWrlUh
vZ6Kln4vpmncY10LE8HPowhR+7sO4NTu8egSd2kl5FmHmH1zWa3Ppk4PhD2dNgQZ
v93Mx2RrKw/oMkU4F7zK+RVxyAtZf8uWeOzSLOrgJl3DAZTIlOVImbagFInFZcUt
EFerSJT+qfU0wHXHzU1o3dLEQXeVqJq4tMZDdgUecceBXYpw4w0ygtNSBO8SZz1S
lFS71dCawnwKz1E8Ien3tIx0UWX8sqZ8upyyO3g7jts3+KD+RyBT3NXdNkN5Fa7L
QgftfYWMamwp1QvtkhtoQLmWPS8b1r+/jk5b9IzuU0qiaTfFFbDXrTAm1npNtggT
uwj3YDItoOkIkMoXbfOmSz2M90KJ8iDOPGJ8fZa6LQg9eA9WFVvr6E0Yju0xJFO5
AFl02+Nq45pVG2LpKTi/h6joQK/8GrnL6HUGftQxo9D2/jJPqRKV7lj670eOObJt
hGoEqRY2Y2C9uqcj9qe3Q85yUanlfHBHH4ZhqLGAswAQSISHbtY1MqvplNALdwcm
kh5aVpsHJDyGX9sIyeoopUSufttqAVK/mqS09o+8nMwXYW2nq/R4jLpdSKyRIfnM
SLPUOaiPzTMnWFeXLc4Hr/73tQHK5znRIiwEN9oqNLNXf1rPKasIK5vFwHNWrZif
YHQmB2yzDXEBBcuFQwAYP2myGCFRlnO3GwPXSscejgh25FFKUP0SsCXnnNOCM+Ob
N7qbf80qQMuoQXnlDUTfNSuvTrvptWAmQZSw0cumziKjNmb2WcI42nKr2U32leMU
z1pl4vG2QiQ/Um0nF6obp5FmCSl+PLk3NGCs4nSWb7yarzBP4TuTlUIQ0sBJbnxR
dSYf1mPRklt3X4UEWim+MR97WEEIqAT0Lu0fVZbww1NgJFo2nXnoffST7KkNS5Cl
HUTevkVTkgK0pv9B4LyKeQRUy7KqcuE8HaNffT6JmYO0/1tGMQrl4Ci4zcMYQa/H
hFbujG+WVIGPGb11FMV0r6L3x8V6kj52jJoLVTZNXcpWSFzUFwucASTXX2vnHCw0
buMmlHAWzW3bFWzyWf/9woRQ44VhogxKi9aweNxe3YViN7Ga848an0lhzd868gVC
iA56hjIqvTyWm705mM4A3yYockGzIqXzOyEkfP2nvMOYdWftO/GBHj8ASn9IyAeD
MWFkPieDtmVktl01WPQpyV/03K3oSon0GZ6XMWH0y6LYQHLtghtn84L5IkTADbC9
K/NP/ygPNSMr5CseCrxCSluRrlS6y4RTR7QY3CDBOCNX1m5m3yf3yvpRvSxt8SHh
4X4XndPuZpMmgvXZOvjUJVwe0ySDJyQaUEikepYb6bqfh+xeA2g854damPZXcqC9
q8ta1tpAp1eONO3KikiRcSKCKXie2ZOuGOhjQMwUsm30wEEH8hcKI0HS8g8hOUVR
DRkp0kBlAmTgFkpLSKdwQpz3+9m30nPQH2GJUL801jiqiKtlY42TBClOAXOtWdkV
qLrNkSJbCm/5Q6Evxce+4Y1EQ/9gsbwpB1k9A1fHXWiJERtiW9bXlmfurA4dF05C
TOXvOxxg6DCcNtWVMHn4bT7zgxBPnvBk1VqPKoZ1IqnAuadp5upj/IET/+3zMeUL
khbym6+SVCHRM/Mh5GA+N2tMhBbsbGyv+l3odkf9F2xpYSCY5etKUkCIrrlsKXJF
4HmIz+oZ+H/KAuDLHg3eOzv2WcQ80nFzZbEE6rv6Ufe8BSo5gI1SM9FqkyN5ouhH
uVGd8qxIZl2Rfry2KNaDhjCuMJBekgKLr/UABznAWh+SXqbOLhBnOD9u2gOGFwQW
/VkBRAfEfO2O1zyBSnfCLNUo6E/Fdr2JlvPCJ+h76cSE+VHxHr+7IkD6J02PGvvV
3Sce8MJkXCCdQwYeibbkPnMSgK0CBdlzf5YUgr38RzpiXlMPiJ9qf2Fls6wz75KT
llKpGFmyV0FA3TvkaEzAHcQd6scuyXhMPKKoZ7NSm0doZmqF2aO45zXe5tX/XCvT
2GN3gXANVXhhViFTPqLOtpLVMWPX0sXS5oJNnAJ+xvStFJn1ruChDgn56Yq1fYtf
l3GmV7+sSXC7EGgA1gbfPMwizUOgswF+QXbm9AvU9/ABTbPHbHleK47UbTSwEiAz
00gZO7GzhTcS7NGL8kheOgtNai59YVVhrwLo9ynr6JpC458Mx6/fvN3I+8IthB2I
w+Q3UY9onyPN86hW0F/nsCPaD8HygS6LtnuAxKte0p1TlqZGn2xsVYNf8e4qGgB2
j21EInV5jAY6y5+pKWB/gWBAM58mH1zZ6+85/IikGBEh+14KlsBxPncUvHM0NfSf
vC9fqhiwMMPbvsRjJApk3B/KcRLkO2TLNZLozwCWTI85jNg3R98mNpJqPXaOAmJx
Gcwp75wTJlJr0PLkZWlfwoVaoC4KZqWcsEkHLurdm/i5caTkhr2DC8ssShnf94TN
uO5mwW+pb13aseka3ERZiDq3NaYJ560FcsU6aHkPADtQAzoWhTDQJd1HgAJr5XwQ
XD7RSF1lVaGoCzo0wK+xqR/5anGLn8PSSB0qe+i7+SoyoxemYw2fD75Pf21FXFqK
/1w5kbtOacSjNrwiMrBpfpI5j8oi///qZaGcsk5L1ztfsNe2AnDfSkF1l5I4L0Lt
vdP0bwpp+UQQx6JbWSKhYB8GVh6EkR/WyzoIoEQqwej/Qz3jLu0ODiZ2ALyF0tQm
6p85lKSXLD5qk2i0RK4GnIyyUnmVSUX7FRB7zDTYR41pYV3MKBPhwKlIqMKTHsz3
dMOQC7DWCAOtuf981o8KNAQTdj8TOaz8spqNF1B07kDTHUsMFCCe5ax4eHnPw7/B
F0liUT57tioNnCXec3QlGihJ5I98TFGIJVRLAx5zkcjOATtP4kQms68+//jBwkoR
bNuPtODZUOfIUcsrF7zP3f2WVdSfLiiFs+M+J59nVh/T6s8gZrlrjXa7HYcofkWq
ODWjRT+SxBfcp+sRjxY894vgohsEapT2E180d9KtJ7YXbASBO/XoguVd4ATGeagk
mf7TqHg2FOzCQzexGm5Tr/HcUQOkAsZqgXSagwpl3kfjYlkKGMwESBuN7xkraNq2
xkyik5yhSLH3vyu3NMrXk6oEwYbZMzyEcGXPbklwRazEphDeYpP7mSReo/7uOdSE
m2ZqPhjqGGesHVS8AnBvQPG5nCQhX4zHP35OANJkhFvTxcIEbruhVNJEdx6m7p11
+2qvkZ3KqQ4xlPhSgs5l0HegsOlXf7CLZAbgkklVM9bqurX/QefUPpqyT1FDfSvX
PEVFT1Oy9ZAsWbPSxDNBbDLWGM0z5dR/OONesKhzoW2URZDqVn+dthIMmRoYfBKa
9b8Fg0Y3fmIvToV5Gi+UAXH2P1j2N83/kLd7zHG1VsFbE1nXD1XXRpnZ4z4kmNtj
rAB4L4YeZQN55Y5OhmuXSfXXIi76JoYqvKy+HCsNtDjJAV4zLSL+4LgI5J4sV7VU
G5Zrnx0X0SZ1oS00awoF2ZZ5mHpr7nju25dO2RAs+jcdZmDsED+PR2Oy7BdP844B
Pi6+rV5J6ruBTjtUtVugTcDfc5tU8AxGViEHbSNAOZ25uJlkUEiI6f2w0GAB0fXw
w1prVfr4sSNrw8LHLkEGC3SMGwFKTC8S/4q1kg/CiJG0moGP4ctg4226t2xpUHNK
W58qom8XTR0tmzUEhGELZ64v9/n7FUf5keKfpf4f01IBkFf2C/8/pVV73IQ9u/6P
bY3I0eWtoO8Z8lXb43QZbOqdBBrgEO7UKzeWt25vs6OS92UobUbPs8lW8kxayrWe
uAMtORQH9Q5DkZsbcnnyM5iinBdSMz2xRxYT1Q3tqjJMDH5ETC7GBKHjRR4Z4dhy
n8koJVUtJ76jjx7e/pANeW/1ZWLcAlL9Ppzp2PETkqvLQvki1V97PKaLANwrgv8K
8cbBfKkleeHWMKET4FlyiJwVEliVkRf+MQ8vPrSta4IqqfD61uWzTt8ipLqkYAkT
AGx8WXEyNvyrfFIJ6cKMCv+M0w1EXDLgw+rqdhzC5N6FNW6dII+ErYKeKAnt/qwr
IV+IH7NvlBWRd4JSTOEtEEYZvDAYp05pskvPALctYLKvG/LPpzsw65n4vl9d+rLo
irFNULchStj0gfiP2yH/OGf5X/AxDZtMFLAtHak3HYHXzAFztKNWkGA7VAJcy25K
3GrKOEZ1H1JCOZEwutqC90/dgMJHV3zWkH5LMd2hF4FOtuEJRfLD+C6n+T9H0Xfa
1lTsF2ZCGJUlz9uGjG2HPjYR2ZW1rSVq7eG2xpZXTEgYT1Y3DeaL7Z1T1pezYK5V
Bv2h4ztnGOEhVXQxL3iJOgBIwt2B5jCG8ydm2A/kXRk20Qw9xkom8PIO/09eG99l
kIGzFYI5Wtw77FimrUCi1WlooEYA9/Rc5QVb9x1KrGYWeUvT200w9kNhqCXqwi54
LVI24EtIsapFHu9Qtf5+mBrzSJQhU8Q6U/2VNHUjb/G8W9BwK44WKonaWC9slTi0
mtG9RCaWdWyOy7/TZ1UvuyhKZnCz4Wd7e3N3spvmjgiNXylvG3o3IZkZCHyjhZHA
ipTpQHS9F5DYTMoJxja0HYlu6Rb/s2jIuRkKf0qUgH9iZbJq0Gv6tr9s2xaMitE0
18rGKqt3+wOs5/NxPoirYbTjPCeyZGQsafiv9CQB/4qE86TSXc1cbcMRGsSMVhRO
QV/W2OBfZMOXv+RCLXsVELV++f+BrDEuTSxX/Y221KkcnS8SuJ/ABwTt42tivSTx
osfNSEbJdOSWucFLMokWp8qQTaDVOBAs054CY225r7tjJdeBsYbANq6Z0wDFnLm/
kUzzDiU6skoS22tdKGpE9+q+FYzyTzAZvAG8yt3SJIy12h2hgV3gW/Ng8Xdg6vdR
4w0Ua7tPWaSedM+m8VxKPV2kBt5Vhw8nq+xXrqVT/psL9AgTrLNjk0EHxEL0Dk2P
HNNywlQdOH1xNs41marwWob0S4iTHJK8HY5hXiLb64ktwNTrXD+GgXasHogggIoY
RI5+X5E4sJjyuklDYF5VTEyvw0aWoBQw8VXWFMXkXwGrSUFXUMgbKSfVArTXSGJH
IbsICCM/aVR8xUvyh8XGhNIJX5FTdqpceTN5vLyLVz+dftDbfvnmvUU2t1bA6AK/
g1CDkEUCERyEXuj3sWYpZonOwvwo8MlH2TKxknPjm+0S2fHcG8WTt0BuNtpNYjkg
7ieNx2peVxHsTh8uF9DkU58i7bx7SDbgK29By/fGi41KGxEYlFUSQ73BfTIb1VOR
tZav7CzqjHKDwPyk/CpsI+2zlH1M6GUPPWeOrTY+jXR8/KzTedv4H6xYtMZYvPfI
eDOZVsZRwsK0HoSES4vH8m6UNYuLraBF0Nf9oT6gbtp6RNtvBw0bfA/maMdvbQWe
iBIMHpbDoUQ8NSpWsEwDg8pQ0DPOFRRoy1KP5++oLTw3sfkFOXrfuGOydiKUHjfU
EGTduaG83UunQkmV7LCkCvjlm/0iAJxpavPoJvJ9LJl0P5GSqiGUdGkbpsj+GWi6
oqZ9QTe3k1EpTMZEAmsyIuc48lpUjZAIyg7mL2k13qAXUpBt9dOxap5Bs5pmuw+D
Ip6OKyuclYknklSqQFwRBBoVfYzATm57hU0EjIc6ia0nyZcYIKsgGLV5/seh43Rj
5yGZVKlshFBceG+gSq1DzK+vuo24VHldRECB4d6G3HvJuY2Zqbp2hdlU1E+TCBwi
UhNFMJGaJnDWPVShJ9Bsch4bed6oQXFESuyutJ+6OxOd+y+87uKFmUYlLsbGjEkS
zAxLcORtvmrjrisV/E/oY7pnyLzYt7h7PAjUAShzn5qB5E0B/d3dgzw1xzo/zFRS
NRCiVbzHG56FZZqHTQ2ix5mYuulexlS8ZI75kR7bLqV15INcbJXkjKYZorLwfp5C
ggYtSg98R90wmkEJbmTTxb6DbgcNGPZgwUNvx31KLiQCaUAbgTvRQMkpTmAslSIf
1ykRwZqVZ0gCO2TN1XfBoaef1axrhZQ6tH5GRyTPQTOwyZEL/UrWt5j9qrH/RFtA
0iuR+D2ZmK9gcXk6oSwTvaUP5v9r2Zbev59pRzllI7UZrEi+DQ8QIFTFeZGIZfBO
Dj9hjahiVSEPLiIZa2jkdlk3Q4aMbkv/rHvDi8GPu4Fatw+aXyEQneDlBwh8w3Vr
kg1aaiGElwPXm/+W8apo78b6txAtG+yi4pUEPWD8oZcViVpMkagsa2zYeYX+AAT+
DnVUZTVVSoAxgDv8saKDesK9Fvs8elZrmQrA6BnW/pTa0tXCkM6e8DRfauxmHlc+
sZLHiezXK4Piom/HnQrOwG/RuB61EwGXuYP8UBMLipnHhzKjzJrAFCs41kyWmrfF
ipbgfhWlJQHOz6IZs81ES5q/JTQPIO9RihDwi6R3RuU6WN5Oei5L7bfsI09XqRkG
mLOjLDLKdehubIPLS4DSlpQAIBtWQmrbS/u7rD0n71sXxrRHcvsxKUSO5fccYGvw
D8eu8XUJCkMMp/4BjvdRRUUa2sXxyPUlaf6j+eHnxLsYHbhwBxjE86K8XDqDf4vx
gGQ/YE1FLFR0gmZWWx5D1W1Zqxzs2huhQin9lcfL9mbZZeEw63/DvnvFAJ00EWvi
yw4gttB1kRMI2W6fnci9f566USnQcbQ1g6rB7iIMWl9e1RIBTEAwAmUhA3XZCnWG
TndKUg1llJs7/ks81bgL8evstPu5pod/YuNd6na0PSo3OSXBQ5fZgq2Wam1iliTw
qkVvdQR4tmi3e2TJKoDeOGqivnmsckRvmMPh31lCG2YdsERcuytmHio2R3vf3RhG
LwwCu3DJywf0UyjZGS/4kMhFKQZlMOs0emklhZZ7ShlpzrY0qa3kb9nNOP9urMNX
u1JyqtLRe64wCuFq8fZSFD2VyoN8bkl7eJggX9IB/ZF38WY5EGwrFP/kEwr5Ta9T
l7qQF/Ldh4pVx2MxX+9KoFikt88bBbOjLC7YE3OKbq8iSf2NkhjqlFAZBAX1gPxi
7AYJUUahfr3van1MltGsXykwpMehVjjzxDLqWY0Cdg4evEMPLQL8ZeN2aBTil5R7
Q+LO8WZ5RaYGZxbUtIsOXhLcPMwzQPi0p637fD8tvkTbEa6GszVia6CqW5peKgze
gJeFDFkcBZ58cmB9x0EdRIXNkYswBMf6lMLamzxoaOGDwtdQaaGPkM72A8ZC1m92
ZKTz+o45cAzD7YlwjZ5W8nFQf+Qs124QfVvpufySOwnh79v+bKsW5+PrWjcGvX8t
izb3oZVwubh7/Bdo/ilwkMrm4Yz9ubL22xdxneTFCcHJvhln85F/25OVJwQm3MO2
0XNAvHVbVjgCZ+7VshkZfLrtiJQNgIeznRBNF6LZ5YJG9J1tYA342QYA9+MsoQER
RhqQGSWv7B8hRdL0LoSCpNkkhUMAs+8r/yzUKsQ0PYwQYipE+sgpCJ3qzBJoP39j
RqL4tVQ10RtOPMMjIAYjqz4zwczLqSDi4aejuYry4qJEQyDosePXGWVwMX64lsiO
jsq27qiuiorPosG3aaMDSC0/JQr/tCUE6sjP2dUC0XfkbdIn81rUDeE8zMVac9hD
LIFUp/HhsT09UyULCiHaWj/0hg5jvpnk9orwNeWo18g1KGbKuk8G6U0VnhMmj5lZ
Q8RIWB/35hHYKs/QNDU6JGavUGy+2xLQ8CmrrXPAgauTMoWxsjz1f8+102ykoiO7
IHPCowJXM3151Z0w26XOq8Qx9lr9y3GeQQ8BgF9x1wahnvPCwtL+qOVGAm4wp2iA
YpARnIM4w/sJ+s6ErL5mu2nEnvSh/ofet+tc+/dkNM5byOskRKg04164W+f4whHE
IxOvvPo4n/eiAg/4cfWGQDp9XwfcNGIdeMPobZDJZ61yZd6z7VCljugez8iNFfNU
Xm8YbXFBaoYUTMhlKQ4WdYh98W/QJIx1ckvnK7RWZMbQT2Aw3BTqdng9w8Hid/R+
+7OtrvsCOAfQlMh+6HoygSkP498vf/Be7P3aYE7+NpegIguuqjnGjWuaHC7+uqGc
0QSE8dWNwIXcJt72gnkLoQUKd7lH68K6/OY1dWIIANbUCC4SxiHgZ5nUnb5SxK0t
gi7OYk4Oe336sbhOWyKQ9P/ZfDRZ/n8uoJmSFpWuUHFq4GpZsfGlIS3YeGEy7sqP
OjYtx7UMwjm4SJbZerrAc5E6zaWSm+whOuAZ+AeyV3N/gEjDp8OXDeagKEpTpRbp
cpG2QijZZyKgv/Bh9IBz3J4kGoiF36JaITLz+3z9BGFAy4Swb5mYzBV9tWV96q25
X+H1EHJVZMQ9D6ptXzSX/ZdTBN8htBaYjeReiuOeWIWs2qn4b4njSYoRorcgG518
XXxE75iLaoWx41mAEcN3obpNUyYou0LWOkhrHVq4CanbuQJ4H9di8tGy1wvZALOv
B4PoZH8j/+FrFzd1QF5mf+/5CJmaiAJAmN+Zr+hf7uQLuhCEejqXVUoqUc+gMtQZ
D2AfZ+gPo9TFv8MOPeBDP2mgy5rEan2lBlIrXN+VJJNVUjv1SQe4ifbDZ34nrjMV
4OwGQkYBdZo9NCJPZ83yEdbhKnGd4rIi9ig5Aeb3Yng/Y/Qzbkv9V30FA0v9DFZt
c1trbEljACu5Gx9UFuhZcfVE09jqUvVIAXqmzhFmShZE3VKWEvw1c2QdcDqZnvAi
Vq1ZBlOK+zjgQKcitaJ/FQ/XGETUHfzfkqymNlWEDrq9sn5KUg9Q743BBkbs37WC
bRaCiRh68SbqH9phrfZitnquCkpag+BBAKTee5RzEcr0HGaVjq9yMR5YMSzj37He
anHKjIRPLV/wf/NmjyvMajqpXNDBi9qCfqEVnOQfslWt9D3hpPS/wcg99rBTR6kw
WRkqiBnAOvbnd69qfgusKkLcVJTVgA29BvOyVzboOHc+AQsG3v4tlLXxP8IQIVkY
d2L8nF7Bm4fr0yQlEnfghCn7ZzL+8mq2ZcPH0mWilQJETfdUulL3YbmH5jvu6SRx
gHXwLKKM0vDGDbdIlt8cscjgC+v1AeQIX9rXPMwfwUQ6g9q6SG6UiUFDQE2QUCuD
+9jk9BkUpXdxWOszDEOut3O1mcIkoaC/wjj5GQ7LeZEjnyRAIGcIK39Ro3FrrQWf
TtKvLuwM/iCoJv7RyTQJm+F9Bm0qoDeObg9UYdXGPedH+edf4QAP/weYn3a7muMN
SZQR4IeFUYcT+35TGEVSHa+S2nPNTkJ+3MjyjXR9Yl/SvHySc2Rac3FsDoftWfTa
OyD5wsQBm+tFk4NHb7PgpdYR++6L/gaFmgcaUdAQUoz4YG04oI/B7txl7g6DPIOG
/XyNMojUMGvRvUxl5UURiGg+im0ZQ1qIbJ7WhR9P7GyaoFt0vyqmUk3QMpII2yY1
1YcpCTlBQzkbISlskoqBhkFKhqWaC/BDRCM5D3cPsIT52HMT/ogAuaa9XEchMu2d
Sm/UrwlUbFfbnr8qBQ69o/4EgrSYcTTpJGdpVxtpM/fj1UW306BK12CjKrQ3j+6L
1SfPQAVCacS5sa2jto0eglqOxpeyGsg9VGCCRueb6iL5VySZnxqd05RhhendajW3
1KhM5BrjyznFghlEoviKS9pbmU35LaUBLz9RN547X1ODZT6Vtvu2Yp2YRcrNJ6Ks
wIoKkOKWZpw9MMITMG1Y90/2BT2PYP7F51YNZqDuONHeXwedJbOVBoPFebcrwlt7
k9p7aQPDJfpJc0HaEcN3VK2zRXMhH9w3JpqGMmj9bxa+EFl/nHh2fNO5qi6woqGf
TO1jhsrj22k9C2EggrY4ap3e7U5nH8H2STNFzAhENo94C/WMa6xVQiZW/YrR2bjT
G8oIoh69Jxoaym4+zqVtw4/nZd+uHTkeoyaDV0GT3VM3yM3OAbhfEIOGB4VLS3g8
+jiU77SCrfSv33EC4dmuLrLvedGk+Bzy/JvpzGKyHs3Lr3VZRInk7LauyvmzeEiN
VG71q5+PWDyUk+6wu/TJ60txQB6oTRBi7KShwu6rPDZcCwVsB/XQqF0ZLUNQHjSv
1Jo3l0K6MFPY6vrk5FFzYuNLpQJkUG8CCtyo9+Cx8PM7wCWHzDUiPMPkHJBWNriN
lxsndwLQpqPBuhaHeGdGqnNUBKvdy2HFTLDMcDRtNfFqxoO8bkb2s2S6EAgYRSEj
vIGcu93ak7arM7U4tThTd3QGB/L8+Sgh33+K1c4YKtOWXDSh9yCu9f2uSgloj8OA
scjVsaWYoUfew0he4gOfAqGKzKGGZptXBc7X/6/t1DHorXUxwZzB5u/FGtvK0MDn
1DrcuA6qwqMo8m+L+CCNeIB1rHtDx+qdadIu5oi+pJC+NTgWHB8PKxAtakyYHN9G
rZIA6iCDhbd0lcIftshrrS0jyWKgxPkCthZ4A1YfD63j+b+aUcuSwxLjwD2d5sOY
E59elKzsEEEjtBNqqBM+REvbOs8aW0F1ETorJ2KfozID4Uit8hhpslHyICxM3F9w
qGk0m3Wu/b4sA5ADn45/uBNw6t5LUHmnTlsky4J/nMBlSu0mzATAsR5pM9HwywuR
iHt6sEYGIHzORE5jnVzIagAF4k+uhDE9nDKySJbulBDUm7kDGYsKU5bVHnyKH4JV
oVtEXJJ+ZtIgqR4LB9TJ+cz0+9ps93Q9wupCvaACefBqSk+ovm/Epn7OdqIIg9Re
xQ+bfueCAfNscnsW6KaKCR8Ua+HdIELPagSEszIOcCBSiQp04Bj9FFpmyuDCdYoH
hmR0/RuF1vH5GY5LNyXvHqU0mAjjc3fMoVLRGFbpRmbQV43GxsLs9ALpV8POY+Yk
JW7/5Wky2wUty4ZxhmtC1iXdaoV+cNPhqMA1sfd3f01GB0hTzEcduys9HIS8ZVGe
3+rYRV8es9McBSROQ9qSfU9QRNjlKbuxl4N9gHZKRSZRDDkQWFXxMCbI67E9gvsj
aJ4TaR/ZoxGdQDuzt15lA6dGSVOak16CUAM/Z2eetcly4kD3dPiuEuoxUGp9tVQX
iY1gyzBsC02dN4s89l8sNidXRpN4G0W/GLvv7cRRatd8cdLJiYhs/7G435KuhWJs
KWsdzG1rUeurhA9f7D/SH1ScbITO4dT4SAwlaucCgDJ71wAZFgj7dKLhDs5RscpX
77AHzgzJjxhy5B7Rvr+hlv7PeYpMyTdlp3sg2RUh2U5hjPybAk/WWMJ/mcNXJnPg
T1Wnf7FNLB6VCUkDblpilAQWLBpb2fbp8L/szISNMs16gjtqtlGZ8xWn8sZG6t40
i+8WNt/5mBx7UMp5cDCm8C7LjNMVdrTpPafpn8uhCK5k0H5foO5OCtJQ8aYpLljS
cakgoB/xS4nSfydnPQsemlHfiz3LZywzbjizkGTZyf0cJXO8blSQ0eDnMqfH97rH
zZFC/KW8c4tUVF+B4zxADB+2Q3SOUh9Vl5zOn49JPh41ZRjJU6YR1c2iftRBQCXN
SLLJolVmZJ8b71zl5nWj/Q3+gyDemTwjNAImLGmS+btWNGpWanQin1m3Vy5m1NbH
sg2r4FL29uNrXqxzJI8XOu/pcGXev7upgE0+xVrXjGy/YIisTdaMzP2Z5P40MMQg
HLU6kl8Esbjm0aKF8j66tUP30jbKwKg9gKV3NwGmRwr+qsdG2HgIvaJZ2A+zKhD3
Sf3YQ5VzLntU4fog043aXh3rUpuddClrU4/4pM9HFYVGhqjxYcVqZroYvtI1OSud
Sa2UGy6CC1EyRTnahwG5lfUTsU5Qziq0aLK4H0WQYq7Wej25vhITZjkkXYLp7ehz
UTOYK7dCWZ815QBOry5EZ9rQ0MxdeSsY16giH1FMkTErcP35wNJURny9f8z6vuzk
BTDJfcRQj3jKPg4tXbCMHXerlEk/M5V1e4zPzsV+UJPm0oIhDFYJWC+tzsP7RlxY
Q7UfVv0eXzFwal/yMrV74TYjBN9ZMZRfhHokIN95qxwMJAAxyI2VcoJt72U21Xos
dFYTiVOgdkmDYr7anFIXgOqUSff9LPRjxkgZepVOSB+0oppPOFNRFWJQQxeljHdy
izhqi5mG2liywpJ76vJuNv0834AQhjx72nHKfzqUU3FjKPvMtomGBnDw9hdSmdyd
XOD6A/kbKXv177KSPz8WmosyeY+tkSUXNLcw1HT5NCg9cotxT3wUg/Y73L40ek71
JJVKGsjYWEkv/hKYgNBf9yuVC11VODRyLr6jfVUnD1rcmjqEFO+6xFPsl6mpZoJZ
ZZ2dhHj76aogU2J+C3mM4Y64C41kyx0n3KBuELxzOn6Px3EyWVtSgI5+WYOW+whZ
9599m7wtS7G7Ooi3aXlus3tFYkxTBNm6ncmtE/EQ3+B+ZH6zriVJXH93JfbAo0t8
ZnBmI0/GjBPkpMj0FNgaUIwNY4CUz8kq/8pjeZqJW/J10sHaTvJPkKT7tYs5h9ES
MqnkA7/xoZsRUa2wuKpwV3soBdVSu2KbnMKr78qEFCxAE7GNDVMMVMpUkVTtpyog
j8lnk30dHOwykJ4379enPWHvKCC+GO3k4jGxdRpq8+r+B7sbVaI/h1ccxN9b2GQN
lTwhul/EbMgLlO5x4eI5qBe+P9Zjo568SQYXT/wWQURNTieXb2ZHLp3UWxFkyvNV
fxFna3Z8EFQfsSJoy5GU73vJZ2s5CxaNNrDnAI0XFi/OlJc75CfwB7BsxtfJadCI
dlHStOfG+6aUAHKFaT3x3/E/oJJoEyFawu/pAVX3JOZaMYcm2AQLEa+Wlz2HRMZr
Q5fSsC8SKBwMQ/zGOzwRSwJgqXBHMuY9V3BbanqmIrXhmgQVP1MbzP4XEz9kBAOc
5lNZyVnGC4WtTiHQ+9I+U0Nvbf8EM799QnARXGEEOB6ZaEf1/4bGRRZCZPbODnhF
0w+ECmO/Vyl9MDVLNkZZrV3qAs3K1SSgBKwBjHosXCFAFbOJsyH3aFAXPpBitN3J
MLOjaggBACor4fNmJk7GkPQW1aibWBJZfERR796ZuRr05IcjC2o56vbbP6zDFvlz
ZHrc6/YL3nXjJsH+rL+S8YnTSx3rwVJxOj4jcVvmExCZWpMgdA34uzfdsXspXD3/
4WajBTDo/2kiv8D+/OBJmf72O3ix0q0F14Vv9CHhYbXiiOjDuFV/KgJZC+sxSf5p
hOck0BDYHRZUeJqzFxWDTtmt4PZkoYMuHvQTXlW6qtTeHNC9fQGo0dc/guCEroLi
9ADkrqb+zhEQui8afLBRJagCrhpxeonYlWL7S8kMDdnHbk9xeWeZ/qHaN1wuyBit
/2FPhUxKNB5QLUbBnHRKOoCyI7CfoIv/XWoOaKYELOQboNAt9tq5LHPEItAtL2tU
GeVL943dpDDDF1AHTCU3r5woNmaqpP3XQ+fuzVz+6nQpx3wxzA4qIfEJP3ogbc6U
Sr+ux2h+SFvOUtXtAomjU0vqGwZvAR/4hpU4/yZ58BM3rPIGTdNSa1jTGIv2uEEg
6hMK6AS+gB0b35EVLORCfBV93s0xsAm7RQsPNtkbX4bVqTJwGdbUFcB7Lw1f0ewR
yRJO7VtuQqPkY0oIdde65WPMwMY2EI5lBZMDkyXMeOKibDZmfYkIU0mIYneGf4Kg
qFokMlKC3hSsBky1B3DCtUdui1niG6QMDDIEHpvHG7J19+bn630W4rDBcaffpGu6
FAxbZpv9KzlXf0g79JTr47yMacdD0772Mpsx5/TdQ+6up2kxFr3wUmtDxL3mzzM9
xMbchCSZL+Vl3j+QFrZL8AhPy6e/l2yfvfQZhAkIbHd5V+nnPuQatJTaye2LCJLv
BFBwo6uZmCXLmFVYxdGX5TEKVVkN2+KbSgytFqIk46SUjpd6tr3MELyDQuuPzhwi
qJkm3vB9Ri6huKx3v9g/G1UZpUezVW8Ft1sO3KkGObs6qKRMtXUpHIijehkpgny/
ebUuN0An9CYJzM71VmgC3+xYRl7UH4XlGyt52l8wRfrfz3si2Y6xJMR+5AUvq3nJ
kOxsnMTjDovjL0VZj4cid/YyMz4Z7xDGrDnZW6cHTX77tFiVXuiScttQFGRbIj5p
DHkcR3pzA1MaTVpUKFPI6z+lUgtTPfUcemkh2etLD31eU1wkok9m4b875og6G3KA
qpajOapVudqZMdgHebHtqvzh2T+zZMUqN5OuvoLxJ7NUskTDULO9e8cLg0rvSG0m
4MZ7W5VIkNg9iQt+R5Ks8u3LsPN5kpZ/eqFita72ORhDGHj037OhOF5MhfleYTKT
4nWcbC/mGnQRnqHAqWnw4UpSbDwPYDiTMN3NhqaWw6lukJXu5i6q6+6WttRFUXSo
LDmho/vhfl0P+JrzjgrpueMhJVWEO5ek/ltXhFqon3o1eMDQ8FxVdPRxLIIareVQ
eYTMGjq36WCpgAqtEiHh3MyVFysd7Dz95VxaWHudeA8KdYEKkb/pJqjHD/ZdC21z
m2uyOXh9vpjGGff33to4XPpzUMyNU3L/MRyMw4ITVystCqlfU/KezwUi3r8aXRtP
mWSCs2vKhRtVkeSMlNqAtHGST85GeLg/u9vrflQTEH66sfU4My0CzuEu26TcyaB4
sgYTVZWZdv6X3J6NAoBAFyfXsRXwqCYycGZerJqvrxqC6M+YH/ELT/NWhGJB71nJ
E7V/MkfSW997FXTQ0AMBGLI6PHFsJrL7C6LzMN2TqZFGPJ+Htthd2JC/1HIQU+1d
cox5KUu+cKsAHQ9bvjfTLDDrZNKvdv2aTT5tW6IeoLTKJO6UKWywIN1N6D8dE5nS
5dKOw2Haoa3q1PU0GJfzAak/KkwJk11d49S576SM1fwLIdNo3bAkHAJHH5EmGbZv
8GFnJnBVxGLhEWl9i1Sx5wp2lwLY0e/18HD6hw1AnPsW0n6KJed37sPDTBlUYSPI
0GapkSRFle0HmflWY4O2ZItw5EcCkkTMBozfjJzaLWZ4QQKt3CabS7kUmprfht2d
Ts8au/FL/kkbjrhvHuRRC+KfrNtdd8bTdCgA7kxeuA0FZkq7d+m4Qa54dNs48cKQ
Zmp4cEy4SSQW0G8awAlcg4xoNwQuZQpw/5+9uOrWpXpJ/zbfz7qo9futq9rcZBf3
vAaikhWFbQ+EvxcrbFm07t2AVKwngvIV3gRKExZ+/+wG53f7V4ybauLyyHaf2roI
N2fdjEkNECEY2zBZKYrozUj3IAaVEZToaPLSOt2esaa0OWxZX+apjusr35YKO0fK
Oo2AW/perclKCg+NcqgsXSquJH3R/wrRsc/0lJmWTXEW+Ed9chmqVBEskg5thzIi
B2dQyRj/jPa+Jr+jf96YQvIcF3hhOUrVO0CAeslNzqnVtBVPIPq5qwBaY/noPBIt
f3m7FEA8oAuR0LW2d+MW4TOiuS79jUyAqQA+nB3JD101zok5x3QsePF/qR3D25GU
EfGIcM8CGAjWdZeiozwaBH5I+K362vA0BYIUpNt4LT3SFJsQZvR+cjaxsqRL8CJx
rLICX6440T0t1JzTIWuFi1hEH/QCFS0AnlJ1U56CsC1gEgMNlJGUyEsPeIbVZHsX
iJ+4wuxD/pROVmuYvtIrsukv7Pd6CPm3gqdelpr16pnmgcRO1nGzQ6HCawQWNHFg
biYYIDgth3FnuQjviqVknnfC3qmvhUa+suWDNaSJNk4Ft7xJl6dU0ThUzPRAzHnn
ZUS94duIcxiastuJWXIBAb8AtPDxzfzCNzJjyXOO5Cp+zjS83owZRpW0VDgEygTL
ERRH1gTiFBnN6Zu6/ZNngzcwhR9IgU06eqD5TC3rzVyN91EAwNRF3aO8sFTEV8Qr
366YJ1v3bzF8DcYNL4SBZE4OldOg8e1+wKPoWFWQHH9F9x3mPPk/SdfO1EKekG5F
dFJ4f1HaW2rcMo/gk8trzrqlnXWhdCdXR3X8w78bXhuhzcVNOAyV0QVsi8laOYe6
gsUgIkTpCPo17sem9h0q5mgn089t54sqyiecYZ4qryWqodMmSgLoCLeeH/KJ4F3z
3nC4Eb47mxIJ9cRz6N9lEcnYvFWV8s042kObvy0Jwar55W4aMv9MUPt8qEEXBuYC
Z1G07J73KSduxFgukMf5jA1Qk6NutJZbKfbbjLkPdf3q0B/kr8qKIyuEhntnuNCr
r+YSPhIP8G/Vz+WdGrvWxP6ZiegNvqGiRROUayItd1rp3CMsaZo41YVKkwNL9B2D
stF3D8EPUmHo5cqsuW09Y5tyACSGcz2R2aR1Grc/raXzWrbi4bWQnRN1855eQcuS
J6GoObFA8zI7Zof5j/WpKYfpxb15XPf2kZ/AD3NCQsda8c6iwvaAxyS2TyQMCPxm
kMep06NX+LOUfAQfqcZ6okZ2fNRlCMxl4T/Sh4mtSMGrGClA+yePYC/LuF78I5Si
IY5s30kXXJhnwE3RVSdJVMK6m1GKPGRrm1iLkZ/oyiIGPLL6cuGXUgdzIT9Bg8ZM
JLkvxXGDbg8Cf8e+rkJepwcJsOiTK8vqmvc8KF/gojbnh9UMHJmg+AUSvfAnLLAc
Asn6OIZkil8p22NSp7qNfAZbEC1KWlCG83yeJ4Gbz5Bydtk07zEZlLzkPfRBgrxp
jKPzOx9AKoD6xDkjdy0i9mHHWSNuwStSxCNRfMIRiQPnv/GOhNuYaZiC4bLNCFDN
NrN1Yqp4iG88oXH80+MwXTZiiMyuNpDrTsLYB+rscOjtTaX7Ae0+YnewLFbQD3nd
WOyGt5k2RZ5y24BTipRtVvwQVXpMobtLEgx+7Cpt3/TA3/aQzbzgW9AYfQ253ARW
JHB7mbiVKe2tJTKxNAi4vvCa9B2ofptO90iRAauia12IOhMCn331Wz460MELcTg1
TpQb3+SErRHBEuQvwhZdMIzG9JlewCNsD4pV5NZBpkbBaukLKtkBtnVAFatFELZc
oCYg/LQrFJ/MF++ZjVuMhJ5k3baBb8rE9LVpscsakg2y/im+71mN0R1poX31/l/l
wVyy9IuhnPpWkRrKWstg+UeqzdyKxeOr48yOuLIAl3XZLdtre5fS4vzhnGMVPRWM
8izJ7VuJXJELNufT8iZ1uF0SS+1kl8kQm0ZKOwDkCUibzeww3QNj7jNNgOLrbvFw
VAnyEXwL5vHAXoccTnYK6NE66Xuasg2AIx+MAy+SgIui4TKYVRe+HCY2wJKeeOE8
GW4ZTwZunm+bZ/HIXG9QZCSJU0ob8kqqOdS2ZG28cXGwJ/DHmieSmgXcSN6MEtRC
dgGOEKcbBN7JBAuOIw3AUEjbE0NM6WKlyQ0ajz753afnAOYJpVOx0+0hfEY2GLka
4mNeWzAMTtzRmzFQDR1z9b5kAk+Go8R2HwlpM1qYgyw2Iw2Bk8xo3IzQt9AiooHW
Snx4H8lLHzOXGUA00H+KZFlzR34Qpx3Yn3dW5V/7inIAhkZ0b8fuzpb6RswHdn6E
Bh6uuBmy3eWX2Hvf+LAJW2cYWYOCGS6K7MgVg/Okaa4LGfj/fT+fG956uXGHrfgv
fAnnzsBVpbelFYtQxswAly/coZpoPUdUQPF/cv6LeDsPDY/OFPBA+TedaY3UDco6
AqfPckCuTyplgB4mMz4tsLN+U4Cafd+8cNhH0LD/+iHuIaXU+huF4NINykjHXrOQ
Mryq1SKa8ig2ft0s+LJ7N+JSRgs6vaTBYZr6//lZYzfzFBqpTbS+vE3J7q+S2yTG
8vf263rFHaaWLJDCH3sFSeoPWey8lzKG5Y+HFV3YZ9po/Ztl/oX6pOVr8TKC7aW1
0s+UIUpTfLFkki4QHdX2/oRBBCNiRmGKx0ogYJjVh9yJrDtY55SD1B6CLQE2lgg2
yFhgWGFHrLlhLPXk6IOyTJ8up5a8HvHimi7jdZ8k5x26kQKvVlc8FoWpZFe5nRaU
8DaqByZWDWb8Z/n2g0TydswVLPvdJYB4SxmJ113ZJk6TQvzLZQ7p9yMItFfPgkiD
a8pdDtSY2Kl+alBNLTiQY9SgHKmcJkWRbt/QToQJQNgtsnxIvafTcHGBIqO7ZDbT
V/GeEu4asfgg06BqusovvEoYB30nvcic1NQRG0QcKhgvadApw0/ZPF1wF+UmVIMf
Kq1KcNPflSIQ16eKF/baf9dcGX9wzrxXnS2C98j0CYo8HSxkqAu8fbVwqRfAVRTI
xrqrdfQZ7yYm8PV4C/r15zVhe19dluHufBIgf4whB6dPeURANfv42ZyNruMz1TBu
Evwfzm7up9ZMeF6SM78u45d4437ITxgocvXpYz0vByXzOYowa8v0ZB1/1YGRL9GR
XSjn4mIkxFmCjec5DarofLGyNYKZQn43BoWGtGKRPle9yNbjIqrGDrviyFthePIg
8iIfVHOhBx0pn5mQUxwEWRjAiRmFfjb79r+SPaYQ2VReSpd/qeBVuFWVVpXwnM5Z
Dw8c7BQUuAfnLLgyrNcQncrKHm7X2PtFA4sITj5jwfK6eM1RnC4sCmDZAQvAKsYV
6x2UBrjg0EkmdU4OndpbPvrwlYgEDro3/dGJRqX99NNBvY01Kjgw6Aj2rHq7K7St
UwfopPXOwL8GFumjvLLYuUMmbczHKDu22xeBsBJakKuv52KRPDORD7zP7q5Z37Nf
bfR3unwnbzCF2Nz3cEAz8jqwvdQZ9vxPWrd60QcT+3WdojXjNL2C8XxysIXp9p3Y
KmqTHVocsvc7VbQA1WtRrH52bbMBXQC+MVTrRO2TJGSaczMGHXAIR7/Dr6lgdQaZ
NR7JbwU7BzleanaMkiFJDoRGqD9hN9C2uQPWgfklH7Uf7ykPgi+1aTYJ+X0+2MnJ
xcr55n9Xi2HluoKgLm7gMsAPYwbcxZjBzI+CNLDZT70JtsJ4regMKYFkj4zNhDE9
MYFu6Ef2iBCjqxQKVCeGwduao3T7jCK+v+CFBfqSjE3QfIeaZIkLEPfwCHTYzpUa
pM+fXNKiQF9hOocoER12IeMy+GGByJeual7ENn8lFcWFXhTVbMe2BbEDzAau19QR
3u0/gIJUMlMxnUKFAPZwFKOX0tAzZ58lxFb7/rxzxfsOdfm8WJMEc8HdTeMPPPm2
Ku2ffNDeN39QSUIGDYtyD/MGga5jmnpSkwmG4vRHIksKAcYAMVgzAI86WyuNADzw
7WmSzWdIKFIq5+246+HndiBDEv2579w66W6c5m+tPd75k8P4npJ61fbD8Dr99d9K
ECoXk6RGQrrNHO0HXhClK9C5fQ1J5LSerUam/dymw3HH8r15PizFenOVPmV8cce0
ZlZVpujdSHw/kgn+W7ou+o9N23G0FbbT69wQhr61qRDSSOlSgXLNeNznT4fTHtSv
EkcjNtDno0mkDbJbLXheV7TSLodnZpMZE/WIRLnY0Gnvu8xxebTeMIGfDSIKvgH8
8I980mi7vf1LBSVqokZ6/WkyqiVggL0BaXC2xw+5RnFwaocNTWSrXZvxtsGe/5qN
VWkNFzgBaWjwhrZWbgpL4M65/8SMMQujOkO+oFEFeEbyIxHFYze2Qz6ojWg4Q2ym
6RHrmCe0lXjoVwH00cnQT5vdC0e5/GtsruPpFKCAOyqpqp3Q4MKzSbWra1xzbAOs
awjCCHDCTZfXcFtrWypHqkzhgZlbwhj17Id1EXV8HYcNtFoGliPzYjrLB8wWL2Kc
QA2gPo2UXG6RfifVsH2vd+TG7HfPIePNcjBigvzMkyd1NQf2TG48IUi247fMki7b
mUYVkJkmAdXIIvYo/RtXeLcpmiwDh8/YKMsZH7Fh/nNNh9MgUFPXyvlVmDCapLYg
Gw1+70eKTo6sYrFOpl811SXtiqBUeXuwq2gRvA+W12RhQgE/z9LhIxMN5PcJuhyV
t3gR/8CX9Em/UZOcsBMv0LrsmiBD0qLQ+n5A7XdeMr7h9LCm1lP8mx21TzAIPC+y
d25dIQy69Z020cFbwZeM4RBvbwNglb7YhAhJrffC1uOAqknUVE1REFFjABhCqeVC
tCWNqvMQiyejpmClvAH0MrmbYHsBfq8y0qx/Pbku4uF1sZ8TGfk3Mro+GKTyXmH3
Y61w3UQleO5hw8VLCN+KVmBmI+tC8D7Sm+xXfkHQjtXGSHCMtMakYdVec+Nf7S18
zeW36lo2z1FlcwLKjVxlhTODhsU4thflh2+g3c7engWhiVsOqtItwK0BKotYyK42
k7fvw5iIkbmaUW0F2PDBKDV0pvchvSUez4DY9wObQIcarD6LNrunR8EmdaYSgft3
grrTK/wpCxEXctiCchdU7IX/Aq/7clTmY03UmDwWLiED7XksMZNxNZn9o1AI9zqb
KSMLIhKq5huLImJspAW0hBP8coGLIa9Yj9x693D15RK+Jy94SNz9ec8mCxKlUDwr
6qf9U5wRcAnpxFyBIOUz03H+aF9CtVqSwQCbobNvg1puj95Hbjre/JCLF70r3ETl
qnE8cUtXpce3KQyjXGyYppl29CEUNms9sDCEhxcUfE9naUkupLaBHYsqZcilJ5dO
BM09dTrk6IPWBhQKynQRrBSoCKLWBBifBM0uBqqnHXq5zKD9DV99X/K1MjrEjuMI
gTTl06vqZ9wFp1S+f4RB6rgCtXzsD0Vl3fVUJFp9rDRnGTzCEZVL1RWPpvgJOiEv
P+s/rKIZtWq6oayzJhKOVrK93VETzT6Ycp2Noi3rjvH2iPJ7TpEjPNglBtoloM0d
CoN5VkQPzV+GGPa1v1ta3nJcUEe8tLfbrsCL6tOoqPuaZdiB0MIjcMsUPFSf0zoS
CyTBcLy2ZoxGCT1wppceings2Wg+Ax+BTPNr2EGCrafiSLvi6qWs4av3B0Fv9guW
Xh008K582o9hguyPnwJjO47Xnhxhz0LdPwyTDTsrj7ZTF++Famrqepj+PIL37ZaB
18zrQM6CSoph4qxfOnhh+oLwOmW40yILkBtIFfu+AHMQ+moxrMcZFH3BvLGVBtFH
CRtnFhGgcQut+9zlZRnm7bb0RH93fzqucaVIahOJ+FNH96s++8v2KUpV4YqkFNml
qyb1ZQlSE1+f50xGVcJ29VDTIfGh5F+Y7QESU/hJmqd4CKGrRZETlH9GKjIcW3PS
PdoRZ30OtJrkWukWjCV+FAeH3Yqtcg3tRpNUD3t0vosi3Q2ZTVYH9RuV3rGRn0Iy
X2AyvHmYAj7/tSYiyra9lfnDioQqZW0YUcabeuqlcyvF3n5TW/F6ujZjIo9Bi9rl
mXuhaXvXPvXEW6FnfNP58Je8oGydntJcpzhuUMeuSy9OUTv7SB7LOKRHnKMKH1eF
IDzYQB4ifYZ6XD/r1ErC8iwlshnKHbgc5p6OjDKxjNURs9SYXgqn9JSK1plks5tu
lZHW4JUEaE103WbLvnSUnpH2TUGggaqQFSyjbXoitE2vdVdhYleIJVtDq2UhYXGn
JueFGPrVIL3OtJo8APn7o8m0+Xo2c8VHLs+wBGjpiAwPYCcr5hLiRoLJt8jGFuGu
k2pZAE5yzj+nhBzmeIBJpXrtP5JYS4gjRelO0vGASZ3jgJTGxhD6uZSYwWtQJniW
iyVyhFk5Mwzjqin4fh3uVkGcW+Z6OzvpIpavKZb887fAxL4LniYsOa8DTLwtDMYU
EXQJRt9ten5SzuTMfNBGfbqTDKSO1Fo36VQs1QVn50avtOYLstjFAGw2+3p+lmoJ
r934ouhKNQ82uGo3Sua7mq23CAhHA57SqB8BXkHi6ZS/W5EfCHlVSiXeP2t3uvZG
JQU5eBoQnITAcmAxvTNfpHlFsQw4RrzqDjX+oeDWj14nXa0+tERmyM0L3I5Oi9kn
T32sgGs5My00IzX/A8EyZnDmT2XUDGfuvfvsR93efalOUcmAISdu+D8OFsANbh05
ccN52ELTep14CSdR5o+MtPBlsqXhifKeUzLuZz5CiBzVR/aMHEH9KBz3u/0Gmnpy
TWM8ZOLiCvDLsXfLsirVgtS4Z7UQIlTDamb/2MAKoVNU+rH7V1aQUwBqobcq4eAb
l6Vrp5Al3AOuGU16nRINSXIjbeVDShxFP1KzMeAKBoue+IzL3BeitxmrRtnNeR3I
Kk+9Mfst38OKlv9/Ypu9ahEQonT63h2TWFEnYRYn3MHbTKgJVdjCq4zoJGRH/bUT
AiGzzEorQFUbKvLMin5e8wxIMJESfuNspO5m3PHZ+z7Fa8RucKi6oVA47TEFLjCO
urnF+fv+zixo0wzvUMbWKWuul7RQ01VK2ot1CBsnepPO/7+5qZ+rJLcliqv3hxqz
H0334wVc+YB//uZQVO+rZh9LjENP8w9A+i/wd/UrvHwALZye8oUkqXIlwmxt1+Q4
QRvNa3G5QFGEBLsJBB9UhT9x35Ruk66FFhTiZjQs7HbZL2IhP5InN69OE4RHtYrY
cTPC9JU1CsTBCj6uKJzZbJUS/mCx952F2+GnCrLGsu9kHlSdg48TybQXn5Wckz8V
T1mqbUsmaWWIR8YP8mX2byEdBsxqaxdVskCIqDqUxRYQCOVSaGbFwgsxXca0aPa7
12Q4rxE4LAReY8NcjVTOJjpf1/NoXsXQuDb9wh57LFcdFPaVT0F9YTRYx76fgmwH
Fi5jDg7agnWVybgLyB4kFy6r+1IJiRJi/hMpe3idQxwY2s/wX2cRygnHnqacIv8z
a1qaGqYzxh+XLVmADrhJch0uKOT7S4po3fMIHbdT29Dr0JVbCl/mT8Y2JpN8XA2j
LelYbSNyVVfuVHkc5AnMhCF1s2wMst6ps1wu4JbHUjfwMz4P6JRtxY161ijpBD2y
VBm4mElhRd4vtwRQmN82psdj2z3LPxKrkNOr+eaJbTI9qRTAlE6/X4TLEWALq/bC
wrT1sxkJrgiXPSMy/JBz6mW5bEVLnzVeZJE94W+ymSO9yuzsmvlcNHn1RAhW+Cfb
Iq7iuwyOZbRlXgcVyPMHerWBtCRcQgPqmO1qbUfc+cnQWkb79yythViZgKilW9O0
V9A1ZUMMrVULkwOMG65Ay5MI65QOhtFXvgWG3G7yDoXo9pgfAy8PQsyTXe3uErGx
5iGJ8rC9E/R8aVfhl8IeM7DLJD5xENqm7q3QEdNvU/4o8Jm5E8vNbt+sH4InjUkU
DkyAb+0Qi7hkKgglmq4hDg8zq/U275+dRsq02pQgoAUVYF9OxxGlL9E6dwxQ7pY6
G3hdP2Frn5lgURaoFBXhD9sV8k5H6dmANmbAea/L5dqRMTw+D3FLsFRF5qpklxQi
rgge9DwsvUXcouW8vvs088GTOFaYXRUphX6PXuO+3mXzgCF2Z+s4sCsd3jCSlxz+
IPeM871rozRkaqjgnUOCNvk1jo21X3O4ff3VRDi/X+b4RuOGvuTeAKr5vxkLr2ct
5ggE3aoANGBB1ngfcNCkQTf0xDKq21x6lPaI5/UyOSKycijWI4+CT9G59BRkJ8lM
6C4YzUaxfjEvFYjdX1HY4xzeqrffCBB7FyC9dtOjEVjpOTVnL3UzgM0/ukAUE8fP
Ln0vUYaIFQ0TjDen5lvap1J7GnAhbQ07l3Mdn323eEaQwgxeAh0nEVPzSw3XbzIE
eEDVzFbBJLuR+Pgx/LGVtyX8z5ux3+tcWGd74G6peC3niH7DDDFB2p26OB8IqTmk
2VtijORDl+JZJfoUSVZSoG1O/pwb2+xtHZFo7Sk6aBCYQULhzZZB3ekeNU1Gi8vU
lRXSBUMnrqIEV+2VkIz4z5cMizvlacEg/6CldYYlWrtK4ELGC6JhjbXkiPESfPXQ
vi5DFKq9p5rDTW8wrjsB2/2UNTm/aa7QhMCZkV6XSkFC2dUpSRLRtzlqb8ani5QA
5GKcqIMZrKB2SXkdOWsLbUHJdNN9xgqE1gf3OnjJkdi1HIJzdJJHyqNi32IxNibQ
C2xTEYOj5IZR5RIBiaQOKxnZh5jCPph37tf+37sv6Altp6N984rbIaIxE9Y8FTa1
JqkmkrauQ5ktGB4gE2ceRuRo8GZGTiG+oLl1pDG94bEvrE0/oQG7KsMAJ0/ADNhF
mRQzunHbJNCZ2OUCL5Qai3Qzmw0CnZF38m3vD9MiyMBsP4Eu7SiMB3KIteOHgKCF
uc2Zr0Tcuxq5lxHi1b/FtFDxm4oYSFYW4LF61HY0vzzqmPal45jgu10XOvmhfpPr
o3k0kjx/E4Uw5yyQYYXVPRmJ5Ki1vtSKBVyvj5mtEVTfmJ1W85RikZJgeAJm1kGi
ePwJPyOpCXVuFqhHTqgfEErdPTbJ9U5MPviZxltxnMqJbfdBcROySx8j3yHzIvr0
pmd2fcqssHF8OUUN/8cJwW6QQ7Vam5jPKOMQZUzwW9Yz8r+T300j1FcyoeQRM2tX
EeqIh1EWA9I/0ASVxvAck49cyDBwKMV0UGD1WOD00P7XOWu85UktGgfRofSeUYZz
j6c0bF47EbXqCqodpwE9Ir6To4YXYH9qFiWDegtAGF3jv0XH8WuLSiUpeUP2uamd
AxNAwQOZCn7hkvmQMZFXDy2X39t5SizxCA82/HuMXQPczEuMUR5wCdC7UI0L7klZ
8geHWMuu95tnFgJNVjHtG2WTkK2iI3ugpIK0f9x+fuQ2qus4OdYtwirfAJ67fZOK
53CXTBYd37NAGd5oDMxMeqogwGFfAOUDmNDgciAVBdNyH3ez0JvntS5L/rRis9Gh
qJBkjSnhZju1hFsJZ0RypMFp7whaZ9TNgXOqVQRne3MBq6CrEEQhOOhCOu3pTmFf
MpWJkMvZ5rLhvtaAzlgX0ENxtvAeXvdOBzFMrArfUDpMtzvS7xn8M9ysCvaEEw/3
z0TdZDwhsdGgcOfzgUya3LVz+qoz4jhthOvcLN4Jfni71DorrUXVOc5d0q6roYaD
xff0cn4kWFTSPVkmX2vQ6iWCcNraz3GvN8JnHOdM4NH5UJB+g2V4oyYXrUoCaxKP
puJO3jdyYPlPWHNIJ5T5Ur3qI5BV3VLcciza9it/Zf6aGFc+fFsN26eQxoh8Y4dU
c7zmIUa0LYA+wwNwgSxgr34+XCbWsS0d8/uhpKuHwdsFtsme39RvEfpZLlt0MHg1
CKm1tQ83/p08DEUdUtszBiBg29iz0J1hhhKTVtXENrxpvdnDKPqfNLd6Y1RLjDih
b5GDyrIM80ykaXJkX0n4g6J9iWpfxXqgkonKTJc6Js6fJhpjwpnL5O4Ocs7/xzPO
MaQ4EOfsBwiPbg90zC6aGdCi72EtP5o0gwbMzoRnb5O8f7lqqS8GGlR9YUmml7HQ
iZAtx9l4PQEkY+rbviWmEXIHyvJumBjQpeQQUp9ahmcI+EiSU88DuG3FbH0EHWdz
iI6O963x+UTYo7s6I1MO7xLWSeI64dx5N46la0jE8ESPdk5XJVHxyJdVgbkJDJWV
xeyEaCKTPSLbRef5dSqzjgM5Eh0wHJeX7DMjQUDiqyQJWPRjSJ1Kf8GLtUCN3u+v
elfC4YDy0DdpPTDD+whQIhA48MHo0k2p8hmdR7EeDKY+abKo4ZLSvWaM5uSZ35T+
IgBq9GYH9F6f72O3IGPISCvNZJ3bOxDJfoFK5USsBoubQGnljLQjcHRi/8L/1aC8
RWK4iu6drbylkdpMsstkqq4r/hqT59QjIWEHOzD/wetJ5S4mja6/GaODhGoVSkPi
DDCUiESFd6cFW90jApODzDiEtZWUgaj+NKLt66RjzvAI/JqBwQuI57VrxKm48DEd
owdTlRs3Yf2a7q9+xl7aGH75wOnDxSYRyo3P4rGAy3GbwkV8rgzddjuzEMDg+hIQ
Od1xl00PFTplrdn2hxXpr2OxCzpnBQvFXtZJD66G4SLEsSVHGT2nGJKvHaOm/K8A
YSchIAVDoPNVavOI27s6jISylC0lvGGPX452JXE92Hqt1olYHbkJpOaJVNbFUzY5
3xYNIzGYNT5DE5RRolwME9ejGF3/D7LFRwuFEzvv16+dBvI3TBdsCgoi/EhpYP/8
fQpKRuSgHDZNsJ98vdHnO6LegdXf6rrBnrC1gpN5xXpzpxsSVIhJOfpW7HYs9I4c
OqaqY6XoNVndxHkttA1165Ct81g7JGSRKcMgIhRO0fnE14BuBeyh8ng+61DNmdlx
eX0/BiFLdTbk5OtLKTJl0D7CVzaKTdExNX/LWF9LRPaQj/NeVOfk6MyGx6KJpVMP
TK+rx1RsHCV10/KFZFLg2AWZs5ndbHjd0RLk3nc6bKbh2gm0aR/GEXFHlPY0zLw/
0Tq0fzk+/RBPB9pTI+EGfWOG0B1FubMZ2TQ7gWtJQXuqxpiacGT4hIZRkVSqsgkJ
sKRn1YIqUoONZuHJHTt1yoJxLiNJw7aeZtjR5TrdSSgB+7o1zMIwQOdvmhueDAo0
xr3LlJlZCJw+Ux1KpPrv3VLU3N61Dl1f0s41JtxLcdgSW07E0FA1vLuKbVtRKZN0
ejpxH5VDWGDvEI7q2uI/5YMSFo66BvmjaD7HVZH6zZVcVn90vkL9vwapYJcF3tTN
rUjWCrX/7jMjnAuounnfQ1C1SfgaWtoREtVkKLytfV0qD/aqVVdSs1xDs/N7vsBP
i9CSlEwiImsw05lJUTzz6Md07SRhTJl1kFsYSu/HhNVqgYN7g3yXaedHJRpL9Xv0
G72L94z8N4VwpkwuXQeYAfaOuqHs7tU43f0bxeaoT6ARpQaXJN1DxkQZoVYhy+2w
li4ifRSSKmTR5Gpv8zT8kdqQgURbWIc9ijIO+Y6YDP1ENZpq7MstqL1Qv3Z1ESfD
md542+Pq137Pw6wf1PyrQtBP7a22CELzpgku0+CF0a/iz+itXAgzBJJTn3uwytuf
Dxp400LZIB7UhSoSKliSOQ6X5IiBneF+3MYbTKYIZXxzEkVBuz8nKmUfZuFfgE0b
QTgW+k6Ybnr/yfkgfwJUbe3++4YaTiEsCpTTaJwJByPQLtuOeOQuVS9xPB863mmn
VaQ8LhAYzfoWC0LcL3Y4DsWtrI3MdH5prLVdI5AeLlBLls4s7hzbP8Ka2xUKLcAe
+tiWSqxmx4bhK/VbIvwKDFiJjCPTjLd02tf8vwGL/LZibT0rHV8n+2m6PYhXbfA4
KwZJhOM/TAVZ28EYYxoYlCyaQCIBOGq12e9POXJSdYSG0sscXnMBNW3n4pGHnuMi
SsKnJpFPLKFdE6eQ/BI7lA3ajs8eyEUFwPMkgaA3dvFS4+A3k7MuWcMyfN9x6O5v
D5JEHnzT4OkgFQ3nJtcmMc4r6fKRH0B8InUEpDWvTBrBPdRnlav8aCJ+RaCjwC1s
6TR0wvt5Uu6u9GmcjVjqe1oOqrl2FzKxIoEYsYQTMH6ZsAtw8MKhe/6g64XbWxKD
Ys+92lnhT4oCiUvHz8xetWEeSRrLqfhNLHhmdew80YCeHOQhjZ56Z82HFTy7XHra
gf+jsK3tXfFVM3EV6R2uo0Y23lL2qPB7a6VWTVpIOpbIg468VFX0+pG0zT9mV7zc
aIm7jEklqIPlZH2u0GfITibLQE29lG5zKcGWRZ9z5GBrRpFUyw3HqrRut0Jhnkqx
VQ68gf5Tt+eUchCJaqKpx8b9/IkDBW7zZgQntXlHt82w3Gf+GZwF1liVYcr1d1q9
s8KN9/6j4xdwuMa9P8BAwGEZGN7gIMehlPy1wlW1gry/58V7aBIqExtprSE/MTQ6
6dVca1tM9FsyfFNaIIF10LuiehhKqyMOXsJ+vstzuaY68A/dvqspnozFgJYBLMoh
hxUX7Z4Km+ntv3qsMDACMCUgB/P3tGcBQ6uZ8yngY6ejlgQ/rKeePYa3LPSkghm+
blc0unaEXVwVdovPwzr3qkkBNzbWoTNY4DdYO50w570EQjBrqGvpowzNVMcToXMH
Awx5s8iQGtzzhZAohpAFepG4DQbylArDZbbqMRENiJz5HC1CodEZXCKJrevbuwnY
Qjc5qh81oYa0ogZ2j+bJaJSALjxEAq0pzrmHphVsnnpWW5ggEyhG79wfaiRh/7sL
qLeJnA4dhy6PpesBlWBgZ8QEQClSVg/JC0OJhNMCHrEEaoE7Jjv0gxZEvt+Sc7Nv
/JFmzz6tyqjFgbU+SQ0faxKwTFXyI/egMkGqMpSybLFUZChclp9nKVUHkOzEnJXY
XIukz0gK46hbxqWvYk4TT/x+7tREurcx4UwbRMuXuK8HdahEiO8irJ88PnjdizgR
UP1r2DlTtp0bmHPcWCvNvmoBZxQinWw4zjhVcjtVSXwxdQsLS2+iNorMvxI12/nX
vbGCgoDTarAnFVifLGVWMpRICn1LJlMMDctrDdHJEKIbrUM7eWhYrivaGZKcricy
C1yoNBClx+P6RHjaGaBknW3JYotbyhIUZB/AmKU3IyrwEwUKl063diXQS1Plktxp
uoQH2YZH+wCRNZaB1sLFYmvhHoWA0RfLCbZx/RdjDEFQ2WdVzE+p+1h5vNfBXj6O
H/PBVR/VBJ8qEzrxVxXOtsm0XXbjMxMxCHV3vgERkHrupFGe6m9BoK9k1j3ZmOlQ
smFrhMgbQvxx3XERMI/ZT8jeLB2ucB0FNSWO/N1nYEETjUX0k/Qm+VTwE60CacUu
9UdMBnNNKQTUMncXaf6dqandRL90Od/80uwlP9JRnUZdPnEzBOJ3XbS4YeWmmGNr
D6ZmAPO/7Ee8G4KKNnELftLJiFAsUzsqsmNsKOYaZxoXoZ94v0HEqQRSU8PTGbvG
lS0avB/vHxJc7WzVWDkVI1kOih8QI7jbfh9Y8TBiSX6y+tZrvFUhKM4ZpZY7RBKd
yUmf91FRDcbuaVvB8Cy10YVss4yegqC1CxTOZdXdO+6t2/z/jX9whdCz+1wfvOA3
2oDAZQiG1G6GoQY7bHU7ZgJqaWsZqCi/2XAs+Rql52WFXXRPqL8DFoVs1mFtAasr
uPB7S/gfMdLvVxdP7jZ5ryQeOg7fsnMdlEkAHrQtif6za0VqY3gKGX2jq0OBO600
ogqU+5d2bTOVqAsGX/3mzpftpzG8jaaIdn9SmWlP5Kxi6W5CduBh3aFSrYwyuXNY
FVqrT05EwQlRsuTN/k+g/tYnXgQdpnJdhP5pCMLLOjd9IFmmXYEzUASWXy+KKUme
fKeCFN39vEf7PppXas6N12PUSCS2XDDHNldnPMOjdc1EhF9rgHCoq4CuOuZ62CRm
xEx3/88G311LlDAJcn09spyGIggk9oTV7m2zkc7cEo9XCvFpNzFJnIM1ZqPRLSeM
m4NHwNKIULGHy86tUyMh5c/pXdP3nhCxzj8fA1iJfFxscU4pOpvHPI5BkcMVNXMN
ojswPCUw7nTaV6UNr7bOfPhRtoNDr3h6z1pXG8r2BwxTEgYq3d00yDjsLPH7vmUK
vL9w+K0RCGTUnJ6pjnqqw43HCNoacImkzDdDByEODid4lrv0J1BagQcX7Z3yzyVj
5WIQJcpHNzIEVW8MhlFaDGwl9NmrGz1OUxx8NF5UdGntfurVv+PGOsXor+3J10US
6rsT+zZeoW/CISJM9j5QYYbf2dcV+47xF9NyUvYw/WavN7EgCCQT9zthc+gDtLiY
SfMn3KMlIDKZ7Qvw/eNtwcM0NBMmLExwE5+cnCXR6O1QOqRbwqAR+Y4edDZAWk0I
rwzQdjmx1uqiZQKNFUQWAImr4ABA67DbIA7FIq5YWsOuL7+gj9JHsTA1aECG4qJt
wKz1FaJuUEV6vUZfH2WaUAGzPTusBCwzRCKrLU7K3RScMqEgthNWCc5Z8XhEKuOj
2WAzJ3hiasnU6rLg3CqBpSC0KC9J6/rpyvOgHqGaj8Er78fXXaDxyZ2YjgS5nBqr
10RJROEL9Y+/dJm4A+gItIS1QWKyG+6ZvXa2FpUu1fwivYst9yU1jEMJPI3yaHDl
PQGYpC32us11yTPLk7R/TE7QhSlv24fzYwi2cHWfEba2gbByV+g0+fmeSM+t+lq6
cl8ULdjeSxX+cYqXuEfBojWpAETmhWUMac3iYZauTFHVBBEE5fse7Kz7fZ3AhwOr
G4/gPQcc3a0Q+FZb0I0ULodrv9mv4aeLL9b8ulqBLXq94oV2CsKXbFPldKA0zOnX
a3s9UcWgpjWVQMWt3Zzmn5kZRxfcmI4GSDSJrBVYLjYWdAYq79s/G0ubsrslMy5c
VctlTuBNxeMVNaxpjCIQlnZ0Eurb1adfsG9jdpYClvRScvaCBJktzQR0mEQAbSA9
uebCh5q+0lhIKSK2HTQTT85ePmjtgkBRl+qjf+7M9xBiYnqYrtiubcP3e5d1FqSy
a9cXpPK44U2a1TA0ATgoPoKB1sLbXa4km2J9DdpqIxOgCY9aWIEFVOLX2qcoMYOV
MfRdrLqpo0Y/AhAkCO5Ze9RZ/SWfdp/l4UyX2R7wD85J0BqPaPtuN/VpVULoLhnM
3ladamUrZvgMus4+EtTamj2G+hkx0kX65PprFvcXGyfu/BNz71N6FLdpzYjGUsrc
NHbgrgl04Tr7gP3oC3FsNAOo5W54xb7W7GCfJuOdey9fSdMBDpOonqzOLr8J0XBe
60pUbmCrQNwcv+jqAz/d01ME19uBPoZlodeAvUgeejzJjpzI2kypf/EG1yNezBd6
71vByO93xUrrjr25NCgGHwBA2SGomrS5eydkkkbK2Mv4kmlslNb5xu+B6NgwXAI4
Cr8fPl9ScYPvZ+eCE1xwp8tM/HxrvRw3wLCLmf+tdHG1BdPJOYu77RI1HNvKT7l9
hnKtGYU1N66ym3NPkfpahdZPmsntfMlQDA1T1UItmPefXUrHdkWke2hfCBXOfYQx
XzqrD/3Hj8VNKak8b2vDkb7CWSSUsKycQwZRF7mu7L7V0Qanl9fONXgV55rvb7bm
DbFFnKWgd64s2dJLhj/lozAMrvRmYgH0a6Xj/opKq9gSHC2dKEcLnv9cbYaAjd1Q
6RMZWMziu03uwqBaUeNQ4TYUbW4CxEgBF1Dfcfe7h5gytYu23gPYouomOxPV6Bsd
0k9z5/eNrznjOg/92+oOqYsYi9U9rTU+Sd61vxKVgTUjQ6Uqu4+oWKErz+Id5Z4/
GsF7UdmlwmwsJHTIQqgW/dXpaUvnaVknZ6PSYGSQH6GaqEW3cWGiCVD4sCvhwNJO
qVf+EHxFbwsJuE73mP2h8PtWhCsVY/u2jnyyMBTvOunxoEphOGXL7cXFHnJ9ntyk
D4Chj07cec/2M1RXWy/AKoAjyOZcn5PgIDo40BSUu7M/Y55yoyUybh1Ou+dRLqxa
HBgYNhLVwM4io+yTb36xo8eBqYsREm1X3UoRVwyRlo7DRs/+COlrprbKn8wt8AiQ
IBuCJsNel9dPpsOezr6vamG+GstCULozRNHOkmApd6Lj5n2mHAcKrPCIYuN8CRHd
TFk8JIXdcKEuG09yey6eYXDiRnkUv8iPBagMlT74hHHqCaAJsKyy7YYGND8+UC/k
pBfHlJz6E9jLzvhQmOPWILBHy1gLiLH7fmkXr+l3mFsmjEucL79Y8MNE0kU+7kYN
9NLi8/m2keWsBidWMuS7UAAe+dkszPgxjLXOT5NSHmb5XvtwwZg4AbqZL4OD/Vcb
EmzzfFfBL71N08RV6q7Mmzy6Dc6ZncMo8Sq5ZuiTZgGqPWY5JNurOMgkH47DlbaV
nTqS4v25vhmK65hbi2KA0NqMhJAFSAHgNa0sB4atxNA+Vcj0Ap5BnhXrEuf+Kwpb
Vgdle+KbfPGzrLHxZZxuDvrkX/HocJL/sa65B8Tzj+zbaUvK02VO5Dl770CDB03z
e7Ue1fY1Bugixuz/Kt1mEYP/59nplK97KNT6GDwUzXu2TalpTqT7kJHJ2qSsKY3v
Ml+2SWD6zJeStVRWFwBMy5gGbaX+JgG1/sUo+EN4rCbObt7Up8ulqsHG7/MpDNhR
hTt3jy5PeWMR5trWDhcsMzrYfSeZD3WP7KqwsvQu/wqIK2UqlH9dXiI0sY/IUTgX
1W67965452/+mPnPubrNbNfr9B5dmjqyY1JQCDoO/5jmUbhL5RAKvm0ASkwEzrJK
75PFFSL2ehtPJXo/v084zea+OrGQrrimBKCm4QWzNJk0+234Yg/isFj4E9QUG9Jc
gEDuIPtBY0Ib4BqT1WP+84bCLzamIUwLGdA+TGmfxcFIrX/rzPVEXAl27XNdamp7
rcMc5EeEqQqyYRN3VYom1kG8J0AWgGHzYx1lRfCBq7oDu7sg2o6SSkDJJsb5dEsb
WWxovSmWDxcxgZDKobNxwPoEypevp7Bm/3Onr4bEu2TuRiqqAaleG2I5fNSIrRgi
S4yR29RAhcHSU09nDIvKybmEoQQnBD6b5d1QQIt32vJcAAsb/JpRMwAb8pbwtKZs
5AZT7U9aXGe0qnINzno63l7ClJW7dqihO4S43uG4tXtk8HdCdTX0l8U3gKX9voTp
IktgMLAl52MZihpqrx88jgVtaazfJkudSE6ulZGodA6hjIFhoeoLR9KTiYkQXw/P
nN85HSW+xlTvgr2yAj8fxT80K0jib7XPl9UbdlDy48lpX1sJfp/cALqsE3RUCSiF
TVZeywtCsF7mu3fFfmA8Ts5pKLBd3ogAOASaNdImTFZYoxGwDBoVNv9+ziyRE2De
W4cDOdSQqHVWruo4ZKprh1yD3yCYYp6b3wVeLg1sMwUgA851yk6hUg5QhU4ykgHC
9IWoGNS2MqQ3/FsbHr4yGqIJXBQ06y1X4kE0L+r0lUJ/MtJOfxxAwz+kripEBVjY
rP1wK7iEBkEWusYKkdr5tceMKzJWi2/KaHOXo7YVGDv1h+bHRfNCN2w8CPrT/1FG
Q/hGGDJ5N7B82LIBeWmhYbkpORNdn/z0bqSPaDpL406Zl+IGY1OHBY/5WiqQWdl6
h0EE++IzFP+Cm+nk2qSGYuyICFWxMN/zCjuoCdxWRzLdvVr1eAjy0Jq1a7IjUxB+
mj/MBtF9xC/gkXw0iP2MMRDJDy7TDeYK3/h/d9mnHUylbzgtPgtKhlqDW1/iPJYQ
jyNfvhTneCW3XBuAjEHZ4S0f6/rsgbSQIo8u0wauxNl74FEucQBIAmXN2FT/jd0P
x2iILYaVfK/U8zODuoxPnj/lT/js+4sq04z50GqsyUwbNraR3NZ36FCfxWKu4Jum
O62QtTArlUA7+XcOTgC5TZeqrB4f2luKvhC+BEpegTi8EJ0uKaNB9STz6zClLRbz
0h09EsXMStc5w0c5dGLGZ7D5O6lCit6Pkb+XmQmgT4RsHP1vFo5noor8OjZU98sD
mVRJXjWHELC27N0v2hboD+WijOS96GxqPY+/TzvvhNQS9VjmNVInHRSGsSD7x9wY
fpOCTHyPq62VlgydFzZATCI802AHssA5lYVNR0Yf92zmYwHmEf9gwrsJw7njmowy
cLpYFSYrePJ49oMAwXWb03lmgVzP+gMdXzi9KoQAccqbTJS7M2WrHKUtHRvtyKCM
uu6qbGiilQi6bManR48WHjP5EDUR84Y02qwjBm5TVtMjLBH+/krxUA2hVuS+q95R
m9nzVai1E4xHjWS/zqaY6IO4dhsrgrRUvY6w9VFfW+UEtNYtbjU97ZXdaSlLT2hd
gCX6e6wnYZQNZiaiOK+ivibTiY8YPy1sP7+pOcpzTdB3PBJ2kNxtXVulEXGqKZSN
3mG9/9sRbNkv5Kyq0Mfk7eW2mnJWaHqOTDodiDJBOn94Nj6OssqC/iwIjs0JbhUW
m1GKibNikgVY0oHwJmxUHy///eEhBTHJoUIyfMEniDm7cVmb8DO0vyibhejTHCuG
OeKtHfoJprmV0UqtlvFLDqGboVWYuCie73BwUdHHya81KsqlfnK9slPPqHReY64P
Ugyj7kZJiJVfX5gxlNyZ0CxvhiHjTg1OatoSRoGDrxhDqC+P+Dr9R0fiW6bi5wXs
tvf4OhGAW4WVn8QrS/tg1kSqKg7SC7w7W9TnFLo+0C42J8+/8dFIVnTaltpwK+8Z
ImAui2iAIEMWYajhw1wsgUwcuVeOay10MEqH6UUiVeRm+IWi1RbUaN63JUzh7OaI
T9mXh/fRoinDPQyd8AzbmK8K57412HE67XS5vf/oWIY7MY14bsTFVRikzsGnVs1L
EcROn/87atPlOHYTTU0sgbxQ+AVAJLHFfA0O4xOabat9R8h852fVZflrQ9IjEOzo
mHVuIhmzi5fi8Hsrr1sdlGWEbijQChig1EOhCkUvebp2qd+Ldts+LjcyaLLwk++O
xf1ZsP6adXCeQ9Rfn65yMTrFbj8BpMtnzX+uWRnkGsya7uScRq9bJqgYmSlFVn06
b0+qbb+0CA2e0dTqdATNMDqOr36zM8dazP1eXQaC2Pt0Ii7zuXsTqmIrVsmyW9+t
S4czevwNywkxyNaBwc8zf2jnW3tB0cSli9lcaf9ixloSfr42ZOyNEjGgErc8RTg0
6pndC7Hx6oLLmMldB90RlDv3G4hvP4jDj20LzU6C+cb1LRdA5Q8eXcJ4Hp3JRqT2
EJNi6ZDYI0ZUyeHwrXvt5zV6Dz9+uTtDCqRJefRgJezVhLYnoxW5XHkJ/xnqvKAG
6yxM+JzneNBeMFbM/sNZ2QUx71h8DCuS7LcWCsNkOIpcFaKoiLMRdh4G8tURFkbN
B1lDmf+y19BTVwIsIhmRJqRfOHffKT61qFTuMv305XnVBKxtE1eDCln0KASAv5HZ
je74nKNVc8oEvlwEI2nG5Gmxwf/fOvg1LbcrFw0CCjxuaHP2I2KwzD3naz1feJuS
4xniH80YgrksJi3bB2KuTK6wUumUkyDGjgpP9S7SimoVStqFUdQQlsq/aJvdCvvj
w3smQ7Ki437g4eCmeji30SyxzNgF9sCxv1p0tqVb+fWDjEZC/GrgLhUIg20+ugFK
wgDh7Pav+O8a9ms8WiRTnpMj/jDNSy4FXrC5SRAHTeMvg4OkHF7gTnUDwryzjAtp
3KGcskyfCfUAQjuKZoTBkWuetNMZ6SxO+r79FarAy4wdiiHEWpcRh7HquftKt4Nn
TTIEEyEARpl/dXw5iwk/hOWdsr1nbxlohrPpbJToqZMXJfY6EvkVAKReH/XG5/3E
0RbhkjOB6AgdW7i1JexcKwvasNgWrfpLCCUqnBCKXOmKr/qHJbNRVPwtJu17pMle
u8niWGLOdZ3Y4FLio/ifBk88gWkEArovv1+9MrhJeAoJr49r8GGoA55fwiI8EST4
wP1UZIcs3Xvwd5YgyM/f9O+lpAk3rarbtEpbyBJFqdjcm2y61ndYdyFSqXnMI5tC
HZYZ1XQz87aFCCD1/8vON1fZlAi0Px6Gc5h2JLAbXo1JxGo1DOf/gNG58Lpcthk6
QzIAXfAfrunkQwhD81BV5m26a8APyWQQ2W+4KJjy1UCUutnovwA91CGEIU5KiimV
HXTqIY6ebkA8rBlCRkogf/JplnX5ThnsOR1vLmVY3toLQieYc2CS9yXSc0AoSAyw
xeQCj3Sve1tVLf5jzofGlxOQ4ZGL1VRV6Xp1KpUM8p25N6QQN/p8BpJOSRpoa0eq
VTKA4GADTudsqCnZrWO0N/J5FH7zd+AKmYKlya1iD7sBuWw/60cGy0KOYr/E/T+c
xKuagb9vdtR7meuQTt63ZS7r9p4StLJw8e8mzxspmOIvc23NeILbJP6UDjUA9V0i
rk8tUAPTiR1ubdebgsQKx1EAqH0hokNwXkgDVUj5tUmRYBUIEJoqKUpblRPd5ONn
nMfBxc7Eky3zlZkwCXk9lyY9R6z+P7YP5oMFcDSYtOe53e8eXD1a/8KlHT1dejga
gbBMiYQR1mm/G1Zu7PGwwbkzJYq6cH+dy4T7wJ65LYPR+xUeVHzzhfSpEbeYVvOq
Ft4zphIwtO25zCKrVaz1FkJUsXxU+IiZ0NRNLX9IdnoRHNqoNqCsYZbFA5yHoCvP
lkvulqa31Rgu1PoPMw7gr6jjLnSBU3Q4rbZfOchYbqzqoVdWehcMuew6F/hvR10+
bVMWp5fG4f14vqq1zbDejmreKeIDTO4iJmUlLibqbO2COxf1+hoRbu3/bVzHcy0m
+IPxEhXJFGPhpS1A4H106795OUZ/vbtjVdwpxCxLSHnIaEEUDuulTnQhcEewfz8w
z/NzQ37wTxlMJvEC6CTEdbPdTF51ceybiPcr3i4FhWzu3hiKCNZMxDMbyHRM5H69
PThViteUaIxJfURHN97WI/F+oGBMOzPfpXCfSvhPzsRqbMy5Bf9xwIWclOGepj/K
DMtN4Q17IL+CEin+np/kfmCSvhftTJL7B/4wcv7NcmWgrSrl6Zbf/I9a1Ao708dq
JzvW09QIG4tNtxdRx5kDlRGyI12RDoVSDQAOasOfzjlLwqTU1D9YCOEsGlTNfyGD
B3Ui20TpO3zfFXVHgjfxhYmucovqAwfSJf7jQQ7LB8ngofKuS5zUek+lS69Fav4g
M6E7jCeUW3l21zhRd8o2TWgftirtoCDyBGFHt1F4zITkYIHNRcgfPFGYBgns8EqN
FKi3hT6Pw4v+V3I/p8EjlzxO3nd2z2qDJZLNHdcOsSkUoBB7+IeyrXYTN0BRPgH0
1rtB7hU4/WCdg+GIUcYOTD/veGSgNldr44mgCZSEJXRao/8hy9dDo2t7gUXeXC9O
Votw4E50K4F1U4lveWaq56sSRMs42N/O1JYkk5usdYIlrcneGBxEodjj1It3BWga
Six1654yopwa2Jvk6JKs1DZDDgUQacY/GSFMxVRcXG9mIdDOAwFY3v71wpwMqNRe
e2JVVmZOoCZJSZtuyt6YoKdz2x4vJQJwCcbxidROXw8Evc97DUZVoYPOQZb2lfip
K2PKv6zLpt/0g8/UIMBxabMVsJJG1BznwrzRY8iSuGPTj7Rt0KOD0xnshRTUxLuA
ABH6SwId5jGYbxjNrRqiTWPxXGI+v3/5msn+WYXMZ2s+7n8dpDLG8pE+TX2929Bn
hLT4l4kvdhl6gguHLS7Oi5P8ZUza2tY7xEp9AF+2h0fGCbWGhQZFmEVFNNzTasaR
tPJ+bmhxB3YWwcFbuG1qn6uvYUBmm5oUkO2zbFMYXJoi29xUVPwZfYa92V7qfrmn
dSsMPCL+HyLjutR6jW72BrNJZJo6nMPLefr9LLhaVkic7W9jhqBGK/t81oquQEBW
in9g8YioIS6T7eOFWj5xD/pRmYLY8pqiHOf5NdRQk0BXVkltYK0aeiavbHUiQA3q
fRCK2wLGPS3Ha+zQPeZTTlw38DVry169gPVbWCecsuciwkd5052LrnD3+/5VCSUO
6IqbgyT2Q/RzRB+qk/meMSQcStHeglCNNsr5S5XKn503bVJQvyeaTWdq6bWpJ2PR
8Y+qiM4Jxgt4OjEm+AXraFCf70vEhrx/peqMv8jH+uRal5sstSfdpVRo5LZQXjf4
/BAY1MCCCAZp868+IqdrC7ofjnYcC6mKUlJAaE849rAxPj9SNL4kYJUR+ep9dpt2
8PPSblMAw2mdJaYKw33AIfR6KpG2E/r76DEaF78eworW+Sk5W01dr0OAZu9i1SiY
Zq5EdC0OplxUyRHxD9OMJ6d60+6PoJTVqP5XgI9pfp2MG4EpaBHsYnfyVawLE8mK
j50mQ++YxEqSK+gg3weFUToG5Y4MeElzHZDRYS/OOoRiUkxO+648H2JM9UbqkDoz
FI8MucIlUSJD7juV9NMSdMXGsXTGDk2IFvKIocLeLQWLDqanDmtr1R3Hr1O1Se6v
q/LD0m96BtCXKrYbrQ9SWDMGbSBDVdZqbbntUD6gqS4hmnhN3WbASu0jim9yyBsK
dnLyNIssPbJytMInisOsfUWKvrtGNJoiQIbIhsUcLHX2NRcpdX++J1R1V+XMxiCR
QKzHSRaOY6l1HY1MV/4+Fm39/wze8SPzRFr2/ylQBxoTK2BiypWEiUIhpHSxHbHa
xEAr8Sh9joe6Ewb5Kyj3NzKSQHy0w4O7LITIPM3WAKd0G0LGjKVlcGxr0reiWRfS
RFLd9kSPxekYUWbTWlZ5zngeQPfVB/0gN0UsYAsYNgv0HmxiOjVhC3I/CbCFLF8z
sNyKozcgkzWjlbHpXQ0WF+pA6WC8Q3z6q0Xv/BB+bEUQSbssfq+kOyna0DTNLNSB
PYNQBZKtIzcJPeWNJ5itlqIMAt8Qc9uwa+n0iDeXd/weKjleMQkVLGlrJz5bfo+E
U8POPWVR6dxevcYn7faJObeQvUzruLPgdIkFog1W1FKtrRhgole5a5tskG8l3BAC
DeKBfAHQTa+L3YClfs01gYpSbPFa1Uw/9Yba2QB4hGSpeqmyriIfSCQXYMfvjppa
rXkW2pslGauLimU8Ku5d92CquqaNNGcY1gRglkPAdS9XhVbsSSxiXhM81mtfdayW
wPC7lO34Qz955Q63EPb7ZqvKedSsWwBWBLaer2wYUKC6XqMoNpr1fCt9b95HpKNj
ToA2X/+P3D1l9ZtGzi7AdBwtSp2UVe5JgZb0l/EslDFiWffoiATUGvmI5XAGEwhg
mPnjTXNrbchqWphBrFZFrLWk3NVWlizxbbkO4/X8bJ04dxynR1vmxAz964K814+M
N+NcFjKjDcMts329znwLP+yChzkw5Am888mjfVLixSt0gzuaOb9mMgXEPI4HwqDt
+/5FCRHmFDi5vHGWx4qnMcx/w/NOzP8LpNOBwj2166draiABQaqeGijs0a1PyGn5
0pUKKPmYYhac8AGpXZGqkJaMZqAJRuDZQXdW64EO1hofO3N7NgTGlfhjpTwRKLhg
imQmLWNHrNZo4AdD0l2lsb3sKkxSaA6L7IakiXLhPNPzr6QTvyLq7xJS+hS7siCe
UsvVxEbImslQBJsCUeJbXxVh5W1GzjyIXznYyie8/INuDp8z+omLyoJsgcptQKID
L1pWzhI7xwnXblf6W9w8MXAtf7b84JJ92n3oev3CqmVjjglI98fWQKBMuFDniLwV
0wBkxRO4S0qjNpBGj5INYEk5utnPYSXNf16r+BC5sFS9NeUpGxKcoictpWwn5BSR
KxEc1fg5JUrFNALUGy/YvjO0QSVyHnX8qXVetc0KSjPuG5lDMf6qmCxDnosjhEzR
xVTS/z1ocE1Z/AwLf+ld/NswsPmHLFJWQiNYlwSIowmM+6u7kxRSw+6y0pS3Cz6s
5LZ0fNrxkORUB8FgOAiZoGLAPo2jMU7pi0y/CXbn5wDrFjaOm+6W3QPlDq/uE77F
fhXQMIPfjlPx5zh77mK6f8TFe0OxHZsn4YGpMvHeYAWMHKDY8ZLGsmjxQ79lX4ad
Wi5QveY4kDErxuamD0ECoPb6THHpkg5gbmvvphMPDlDiZ7jhcWk6laNoGgr3wNZ3
807JLkQV/cLEAXogEyhXuFPwMp3dtnqQkTKRaekexlu8Lw5veL+uRJMJRHyvY1hE
Ubi/bPeaYiMoiOqbNGYsPqzd6jDo2bGaEzRLbVq1IZi7mcX8C1ljdbva9t/p3wWV
7Ve3bhuuZ+nzosRbB1l0jce7OtMnpWyDRZFfuVxMMo0pLmxdxWU9MFy1Lvwf9aFb
oK7PT+JAePXpITxMTSjUU2VuBfoiOVP0/pUfo+Gygt0YQv1qY2RxMi407wK7maSv
51663mytKpyu80lD8bmD5N4PXdjOLi6vfoM3diOIMgKmrrzmheGbkEBPyz7gMUu+
7M7gmOx4gMn4za5mq/IyjW9+97FmtDTSUNBzjLdRWbNfUzglrOhf4hMfk8S0pFsi
Cm9a2y6/nlRh1flQN2094sqJkuWrVyAy32C6v5CkRrk1YNzbysDjfGYwl08xait7
TmVe9FngnB68Vh3DzEDUjvI3a86+EuwS0TyhOesc9FDe8ntOqJMHs3+QkVQ78reR
5AfMsSIb13S1cRkRzScrd6UN2PuUvsto/DTa/wki7NJS7pM46dJ2Cd46VI8LmzHZ
PxSXPjuZoUpohJfur2qT6gaBYVrGRCLT0TjGNX+jguj0tRyCNc/XICkpZatRlsF3
Em/pU8HguaLuuPhgKIiEzqp2Re+0RjxfJLt5SFofNtZYbeEU/4BPACwQTCzPEr8c
ZyW9cNfS4KFlVHJcoYtB7WtnROkRH6/ND7DE+YgE17Sv0qKIhSx1qg0ADM+qTRfp
v9t+iivyMw6y5O5yicp1bCq9Gr9x7CxqIefBJDSDlwxF4P3EKo0TISOTXKQotrmC
jCplPfERIlAMEvFLmPBtLFCuuZ5xxWknRod8r4NutfduEH9vYUegQQ4dlg8MI9XJ
PV+6YEjBnSig/WSkluHpuuEwTmuKASeYcYCqXYxyOQrkuTcY+j79TeMVJNb6QOR4
zjlkP1whzJQCf9gnMdZl3ubRFMOhqJQBkUqRUinlkLL+r9k94mzhhJ78OvjzEZgg
pX5nnzf2Sao2P1iSOUb+sWgCYUwkp8tTaimsLN+/8EDTJT/JCu3eh4VmO3zaaetr
ZGhI3fFZ6LTvxyKO66e4d8pY+PjS+r+ubI+r5QpnyDQXDOdxBn1XlPgwzO6/m10G
CYNBPZ5guhrNrRUR5n9QeV3VrVADXAC50/ROe3SMbHjb3Mj/yEMRQR3ncDfbRtZB
Y2M+FphQbC0a3HIfICg+qPYXPbPe8oVd0PV0VVATSyazWz3cG/6UKYrDc78qnrWr
TAzZ8iekAN5CInzt/7hMinLi/GLg1+GwGd5Yxbbx1pWRaY7KkTSoJaD9TngwcG9x
YTLiOGfvJuZjc+sTFhLhmdREasa7ky9KR4QtTKsEyF7mVKAG+WyG9l1D+2+nD0DN
ynuO4gRX0+7EdDhZsiU3RrcIcdApbUPl0KllvZpHoSNYuTUOu4Cwi+HCxl6XE1ST
aBR4XkVYfBALaDc8jzo4200KyJQlcuKAg/vo4BV/aBwEC7II9a+wFI3HXfz+mMqX
Bw8oj6eDNlIG3qMg1EpT/k1saWWte5ELU0AuZ2vjMt1wIf6dmj1CtZBybU6F+jF/
h1JUhOyTtXQaz3xQWywW+/WK+Yp4Fvs/j/lfYuon52qQkCNCzdY7BYUmqRtDF3pW
XwemAq5JPKTuju+mR8k+pvfv8dNl6MzdWK7GokzbPcytjeURGCzGZ09LQQUKGpCb
SAN8F9/ezlcyvGzocYomuK00m7ex8wOrXJpTqnMHK5vAiVRFpxSUbVnuTvK/qlYe
C6cNpfxz0GnD5GfkaT7224PlzHIH3qm87bvgLzy+P3lLZNKo7M1GoWwG12jlESgI
VyiZwR9v9EvBCsaaIBS59PFRoluLLfeWX9VEjAGPscEehykrGAg0JYxSBDCKFGR1
423J4gHGkGBLPYYxHIyEXgMX5b5T4iXsPlOMHnCRP4c7xIlkEbIejtZoJzZQsAGL
RaHug8n9TaixACENL0i1pBTYlE+3tSicfeohBWrkm63mc9F7i4rxjlMMiyBZMlHQ
RlX2VTtGaKycdyxLIr1KMWAitfQf8cj0S5BampsBIdMIwSFxAoEMxgmiQcFFwe4G
E5Z/MEmgNlV0Ig2ENkpUTk5ILi1PLwv/MpeDi+SZz/vwYQkhz547Xi6+PufoZz0u
OmKJr7un1yitHo7fmxA7ZZnt37eOufK9amk3MQzUBxTmClCUIMu+B8inYGoIA4o2
/8LfkJnWCKapT5f0AA8we6+EXXJz09ox9ydkLquKjfVFdl9Y5Xr28xoMEf6GCtti
WcdJiObUXk6rpP8sdGAnPvTY560GNE4uWXHyH2C4pso7PqGrJG8XDEcjSRxa4ujK
HjKmfYJGd9keTZuFz6omutgfKXvni79bAL3678jzem2UOb/dxypF7CL5KZcdHdpr
Q/Na8q+iVcmsBQ3q5/Iz1k1NS2d1IjbCvcuX8ykXo3X1uEq2yrO5jw87BRidDRqG
NgbAwHrWUYGkSr/YX1V7/rIS5jJWdqA8HNzxhrZwK3ckodyJx2tsX0+j95YbIOcQ
qsr3EDpGv6/5BdRyGdCdMaLiG3yJDZiThH8OqlkJAHekYqjixW2NJFo8MGOTCXfe
vOGdxb6Gd0H3rzgQN+0lzYS2HxCOawKUOOaXkGRH6WS7Sbzb5aDTp1k1jkA4Ne6J
9AZ7SkbjgHriFKbhDYZJHvOGOtiygD4aMnhTdt8lMaLGcJVQb5PAy3VTjfbOuvsp
pbV3YwuBVWmM/yM1fIVUb991yLDBHoVRqC80vLb0O7JpU9qeOm0tUFx2moqPPjrI
eaoq2EXfm0ronueSRmNAhRxPxb2AXBX/p5vvoGDsYwPNs+k7KYNoifJQ1eDjbVvQ
pROY1SZ5nBi1jD8Pu5+gPo319zRIYFM09GC4UDIVbY5MueQ1jcvX0ajPGE5V4wT8
e1GoIxAm2k0EnQWqIefrtTs5UKx6+9MXBbMvn17LPO6bYE2ILTnTCxHBtoFCtd78
RX1tqKMdABiJX30jxvZHFhRzmOFkPoauKjYwf8srn9LwEo7ThfjoG8gCISNrCV6L
oTodslxs9Dj7xrzmw/+N0jI3qx8bjAO9oLJa8klb2vHdBoUPtwtks3BMFYJXPNn0
ME2hVRJW0NDgooIu8fueuI1DsJOop0UUqHNQXpi8tTVTrlgZ3ZHQ+z9uUmMJyJVh
8nHDTPDPRNsNWKb0JCFGOmAynjxZVYVjtkKE5/TNtuaFLO3cpO39W7ani6C7Om71
FTlvGn5SAfEeZBJ7PRtrVeqQtShsqRV9mck4iCrr+zI3NHZTSP3eHhXj+7hPZhS/
41b7qnCBo+3+mMllJCrpVKjnT4+SBQ5uzQ5eTT14h781dEUKhNNpFGXHw0FReOv8
x2+WmMYvl0N4HtgD8S01WbD3nEIiEMWGWfNd58yaUTm0ItplYzXgbbtUXGISxVnT
rH7n+8UY8KLiK51LnKNSPMqNy9jwmcSphDhxFNVjcF57YRvzhHk1Rurp1Zmrw05r
GdX6fLDE+UTMnY0luQqb8SMh1Qpj3p+PCwJU6490BsM+w4JqVXzmIvh3S5oo50mx
xvXTOnefRiHuZIE0WLijVlG3UG8rN05XV0HvAz7Ldh68ylEReBtdAmmBehb4c8L4
L7HCf/NqXqpaCrLFreScQQp7x20x0NZB0p/sXIdIuhJ1RIg0r6njSqwTjCX8u1W/
10OHiGgZnJ8+d6RCUkqJ9GFA1IaoJHOpJDWY3pImmtbTpqlriEuvVg7iBhyk4faG
MnAm3FsxhjkpPJzHcQBOmcVpZdPdRzn4HNrcpbbskn66LICeyW3Gb+zciimljmYY
AVav2fURKpOAci7U8MyUTMI2nGxIKa8aYnfh+8w6+1nUB09KRrztzUhLhaZib2Dm
Iawt0sUjud/uQg960Se5QUt+O6p2TK8IbFJDCiILxQJH+pdJQ6KhNAYs2PjB9N9X
YyXP6C1Iyg9GS4KIygvPaYUCKycCPqL3sbdb+Ag3Y658UApJTjdduXxrSInNaD0l
PyFm6zpXsZF0KO8SuMroS5+Ncz6SHvaDHrJ6ssDSet14lzOMlS8SUwSOAL76ylBE
5QGKWdjYctMduqdYj2O212JlQtofZI1TsdowppTQdXIWLqH7qJwbDIipGxQZR/7u
lypXxuynDtKT4fO/d2UweU22t8gv8Ri3LJPYXS2vmohX64atNEDkXhl7BOg6va6F
GAhjpOv1K4RweRWjNxSZx8we+KnqCyC1Zj4RNd7f+SiVpdwnFKJ4XLGtO6hzR9Fm
OfojGfzn1mWL+UzRk0Wan96beqrabklIGVS1BdgefwWPp4XJ/RSh+YZEQxp6ICgm
DiFa3OhiBPbiTJW08ED9E5+0X0/gDJyir4uzLXbW8PsaQ2UXBjgKKxp9svzOD/wn
udx+nV30x/qEvF4jyYZshHHo4aLk+DEZWSeX3VoRgM6AWbQuXBgO2QhD3qZPIje+
CDg1H4cKIXpy4CDskG3XOtRgCeX0RgRjJeGM89oXe5lilO3hU6oTiswbdig0g51j
FJewQzGiiLakxWZ0pbEeB1urXZ8tDUTk4MwMfmfplr4zkmE4/VscqZ+aFXmxFI8I
YubLeqUiTin7Jd2sCfI26phQ6Pk1pRuoeZmvVW+XowN12+ojwkTR2kajA0Rb5+IE
Z0Cm4AhXXsVYL78zwNYAxjEMolhagjkAScLlJY+Qx6NIJRS+nR+irqHGKHeXgnz/
QuU4MMPbat70hbiqW5o3lx59GolTud9Mxh/BC1DGXTxveV31bSnHrtmtZSbZHw0N
tRP2k3oux6bcEOAVrr4w6yGY6qr4Axej7VwJVizwXGT0N4xTV0xFK3lZvt8RSEsr
Ge04inRN5paihI4SmS4RG/PNTfdliT+wej2SAp6hdlYlaFXR6KAW7ffYMQpBmkQg
uS7NrtwGqVHuvKIDeC+qs42h5BkPkD5WfN6ukFz5gHPjPk04AxKlXTvDmWhhsw8C
6Tago1wS25c3U5tqCBryXbWW4lRXWohXFKUiuncG1IHOH1VvsTII9oRJ4Ye59DjM
knIZFAzSSONXQkpDQo0aO+JbcBMIHFrX+kCp1miYWhnRA21+5mIRiKBFovGQzSzh
liycXU1MaiGXo0tFNYGzyKv62axRhbfdTEAum3+bNf55QeomTo9ARx/Lw3cY4t86
gsH0fAY8CVvbh4KOaNpzZC/wcg4pe8+ED6oyKxQuMGoxWY4EoyZFZwoZX2dKpxq4
dxB/jyh0CwvYTHYt5WrnNucuIWmgRiQCXnyKcZaGKchVjbzco/MFslRQn2T51cX4
tJXQpfYlfiDvTeSZ6zwWI8XxvNtaoUqf0EXfxwBa+8nRDVjvRX8cJu7ayLYs3cWJ
Tp9YpDVwQeSF1wW+PdFV6tOR2xtDXkBgtizXn9QdC2vXeOrl3cJ+twVNdeZz2R5k
VTTyMSCtVBuXks7NZ5KlxuXGVjm00wLk2RLCxY6mjiuwHYcEJXvIVu7zIzbr3Lhd
wnLhXMDiSogzrG/nA/qBO08ZMl6eZ7YJ3DFCG9CJif98uTSWCTIBEUh4HUFS0KlU
nhr+8J6tATVQMAgdXJjsDzMtxuoVTokorncwag7u/cbCvyUIHMD2EBFmodo30SiZ
1qJKyWwyt4dBEwRlB3NlZRU/OvlHdtTrb9Q1pfVkwd6d+stpB9zUQdALFZ4gubhb
jNj9ut7RgX+WFd3ylu3OljegTzYMb9GZpQrKvfUAaJuuw0B6u1G8FEF305mDSARh
HDBmutJEAV2epP8OPMrEPpOaQDm5kBqznVgAgvhDTXGPjshXY925pzqqxaZxnAwj
fq4bNU6NixR3MYlUQdmM80HiVbsQ36/l+NnUyj6EbBJCznNBwwcd0iHzppxvtUNJ
5v3Pq/gsEaGryqmNe12LQez1tk7wsSJKdfqqvfPwKWC/tnl1XpkpEoe1Oyiu1Q/X
QQ/xjFdaKuntUjtpX5FoCU7aZlwpQb6QmmeffDm3MqyL6JpUobxnR4gsCFU/OQSI
XmptMCRFMJfrWw0FnQ+pNzSpHkE+N41uTDAfG3epYGCoflDv62Xd676C3nDMMJl9
55dL14fm4KBDPXBPBF11ofePI0BDxu3sUjoOOJ8epNjiVPfCCIBRt1I0aACjVpVy
JITBq3RNB6fKw36E+CnJhvtdHK6oQkZTjxRTt7hlnJj/nbx8kK8t88zVVP4TcRGj
AiJwD4PwCLZQPGwsh+dwHZ8erKFWVnw89kFNqEUVS6CHAo9cWtpt1qrbGFZSYT6z
3JMCBgDqBhoSn2JUL1968lGveeg4E7JEskdGDERa9KdZG3liCq85suNFaVw2O9Z0
e2NncM/ZxTL9bXWtajYvf+JCj9d/QJfnbflXec1YHXuqK5QFkaz0crOMgGLh5Y3n
uwA7RFQwVA+zmokCgtAfzWi1zg9egJSikRWUi0WIZE+ER8rP5eTw6y1PBV7e/7sH
iiD/cEkTdR4SoqGssoAv9mDuLNSlYu0GxJ1WHjrfe+/P9yR81nlGDyzICRJAeW4t
AQe/7kRXnU0o1+vSBHpa4GrXaTjr7TuAR3a41Y80fmgMfRQvmgGIuvc283GmY1ru
2clsM2vGGlxYnX4jssYNqJ17y8aeiwwCLaHXBdQFnNY1B6qxaSM6f/4r32C8/eU/
ILhqqM9jsSvOZGyWoG9pD/MHKuRSuQ6gDzjNy3jaFJnbwJLywz4XDl/PWa60r26N
9syK/soNS3ywV5PUf5JP0sClKwQO7ZRmV+DYx5FyOcqm8iJsPg6ejR6eNeD1M9KL
SdNpyUWheLpCvOL6yMhiZEDPmJik38Z66RbzEaggwSJgE2ZajTA4T/S5UWegzNad
hc9EKTYW/nVS6xiOAl4Kq3e9f8SM6JziHwPj2uMZu9nLEUnRAoeaIG/6iAjc3bB2
L9BEEdVCEhOgB1HeJVDYW107IvcP7iGSEjv0b+Q+iVNBGbfUVepDll4vJuW9rF5c
z+PsBVMx+V/TOd8y4ZNJ8D1oVa+5Pk6WhTDQZ+pTlsN9wLwNXrOmKnT4pnXpzrDX
6PswFf9tEc5Zu13F7TQERQaYf7QzcdHTwRAk+IGZERtSc9C7ZkrnRLnQqhcd3Hrk
LEVy/eoKZI5YQiAdiZE6XzYE9hZtw3OXjL6Q+cYcKe3cWX9/TPARUL5BaN2ptafG
epVpdsFQu7Hnvb56ByZaPKV1rWZ5CvzrCpY/KXx6J1EkXUYmpkvhMOTFSaHET1zK
za0fCtOlMF28zCByBUgi9yB5iwR8n6dRkcZT3J3CKYtcCGw3NazR/KBe6dy3qcZ5
uQpv5BCw+ND33ETTon/8NOpLVFjeYubKmGLyeDrjraF5gPhj40huQw+HaGnQtJNM
zr3vEf4lnkHPWIZU6PvjMYE8j5yQbpafadeDQ0xB6a0WEskFwKPl38oiQSoCH4Qp
EKggDQOk8UNPvr/5s1p+25hslRE5SDtS97dkAyNhGIe1WHPVp8hFrEkMRLkjvU3M
68902ZudWEHEnD1zrQ0yI6boWROWuYPlgeoJwjVqqulndWz6lxw85wThhvWpnNku
l0zHK89OG41fdpxgQo/mD0czNIAOHYcv8auVYsYb000c13A8K7TdeKCxB6loRaYA
Uy8royBiuXNbkOm+gsjXQI187KjYfBuTg4U3O7K9BQF6ZK8r3z1f1hToyVHGo/n9
Iccsgm01G5J0Os2a+x6ZN9gsMRNKF2dj8p4Q5vJRMXxqd+AceO73L5dIIswYY+rv
SoVe0JVCSxtTkR6jFBJzYnI3TFpngzYAmXPcd5eKWeOD2SHYA5SLrQhALP1kABZu
Zm3Bd/8nN2RsR/vMKRBBQu1bbuVaMZRd4qOeAQaACnh6p2mRdLYUw2VDKdGqq7VZ
71063LwtEj32uUVJr+YFMWXObfqvU0LSqULaxhN2QoeuJPTHsAVECP+DJgBqMN/U
kdLsWGI/LgFkHDy4oHqzxtGyO+nPn02cSLG2viwQ0ZcPcYW01HhyZTZSI6GtlrI3
fGJCZgDlpSY44fXt/g2YTKd0OW235iJjPFMl07Gft6md4JGI42eTa9/bXrCQ72SR
OksIWyt3G0h22gMC6I+KBSypWjk7oeydYbbCh9XHb68pMbv2OXZf4keuXTgZJyXb
cjLt6dJ/MYNrLmtGKhVOuaOQDlVQnCc/KlO12KdpWL+PPrfY24aMUoCK4475v+/U
CIkrJK5i6N7BQpmbHgfF+XlNqpLk6nM4vYLVQ779X9txV1N+fnyZ2RE2hDMLVvjk
F5gyh4Ysj2V+V6ZCaUcpe6gds1tHLJBZrtsIuNYZfH7mYo18QnSODMV5Wlu0wJXg
60cnInA2oRBlOEpKQxSrNHdmDlOXvQwny71uBRfnwdjqdbIwsYysdFwbu26PtG+L
wEGjX2dno45iKRwMlqM84rUS/TKJDe2KMbYa6Xydg/UnxyPwjmjuDRl47YzF/pRl
qjPCl8Q57PkfmBR64XFoCKcdr1XStgMZ1edGRMX9D98NTimM/jzW5TlgAgyezDS6
yLJ7Op5T6E8v9psUT2dLtD/1qc9Jx5kPpQbZ/Gpj20rMkmKzahwiWSyaQ4VTv1Uk
/RGGkS7qq/L3HIbdHV8DyGjXpJk0LWDo2hBLMFq+whWnQ+a4UM+2GNxhwpavR3G+
D3pHaiHwpnnAs9H8jsUZbjG1giXitRqqMsunZqzmnIz5EP4UMzfxrc9ksJYuxZTa
Pg3j1fwIsZefYvY4F6FkjkU18vHrNYq/f7aVUg1s6MC6Pm3BVm/r0oRIkUpKWiqF
sjRTPRMx4R7zEaPkKENSmaxWmsXsSsyipzBbYP9O5P0E0C67sQylnr1HtnRgbi5g
nKr/utC+n7JYVWSmAQ0np043Igx57sGK2Ka0XyWtZX8ut4bDnnbTbC7Gr1/vY1mb
Y5gf61bFtbBQMZAYc3IeLmMGvYeEKqO3Wod622/oBhP26HtRULCH39/dVJxjVQCk
TMUEiOKU6zksoSaBdi8VBxKyTqLgy7zitaNROMlhftbv8iHKxgTmwyQnrMqiaFWT
FCCGIh0M3tKDqM35WamokY09KlDr+jfu3pfOtPhvPzk5BdUxdCPfHWgy0zAEyvWL
5aEhdCqq/6LPlPlgepdH89e7q48AtoWKmqgAKxZcR17GfP6jhLZpvGz4KUn1FVvL
x+G8vwVXRPF8X/KmpqqG5pfGwjzThHHsAWDVtD4YG/mj3AY6l7aiz91XTDLgwIVB
HmNKtyewllv8NQxxneGXDg/GZv0xfPt15UzggH97mT1cVLVGvRcceGMwEH1uIqUg
TlBHYLNs+WGrcsHdvJkR5RLvPDOytBWXiGQLHGRwD9ll7VmpM4YVZFq8dQtbf87E
ew9p6+D636Fb4H42OCdIoQkneCRC8rjvkMySx8EvulC5ZZhmBt33abHj8i2dsnu2
0+GmCnkkXHr/bEgOBouOSV55jVu1uj8G7HSCiR7Tiy2nTYxxUA09splxZAKRVRhP
8RYP/6nUQh18FFtKy036pwOIFMMTe2kwC9LdOwWgkXcIyt+CEcFd6fFSPrxkvPDn
KLGycVRSjnlu0ZLYDp7pV2TII01TC/n4Dwd4Wdj4cETBZ7aXihEM6FkUajphIr6R
rMKJc4/4OebyB+65Iz5kLD9qqMxo2/JyeYbqTKH9NMO4ko8waSuvOPpQU1YnDl85
y+yY094uKbLRl9q1fo5roFZQ+35k3QcPR1IzMzOJaT2lwt37whE8TmTIRBeDF2b+
ub41s7gk61UmPhlEFdfpr2yFsSk70Ad0kG7Dw98MYexhMFaPvZTeS++N06BZs21F
hr6BjC/nuj0eG7AaKcpPOHaOEzKJ8xp2fkq4qvUn2jKTeQvPehoQP6RD6Ly2pRHG
ylEgjiSj7rgP0JHm9VhgjLq9m7ShCkG/5D52MiOf7DUAmdcfxzSaxeHt/701xPlQ
tHf/qOKUn+kkF5oTWL7MxbxAAXmh5xRyWQp66tEb3B+tSJJeZxgxjbR89gUI5pHO
5qk+ji0uca7Lt2sIzNayKjJfhT3gObsko9piShHPcoFEZ9942Bbgo225qQRytmCV
PrSRP2wKhETEaYAe34qpftczfVMZ5RbPg9t1DL13WRI3ZYd8Qto6rQbdy1QglYPT
sFTbQtiONGOUn5GY9H623xjpXHhjOv1X2swwzuMCqyho1qq7rSI4HWzGB7UemhP5
XVK5ccJaVoiLciSW0DzuDA+M5eXTgXq4WtlQQHkOmprw6aB8+JuivqIUIhzrexJQ
sD7mgbrVtN1UnvrR4/LmI++emQ53xLQfL/0HSQwOPeUS9rOZR4W45wZxJo+6rSZs
PGxxN55Q2OW5XM2OeDdrOTYp4LMxr6S0iMG8XEtyS7Nqe1T7SUtnxUCHObaTil3m
w4AdzxhNIpAmgcZDaxGGbMCtp8n/7bhHCpeN3j2ypeo0dvyQJskBt49gS1wMouSe
ia7YFppCEDA+dQRS6nMVvLI6ncLh526kljx8fXhv9WAY9cmu308O5yB6WijYAdlk
m1MQAvW8wZBeFt2Ed8jrqfYU2obgRrjGFVZUcgiV+Z7lQrZrax4xWp8JF7lDKNvj
joejamWGHqSCHBgvzaet58+0dQEYICb2HhIy7RxxnaPIS/4kQxQJ3VAi3ZmBngGW
Y+K0GJFrC91PdWOgKAfCISSSwjThQ7SeA9EOwOP+X0D+tlyQis+kZ6vWNWdeeItB
LoMI3yRWZVmH198eFCw7tNeiml9aFBueoIut1vIPKgN+vVvGPIiLj2XQ2bvo42Sr
P64D3ku7tgjx72gSxavh9ItYTfESO0zknb78/0AL7cSBaiKijSytQri/YaT752bR
16CExuKlae2RsaC+xsIalkrvSBToP/FxhotL7eitKf3wglxJX2ZcUnS9Vtbtd5C4
Sg4aUuMaq+4u9Yl2R0h0L+/x9ITXzbw/W99a+MkGrveCpEZ6AirAf4OSy+3VsXF3
imU+QhQxTcT4vzUzsmXKWazDxW3UOsGAzRcfJVUqhstF3AkfGg+iOUgV8Yzkker7
FsrC07c1OPnOR+4XJ4ySmn/WzfdWmeiVIDMptntzj+Q2oN0V4IEWeXm34oVl4+hM
jfD2+Q2KIP21XtxiObQjR+lryAy5Q4X2wmcBjwgFx7D03oLQsvKW5w48ggi4esLD
z9AXM8SPMopEQGncxzS98aGwjgjKMAm4la9NXRUhu6acsIOG2oI/yK9XAarrKEbL
YRaBbCf3qmHJk+QYfj2IBeSefbHlAqMgM+6uVIyMYcrrw5+xaXsg+C3AI/IEOQ63
gSn/WWsuk/t8TKwKCiT90RWkia2fAM/LX2TSePN2v00y5JVIh/TTj/PUPlvDp/Sm
gfCYVWYFWSaeS7a/VZLQ2/QS++rh6U6+82z2LzhrXUe3ctEhvo0hAHRdDodq1T4c
6Fg3dBF+9LkU4tXHEKWy/ZtkLfvnZSI4cFanuBBILASPdbuJi1fEwhfaDqnv/5C+
dTQsfkobfUqUSHeyqCCaYMJOR3Bb+CYRb6esvrr6h28F899NXe/p7yZrH7wIdaRK
6RbC1pGmBYvKOTr3OaJB19KkK9NnXULmH29DFl5PL8FEEIxqOWFreA6iybTkAiKx
a2x0Esqh1X3ZHimFw+RSgawt24NFepFcE76x8duZgPNPW5NBOpDbg3uKZgwPx02S
wBadK+04mbu6sqI8+5N2o8qZcQ1ifdJgULCwa9xZhhiLSxoAaeek741tA3GN8ooq
i0owOhPYHzzqKuCbpmgso4mJHsMFpmqdXOt1W9MBzPj8CVH+X6bh72rWiyP4Oe9n
I7kK1Y8a+a7J/5twE1PQPcyogUCUdpN6h4/+LtoR2iq4B1LNmHVtvcvnK+IFxKJm
dBD0UOpiPMsFkD+xgFjCxhner+wT3ctW2ON4ApDwqw72VQYFtxNk2bUNYvBmUQen
L3SHVkJ9MRsSYyeQVMIiAOfnBwUNg3n1E7nkj6qmN4Yd6lGjpQC8aQeaAew8P2Gi
HB/UA+iAmNReVs0INdQBGLo+XLgFpI0jhJdht1/vwN+Aho/IKthHNBVsPvtGQSZh
47scZhpfJ+ATj+Mmz1PWeJNAbZcG+MYHU5LtRIk0Q4C0pn4J3CWWZI3s1uek2+dr
l00fUSlTDTt5at8f8Orsa3hPphf4hg+Ne6vPqdNg9HgUgV5Du0ig0I31dbopw18L
7oLVIy0R6hQUXCMpmeLR7ALP6sMcMPP6VOGV4te0pqirj2OIWM0Pcr9JNL+VSJlm
KA5LPSOyivfEl+wRU2z3Ke+kS6qYX10Ke8BmfpScR5m91AVZRxXVfgDN21ifUDK/
gczMp+qFSX5c/rKVC3sjFafLDa8wFcILGowWPZSmKxA4feSAzZ/blt3yHJ1pMSVx
g0ZjAMJANTfC4enW2b4ufiwPrLbkFA+/BKxTmTsizGbEPt1F3x3RFPKi1sy7pmBY
L1bvdGulkegjO8g2J29WQzlYTPcEnQ1HPNLZ1H87ozDfhaFEVaih+/GuOE4rCVUU
SjL4VeKgU1sfugMKubdArnyoq+csGG2U9cfsHgDd5GDREkSAcUxLBS0+fGtQb1VG
2j95BPKMnup8RSuk22x0IWShUrX7oqmUoCj8EY0wnmtdoDkc5/y4rQh1nxm6YUc1
Q90NtvRk6tY84VhLGfqRuPf6nXQlLwrBhmsdAgT5WDXM2DD4f53i1SA48e8OxfSc
Ctug6wsdY+p2v8DumZ1N16LqVeOS8Zuwy3vHCXOqy8uawZbykJmyFgDxb969533N
GkUOg3uopssu3YJpuMDLjmUkghdSMz+1BUjkcPW3DQcgnkiItOZV06LTlP3mlQft
f+ZiH/q2bzhTDvbPMrw6PwEBPDF8xvTu8UmE6WXaipGYI5XE4DP68ZooJDaTaPVV
yJj6FXoDSGhy4BR93buS3KtYh2NBxp8GcKf4sp4WjBlT37xlw5urmS1eRQi5PyD+
hjTilK/0DcbeKFFDi9ZnH9mAAuJmMWAeLgtdLXeDC/yjnyAofr/ynE7gN4KFcQx5
pA1QEMLO3s844T4CSkgcsJJ0yo8+okrUaroM00OpruhQHlFSLsfofrUDh/ZP0uNI
4n694oDUAvFV9DJYxxzL2MQURY771B02SfAxr0vL59ivLIihO1P4jsh2ui/AoFju
CArrUyaDUV8Pp1Fc/u9BZqCwY8KvHE+Tw+yP28/nKHXCQ5X50aFSa5lQSWpbqoev
w0IPINcevXh2+cPXSLdJg0KGJ8Vszqnw3DfY0soCZ7+EUbIyXV16CLZa0tVQsU4+
CJDJb70y2avhgwTp2ACKlY3wMEO1lNBtbO08SXB0rqiZs8y8haaP1/NwIKpD9rPF
BvzY1MQkEJKIam7m169QEghTOqXEIkdV9EVnDzashKiU/U78Xw9KWyDFo6lzLZ+D
sINzXIZRcsZLms7DICCmwyBbcYEpq5YTZCpW+LI2VHjs0W9hB/Ixvn3IK9BRCmEk
oR4mVBr8IsGOaxd0GgiTxfeISyr0koZEu4RETHTc176WMiiyBRnRRshczjIjFIvj
KLUJ8cxNbBpA3/xRVLbANCJHq0zpSkW7lSE9QrL0kHnjyofzt2wBPA6OC1VW34Wd
WagGBzvrNGIVWhg7FsHsBoHA/tGCx3PvCmtDYzgiA80vBJrHSNgYn4c81wmBmR9b
/md5nSoTZUvaU4ppbOaLb/5LN0UaUVX7QpmrzDAog2ZMNisOI7dOiMF4RR0wQ5Xq
Yemm++iQaKcczW0n7EtY8lAqVFAcapAWbaf77NGtDrQfDIs8i9djgswITRQhIzeB
hnBh7w+FOQ0FiKIlZMCmJOiHJRVDBdfGWkqs46P8LDQxAhU7FFv+3I//ukudZ15r
fX6UdFiwnzQCj9uB9O0fry+oZtFnXM2jG6PwVr+nm3Rnu/UflqSH+rBdR8vxseQd
81Ki9Jpn3pQeZyxls1+BaSgxKVO4Q2s6bykQVjkLDp64Vwg73RX7dVdk40bdjmiD
LB99bZjN2aSd6sKRBmeqORtp6lFu7ET0VPueLw6+W51olhuoMcGlpEslJveRMWC1
BBX0TnOGlVD7GP2w1Co5YfMXCw7hAV0N/7GTjzzs1RKnNSl0lm1fBFvp8vf6iy/N
ckB/otojGqXDCpULInOtgVMokdo47YmCeY1sl1OPN8+RWNjvG59vShN6Rh+j+Dts
/ZYZbBFjy4Sw1ryg/qfBFIT6Q+xrnoryUVnQJ6nRHk0jKV9cTY5CHAFHL+luKJ/o
zDXFLszCcgrwLqhSHlt4NCRCOuK+Ke2q2nEPZmk5YMw6nn2OW8i1idnaXDspnYWy
9fnqOKyN7+HD1UHwXEUh77ucyuB+MFNnNtBxk5Xo/+iFAXVR8Ucl6ziYcndHl/gw
Bs16y+vdFXg8LNy+fKY+haxgbN6sn7tSd2cZuaoIYLrLuYX8cvbl5igvvAKrUlEt
XljGRxmCtmdGr0VxSEyzpJiSCLh6ZPciIaqdnWI9593g3y9E+0oa3J03vFrk1dZC
HJHio81vYMm4e2lUauzWsqAf+jYfanbFxz1yJ7gPfckmn8Zq7o4H9JdU0uBQm5n8
qWpaDbFSXN0aoGGvVpngy8uo3+6a3BcNnnbsuenEAzVyC3gMl+FPpR5TtgQeTFdJ
33V2rw775GLoIEktM8rL9cMgJRJXOwzlxNm3hNxqh4yIK2dqgyZJ9bMfcRUViAXP
1RYNejpdBhszDKy0L3G82DzamuhuyKu6mr5Bq+8i3Ou6+Cz3v7bMC6I7Cj2DTCxm
PCmw8qTSUB1NisVE0U18gFAJqfzQ1Cpz5ds3/zCrC4BCa4tB7NH2lwHWPvHmzuyl
8lkcCPxZ05aSgDn6tXeYuENOG+JOFk0taFbcpaIQ7HlrH6Asp+rT98qv6MmVtPFG
eIGuEQx4q0XUXksWZ+8lnRBHqrWE0E/rLwhSkU4jGivOPgbAScGsrowOti8bx3Fr
6UdRin0NU5haVmQjiSjytvhJ1tgEf3aReM3CqhLb4KqGg5ShaXBvsB7g+uAZTAN/
ct3MiVaVEww4P217JvdnxEUL5NPtTWiF0AKDj8oOKjYF0eaVoUjwM+gOZrMGPXeT
zFq4yRfzZQOj650+zowuQWtti9n3K0Qg+Byu+0gYZ/r2a6x4a4prBc1pQlkWvVBz
dbJyA7K9mScJHNuWpMexPaEPpSrvH7zz4iap4R/eA3L7vmpK8gXyf+322YjyRnGV
YHVKDRzppu706tS5j2QWpr0BnRUyyzlEOtZld94mSQLPBCI+s96wNGMe+nIUZHw0
98HbqB6Uf0HZhV6uKxVuAauHaynRneNQXx40Gjx+q6/G7JGKHTpEHilnc66k5HaA
e22t5a6erIUrsFxOmF7jiefQ+yxYOc+D8gpOfLsfBwRmU/4y8S8WT6CM0KkmSkV8
2h5HaWJbFmwmEJFsUnBXvHpcSKiupCMljJQZ195dlC9xeOqYBafL23p2++3wHY8z
nfa9bDctRPXFGI8EmIE/GaXBXR/njiGV0Gp8keh72ArvTRMTn5H5K/SfbUnC1V0D
JVPlxPYcIE27lkzEWOVjFUfu45gzD5IqTfUHyhbhc1PptHf7gGgkMrzQX+BRqSoE
fldEFXaquUDlaXvJmF4TBkPhbThyreE6YJ6F4Enj0/zHuEFRtLbpHq73sCGRTyUB
IWvSu22CufiNZles6Vr6rfxvIhT56FeIt96Th2g6hFpeCSsUpUjFquoNRv8jZmcF
D1m4XElnuGz7tb9vPQ/7ABbO0BP7anv/BshLX6I0IqdfKtYHYMLBD3OLu/Z/lySZ
AuU7LAETlglLhBKh7BLmgTxXJl+Wp1/F0xbSJnoXIvfLetpnf26yVWCA4gtbvcwu
eXR4X9EJquckP2vMUsS9JVSkCRm+kSOA7kPJCNAV9HpBvrDJZ5odz+foAtYZxPYK
dpb399ESD+yfvAmSasedJTSYpGSbDXnBPuAimbvRKARxEmexkIMHNPfWcED1MaLe
FeC55tjqEu4OSigDf4DIyN3N5rYZAxnUGvn7Ocf31hfJHVnHkagqIK93ceEdyC1+
LSgIMD0BmUmM4HE/4Iareg2BXbA4d+yKt8qnkllP/FyZhKj3NYAzoS29FgvLcCQO
/FJbSHi/297fHsDa5fCj64KuTajQGoHr659VaKCOTiaHpCMNFYUGULO3B3JrRYWL
5ad8QWquusciU3QmIfcdv63GMsh7T7yPPYoexFYqya3CVvY/qejfPLHtJ6WZ435+
VQnslZ3cxURNQ6+onegf/lamFi1raJ9Cd/PD++C6aFk5BDGxhGp43+xNjln0DHQH
ln3YBbk1s7DXX+w56UNV4zfRYKskNfaSbq7aXPiI1c6wAXhkS7Ubat/PGTVjxsHX
`pragma protect end_protected

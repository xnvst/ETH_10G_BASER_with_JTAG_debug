// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
S2aNLx8na9Wq38C5AFGvg9cBYAj4yIPaQUEMW0nGKzQEfXkNoHSEtihO0mWySVJWwn+2lE0tk7p7
ff4aosT3d3AQUuDazSE1Y89WVHauOwgNuZeJbqD2CjgWUue8ON65gnsgl7enEnziRGHlxltUqMuB
sOehwpSSSpXgmF7jK4VW74h2B6Y0mRe0nsIglcQn0WsFSzGecdQyJ/4O0/RSwrkUVnYGFYlz8MnS
m4cuCAIXS7hGWnqe4Cnvc63Hil2M9cy3i0tLz2vcDSVTb9gUXjldZxvV37ZtwyCbpl+YPs/cWna0
SwTWaFrFwVOVN88yZC7Qkix4iIbghvd002Krkw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
hDYcB/Kwi7pCN2Lp5cLROZffCJVNw+hP73fp85q3oBX6LAKbb4+BAp7dnsRqPzG8lu33r5s+rx3C
5DJTQOwmwWxdIL1C29K+qi6LYnNDqBr+QcvKFdVFq55kK0Yhadb88GvesJZjobHpUI9n51KCcdmy
OExB+thtV4eB7yVUoSYK8nlrA6DBQ5K8JQ8wfIcYYc4WtrxuKd2NfPD7cZA4dAucWNV9IKUdndMC
lJxE63lZgLo8OjSwpGGOHRu9QfeFW7Slsg5nlFA1X5XQVgUJ2EP1aCwRqJjeZRiHVAotK5gCUdS6
YlhtkzdvGC91zWhGbF88HsuyyUqnB16wn/yFui+k68r95eqI1rhI4GImmFuy8WwXKqM+cB8wzyYh
gilCQEkQY2bA/4lknwSdXVmyxxsdzCiDvgwNEcr5FQykyKmLtnCOtZ6PN2Pu4wNtKLO5X8JgNtz0
l12phwtkf64UCp1o3JA6A+J8kOAK5lbqyEwpWFCVTBYsDz1btOFDGL2JBGqsLUEMWEgvJDU1qe/+
gHIFzLC9SAVTYOPcNsALFr2DNx6S54M5mJiXxBJbHzvorLWUNkfAwV6MzwIvrmTp+5bBOtYk1yIo
Q91jg34J+G1nsvf8HDVEdKbdfnCJ/4DNguqP86rpUTt0HuoF/8n4BJnBA9yMG5IG7vc6rpSA6mDs
Os887cT/+oP1Fk5PrVN63dD7GfDNWVET51Vw0edRupRPpXM98Uq9Hx5HQHtSXskjtKJIkEthnYEK
WnpHlzOUgYAX9YddKE1D2zb8q3TuXKFo83ynSeXHFfUtBJuTQXQsFwB6EOWV5jwo3Zwc3xQuAtCn
4iYfEKup2r9c+zoB9tlewZ/Ic7Z6ocZmDDpydtiZWe6FUjk21hzPKiSiLo8f+h2iof4g0GXjSVfs
kK4S1qSkda5pZRjmbUmvrDFdhfgdSgA9GlaHoj0B3z4B1XG6cRVDDu87G3f0BSXUrfnK55esa1Pz
ZSBm8SZhBPRbl6d1xOsTyfM46xITRnPph1tmVDmofJCZ5bUg0PzYmLXOsYChQ6WOoOR95WZ33vAe
9htRLhAyxm2dq+Qu5ERL3NaEjkWAdiqttn1zbIjTU+NaatgZkXGDA+l3KkBYSmF2K/m9L6jH5QvV
dIl6x2vO9PaxJXmbUaL96KDZQwJFYVr5raf8JZtFYxls98oMpnKUxmvyl1Lio8n0JoRMxJiDW9ZN
zNZunXuatf8WFcLyhjDp/2kyjH2uOdVoIZAiHrvAWvSf36H74rl7g9HfrF/vvX3vid5s96rp320O
dM2A1Bqhg0OvYSIPw4tDNbjJd++T5ePxzYFaluTsdruiaVj7f7NA2L+IDAb21Ga2rGNUSHSAVCFz
P1oMXubKgYJf7lsZGW/J7C96PFtRIbUs/yDPh72zGVNqtcp1sFrnVzJkFn7QA+TOx0Xi89mTBJJ2
QTW8jDrjrcvib7Aoh1DBztNJvarA3HL0bbd5Oia4JoWM4W1MOcEcO9lek79cO5CDbnAVEehT8LcT
8eNCu6vo0VvMVt+6RhNoEClyHDvrD8oJUBPeOeTd90ViLCbL3lYd4kwp2RV1AfQqoU/iKWC7bgFS
pVPA827AwU068mpBJrYkThPSMAw+4Ovk4c9i0sUA+Pt0nwmcX1GJx+zOHv3tf5JEk0U/eNL9vTq4
40QJxeMDIUaLPZ3sJnkGuVLwBqeiojJi/MbJO6HUpt+aUPYv+DMqVY7xkHdqb1QMALmKEre09aSU
p87rL7KPGJzx54ZuRlRFoW/dfF2UDEEYVZEPwVQc+IzhOhL+2XHmDT7a6QONZLCqv8bZlqV6m7vC
Rl0hPnKdPbZcvzp2OGq5JywsAVdF4BD8QVc0SOAb9X8SVtAquiGuGu4LpROWwE16dG3Dv1/Y7nuS
rZ5UXwO+UTDqwfDUfB6iOKAFAVHqs4S/o1ZbaCkPAcq5SjD3boNsTfmMRwrxsxoLeOcA4eODCOrR
BVqfCGbOLRswb6xro5XnrlmCf0q3nJIGilQVbGyBUBkuWJFVyGXAHwqEPdORT7W43CnWSmj20ECh
Z4GrjjSLQT+mOnqy5WNpFO8IYd/hQ1m+OyYXgFBlWdBdlmsJjVsstF0Ygd0uokMgO/m02OhGedX8
eLoeiOvXnZXJOq9dRw4nL6f0ESmao2jh28dXJOKPGw4eDZV9AIzsbj7Ffq1+RndR0sy1LxofYYWX
6rLCV8seHCMeRZGJ8Ubk6m7Sw+iTf3UxItpSvigoGEBe8ELuVHbkteAOEIDCYXE6kkCGnzNFuY7C
1u97YpnB3ccRXLU7ohs0OpZyTxTPwl8znShj2GgVGfPfDR9j0idsFMsAhxFA3qZ+8KRL0HUKsb4M
Hzor13e983vQHrwemjS2ouILz1wv/DQpJ0V7US6BILq2nypPG7zQ6+g8jWiCbUFxMsGZr/3pQaCn
CYiHVGw1ndyE3FAOwT5tFjrsICZEiBamv/XUljG0mm6UL7WMVqhIV04UbtC3SVFKqWevqtJ3K3nX
5wguHRNsfk1D1zO9Cxub102ZRp+VzFDNFxkcUHDtUErBPuszjBJ9Td0I+b7cMsnuKbaBbztpz+Zx
OHSD1U8/c7h5nEZ73vDBt5ZKJ+e2Jrlhqts21MW51cKGt+yN7pAzeVASSfD3ul325u5uQUe8vQpZ
rRq9XFRqBByCCu2ml8JScfRVJg/wU4HFVJMnyJMliXyZo/trMFOGROXqZHbRXbaQp6QK08NKlqGD
IJNikF2GCrV/Ed9xzDcX9ADxkXzCbQzDur2kwSb4HtNVoeefZ2w95ue+Hr9MkoWdz9cmSlS6YOVx
ptD4bEC8FpzWYn6n2OtVSYNZ4Dw1OJdI4/NTqvsv0JI0LPeZcjFVt2oOvOa31IC/pfJjKsnPMk0P
TSsb40B3O7J/euTZCdOcPrxJMDybtPZkIfq/MuU+UCIiOeta4FaGGdx0uI3Z/Y+1rfRN2bk2rmjz
7iyOG0BjoYyjukW/y18oNQkRCGYDzTD16bQmwcZpo6OYZ6TCKVGcJJqJhIQKCo86/CCNCHQxN1Ng
7QDdNEJBsdEDRW77U2cWdptcZwwLI7eOexMM8ZB8Wvnj1ncijkMl4FqGZ3gBXoiVCBWOGO+tvXmE
B/8FtwPfIG4ahucmjqO+a87sZQ43cf2r6g7CyS/dRrpyBAyVodq5sLYVVHhCm/whLpiRycO2ECze
+Aj3USduVF6T6TXBVw2RsEefRChALhfz8x5NxT1Uk0bdTo4RaGIWk6YvCTUEISh4DFSCsbcLbsXo
4pjrFukMqpHELhfzfQKLHM4ZiOQQgUwt3l0DPkxu/d1Kx2RswfNvyEYQlFc2PpfykaaMhixFzeVc
kYAAWUXhuTaq2cKmMuo4sDSdUgn56+rvfRaO+lYU9XjAup17ZqMC7Z2L+ad8JKYEi9y6ePNruCs4
cbZSpCftbl7pqhW9GZkFC/4Eikf+9Q52b2uXRHGLyNgl4N2LOlOnNBPgQSUcccDDWAgw033z/C0D
HPU1FmZ7aNxUAHdkevBJ7bcWng/f7w0GwtFK7MltTfg54ZjOG/FJbpr0oFlxKv/Szeg+VHdHfZhl
mBFe/4eFiWLYEMr9rIWHChovsEPpmSA+OjQZrXoEah3PRHd99e2ocmzcywcr1nzmR3W7ScOYVULn
6YZwQQouVI3wyWt7g8qgEPl6kgSpG7jYoyjgYvr1p1OVl/OlNJykRs40zYyjVFhNGhXtO6Dvad0V
HRWAKiA+AHw+7cXJmuSnmII6RNuipdEZnc/JtTDhI5KreS/ndXUP9AEIrYUKnuuY9N4h/iFgMLhC
sTS2Q7xX/le2jrX3xKZjH+5MNG1V86RGGFF89pWPwCFT4pELRjElwbGkVbcLGgElP75jgADlhMNn
lax882GtQBNw4DUiB8R7rVSrRQFXePtYbEgME/2ItZrh0CE8NxO5TuxqMpYJIHtG5VT4uWueHblf
0afAn+jeMTjVYVPKOSZuByIxpn9oX1IDycx7ojWgUTnMAuz47Yg8+QPYBtRwi08bYaOx+IPykpnL
ymGjqoe1A1+Xu1TtZ2YZzd3yq8uIYTNKdVRxeS5PaL8VVYMjG1qQTIPM8r1ZvdBxUBsoN+uPXOJC
AyCMoAwWblCVA3GNmcdT7ADXXDQw0g24QxLNsqfi7aGQFsc+Zu6CbHwfuFu7hjWLVsl8EIsnpqr6
/dV4VAMmHWZXu9XYr7K+sPlQH7I+qWeQ6hStl1ClFUx2bnjwzS+OruOPZ1C+3l50FkXhDLqyep8C
fri16d+sVulzTHbGm/NXV77atz2hIyXqYv/FffYNwCph/D+fN9bkg9EC/iHvCPlguoIn57DxrZ7I
xb4fvzRPHlN6C3TfGMWUnMisfBcqvkB+ylzlf/ARUWtzuUZsQa3mdpqWK8FyNlYCrv4tWm7IcpB4
RYwsHH5vBmoGNMsKxQcwkjmxundr/SAz3fVBAB+4cdd0FNBtNaK8PyZ80z3PpRY18vTL2xHHzrjX
Aj7xUy4MTUGVDgyHiBoHwmPopxDOd0sNLswXc11/inxRrrr9g9l0yb8KrAfUvycDUs5DtcFkdYu7
wAkr4WeV0YpvdFgXJ49FlgDP0p1c9jxi4jWpEkgyaeoIb7BmGCk/174mY1otK4EBj3XO2Z/dkgY4
yLZb6B9ygLXwqnn4chSvopjzfVxlKHuTjGzFNFqQIG9N7vDJ+J7ngIeTLvSV9N7lHwmupuDqf1d4
UqldS2Mhh92KWNOpgQnGsJ5Df7AZhbnBrDhyhfIAN4TOGMO3WKsMNCs9WEEN6rJs9BWxKm/FSuid
wTGpscd0h17jeKKzpDu8Xhru0eRwEu23BwTDAF54XIQo+0sQuAmvsal80zYn6QE0+erEK/b0vEQp
ZDqEy52qxld/61vSANK0N7hJwnh9XAvFFE2nw0hUEQNpeYVhahNJIISNFghShpmsHEC+udKp5dsH
3p07hsfEIBBZVoCHq7oP2tlINUzwW2dGcCtEJdVeyQdrhRYzbJxYUQPmrXOQhnLjvhQa8qVeD+Wt
izvxwQxeHn43HibTIFl8bXbyLVNEHolzvNzYnkbUkj8uuoeEQiCDYHku1JbxMeyRp/Us8KlDbSVq
vmFdd6fgZRNX3W9MNbgVcSNqBeJf2OGgxOZnQwH2FIymBEUi0mka5Hrk83vi4kk/AOf/E/j26kDi
x7Tw/dXcNzsXQ1F6yKy3ksf4i8a65lhL8myFOQQZWyCau8qr/hKz0CdoOmw+TX5o4/lgMsfw1jIF
G6yUCytX5vE5TIkKxJwQJI0b4AUxuMBYZFCEyEyP6IsymavhzbCkNBJkLJMn+lREgZD4qMLuXdWj
dS69L0PIAE/wkFKfCEc3JwC6NKAnLanbCc4dmXMBHglV4HVltNl96KeNZB3BN73+nokR4luSQTEu
mvLrNcrMj7DqpBBGYp9OMbw6wbwNyofcs47X8md9Ip9oXZIoCYLtnZOHGV//OTTut4tsmY59Fmup
CvTlEZoDNn9fmhgsBGItJ4mzBfMiUxCqnoRrVkOml7H9LWCucjOUpDFXVi4KAymHZlWciIosMEpe
paefrq71Q60aXBY9M5EGB2aSmcIc+WGOuJNhUGzQRiL+d+Pa3aEqnEqLbuc2yqUrVXxEpgOV+c43
6FdAZpvbsPx66wrMJ77RtGFfAxTjDZYb0aJCDbeO86rwm/iVilrv0QEvFm4+i9B4D75sRDI9ytl/
WOD3ilghTy46n372XBxa1qrMICh5orM5d7fSYIL6eNJZntYrttb0bfmT5+R1wivA/faxTkilDM89
rII+3mN+QwyJWpsGgHJgmrxTyYPPk5giBHwm1CM8K1+bqOsvIZjKWwAVDr68uu3i8JwR5C+t1sbu
+F8Vx5KYelaV2EJAEASFykGikv+8aVl89tmhSlrmJ4nWH8FXNV5Dr90tEsWW3vKCaeq+NHfaGBp6
QTGC/2bQjKjZbAaX/XfNDRDDbWUeH+NGjxsTdO3vqp2OD6kgRsG0QK1gxIR+amfxcku/3Yxm9m//
pwBS+zuIBE72e5Cj3VIOq+Of+bERWoqbBS5VqY/m4nqJ8D3kNaJOkXrI2Icn6i4X9xazAFxMeKH6
NRUHSX0qqErBb0GuXLKDSoq6vIcYVLeA+t1xU4xp9xeU+A0eS9Hoo51Vrl46qx4ZTQv/DPmTEQr7
4DF2YqL4He2lHAuPBWs70VtxWlgxmo5LaXkJ3NghIOKE6YjL3WD8JimFNXNuo64IuiMTYE2VpF29
/Zr2GGkdtm3zDvoib6BcAuK/bZ/jJm3C3N/xJR1m/7SMVhvl8+sSKbQlJAa814B9ScTF7FIDKyAV
uCdcWlweofdMrP3Rk4od0lkXcOHE5XJGnOjJ1OwVMwESyFsRtsTZY34mm7YaqjwOh3G1LSZ40uJV
HdDQI5Ktq5EVWuUEq/7YiNenqYe9FIYG0cT3Nk656y1Vo14tmY7YgX+fU85J584jhYDf7YScqYKW
enKabFisc1R2y8raFLDvHRMuUNFpfQYDNwVXzPaeRUgGXK3nvpBmQIQjEYo/ycvZakFZh8gtgNkg
iMU+vpH9rs6BEmbskcRDor+Sc1bOkG5sITiTH/yh4qKtRFbtz0iYR3TdKo8TrGcN9QaoFjCBMi7h
WnSbvvEiLrBaQnNjD5l7aCTdHSp9u61EAckGeFR4CKS0ZySlIRc971yexLN3349Bba5I4mOZydVq
xyuJ52jNLUPVesEny0qOuHcbNeKZ8ubgsMbwV+CRK+yOZXCKYDrvBUv5ido2/RmrilujBL1daRoA
G9YpfO4YIWW5ALMQnlLx5eiEvRCHCvSSnA/9PQdvgciCExjw/glH0bIbJqAGIAHypUdv9tQRfZqO
nzE4/c3WCNBwtPod4C5iCG+FtoPpfAgdcIYv47r6wt4j6s6CXW34IRCbkllH/BJ03CltOubK2fOp
umwZN50X/YcfE5BLZS+UnAJBei22qqd6XlJZfyjBeY6XA5uOrgVw2RWPPDMlsI0KdERWvb2FvUwv
1FtgxTC3vdB0r2dv/15dA7bE51yQOZwm+pPiHItLDhRSSTe1cQvu1RlVVbMEcdOl7E12Fm4GVeJ2
+5qaPIBcj9AWWMX1TjbpNHypMUKM5sF7PHfoGM3tPy0H4IIqMljuX7xn2mlFIrYatHbRiZDu37V/
CcZ7QanzcJDD8ThaculYMJWxT4A0nm/A8e+CvHRq78vMTW0zkz6m/zEqdKCLWXiIe/sZmzikyaJg
FggN0tSeYTJxlhRdlED2ULbNX5ujTQwi6HuSOJzS/8FuY11O3UjdHaDhhMIbnFSzP6BTez13dxPe
m49KFwwIoMqXrYh11XFy3P1t0iVVRiSMQ+sExvtXpC+eli1dxeeFCkVOKuzf/gP9IpJIzoz3zydH
Tg3nYztO4o5N9Z1HwDk6NQDiShxo3lYnxVFw/MUbItPpXzyh4inwrniV0RYU7Egaau2ByvGiguHW
jF0UdpbbiUIRb9zQLzFVdMHjJlo3DkP327Xo9A89K86gMGLUGCTNgukCyalaNUlxHnFk76a5A3DQ
3otOyT0DB/Aodz0qFAsQQyJXt4eCbKOpS6ez2Ax2rxy1X37nxNHv94GPsTy4IxarJEUonb5siRz3
iP2FD5VUJG7CGpSrayglzO7cs0qhH0Th+b0fYr5B3Xs2yWz1ZG34Rfwptg7lvKXIERXE8j/XZTJh
5q9US01qpDasMxZVmvV4/sQKWgV9DJ7iTCuIPPlra3HPWL/wboIqiUcSzQivw37cM1kMwvxw0mtY
jjEG3UI+jRJ2Pphm89Yy53/YVA3WKermxRKJmaMf31tawFpgUe0LypGJQCF5FkCGneMnsQZziNGP
lURGA1zI7k+SNKgMTYzNOqOqjLTyPrWRK9Mlfwwx2Hbb/vy0XIh7G+NAyDH0Q8AWVtQ6B3tzWTtk
q+w0nppKXowZMCGmdi5Mx1nJocaLKC6xOZMHO4urgMbbuqPUO5VVJvjlzGDhDho9HR54BBFvuXuK
l8kBfdkBccAEOWE0GQrwppTYl2RrCe9EzSMG3KjVHAqnal9XctDNEJq49hmph64Khqs6lKnddgBi
pd3gVF9ZXov/Xn6wvoRAtt8tK1Q3E1xdm53doc3g0X6Rj+X7QYKo94oXZlJ1h/zPCx7CXOeMTzn8
YHX8sLqPCLUWjJQqs2Kr0fbaM5wmJVj6/wXRbPnnBgHzcr1NTRVgr9e6EgXZ+9BimxzW0R53e/Dd
A3TrzOqtK+YVZkHAueUf2nuZKCqlBsa9D1kvLAmn7chr8tItsluT5JVXeX3s2+j4JHY+zXjtvkBK
xFsD6iCOJuscEi8TQr6kzexhKUtLqyYQrr9VZ5EBWhF039mmfHhe31ckoeO9PH9gYRfPZBnkpup6
PPakjg3y2KIPzYEmdAbPfjiXKmW2H12JMzKMUrjM2t2GJ1iP2R5QrLsynBPJhyi/WWSJZfnr1YFc
sllEDgkWItY+INhn2m0naQJ1wAIFq4mrhpA4kqL+zTc9lx6beQhgOMoxuJ0jbyGnP2dzdKij95lo
3L7/pXFfhcN1oqsK33A4VoM8vvqy40YABEyOtaatPclbmRmHNhSUihCMlV4Li8NFeScsb76KYDmF
FyNaOMfTqDftzzEONqcXkMkT5loPh0g4jCSn/i379+tZJDU2USJ24yMCHUKfJWaty8wNaJmHWqUb
XKI7Vi6U9KU+anWTRsgkSMiqw8AwcoVITgxDHEzhEPXbuph1wtU8lFfAF2h57w9RTLKfXZMoaUye
V0Ej+NJtMsGZRO0Q8zOmRBXW6GGvIHO1wCqGi1YdTW4UruJ1XvokQOyeXfLaxt0b57Tklco/VyqY
CoXaZNgpxjazMoOy5U2RdGIl808g92ow5v+dn5tto8CIt0x/g4wbnEqM4tb2oZ0BuPzhIqH+ZK+j
A7ewc1wY1ZhO3Wv7d+NLdYe4G2+lQ4SaiM9ct7sZ9PoWjtbVOkNs0jCEb9AKzTVlgEFXALuXpbBl
ndcsrSK1IxlZeMZw3LEbhD9tenikyO6Mu/SwLxOPTBmYpPak/l5PelXYB27Zpcxji5M5/xrsd3k7
diSnRJUNxYjuxqGU2ymuw5+Yw1YRVZ/EiZ1mVL2reSWAi1XznX+df0C1MX7Mlh3iCEt0DMH4m+uk
ri7jJF88oA91i/uAlHoOJr6x7GfJKe+HazhweDSTE2OBUnN6FDBTCBPAhRESa3lC/BbhkOoppx4l
8MYi/Cq2QuDuqpsfiwzWnD4XA5msYUiKRSBvI015busDfyrf9cP+CEmaNOkY0la/tVGZNqcGnlXH
/a5x59aCIkWHm3L23Y1Fd5wlCBO6VYW9+3hQWcfpA+HhEUARgWBBg8NMi71A8gS1zlkK22XHuJFd
Qpilnq3YDdwOBHlchnRLv50Yvvrg7xdsp7d6qz+XFjDm1d9laZ9lDBrDa4Bek1TtFE31SdaVTq4h
cs4BOPD1rS684+kgrauWLtD1+ZoC33U7IkroXUlXRrPdTtVNNWx1rBF/7+yTc1gWqKm52m0B0FvA
D9CLKXVQgQTl4L6rPb+8+PMKjfAFUgHtpY6CsLtBMPO64XPZFgUcH5J13LyOtph1gDn/OdGoR/OG
YXqaTZKtqylnzocIP4F3GTOTbEfg7qENgaPCPkiuji9nJp+mTsoeSdRiHmZ2VZPlalg2Ill7T11i
/z5NQgeup0GI8JrewEA1gNsz6bFWyKQqFIuhrJD5OCewuxIvq8JvlNa7w/S40XKwiMp5OI7K0OYi
t41WB1nFWkVzpwo5FldEeSxjmMXKRfqDgvXjxeu8F1mAmrBhlMulRnLiOZNk2wNEhXgbTTZkUiJ/
PKWTYKmwADCELo1Ye1hY3GoEMyEiKZhR094HHEW1dz/bqMuSsR8a2+yihj8QhzL5ngi6Q+WSCMkE
p6xomwN0JGn0k6Dt/+xmiynlcZKH8rn3vvND25+TnNGWmGQtRq5CU02XpRLkJHl256dGHAzZpcaG
rxYZqepaQMXTBZBO/Y76VKIbd5x+/3DcVGZK7+Mf4Ld05bLFmKIr+yLaQRtbKM4bT04T6AdtK4dg
6/B6Hf6A9HAd5cyDGnYz8I9fSYglsINmyNbFc95tQMcLm0DyNNalGwnoAd1eWL1SqbJQpC63BD/N
png7i4dF9S1J1QapNVPmgXL1mb8xqDFtmdG7TMnTkmSi8jWg0Y+BtKUJJdjUOgaSB4yhssmeI7PU
NvZ1M/P638g2nT4rQYtGsR9WUCrIFVwv5j/PojX6BqUcC+650CMTWpuhiapa026eB5QSWHmDGKW0
o5+gixhm0MtgrI2t9Zn8Ti+GXiwHCXMfk3SQBk18AGeVvH/buWBP6emi0yihqE4Tt0Q3kdRvYo0T
J4xX7bQOlq4NgypSiicwwfDzxP+M/FImrGZtOKdPVriRr+K22ANq7xue086ccHyF3GzB+sPNnC6Y
UKruN3ptabakr8prL8+c+cNsyDm0sQZ/W2GDKqm+Uq+WU/WLtNnjd5MNf7n5Hzd/Vos4FfD/+pLJ
Ulu8yeIivHGyXRoHKJAdE/NSrseK0EQEUZ3UWSU+c/FKsA22JeziicyG7f4vZKijUChCv/GeQLb1
OA9haK7956FBGR66hp/TXa5LqW1i/xGiV6JIwJwehtqqBlQC8ifbP+Bb8J6R7r8Db6KC0piCz0FO
y9YoAM36IoXDd5TvTpqCM+p72r3SqqTYlx08AyqpJ+kVptHElOzQeDzqVGRB3qJFRAsNRXZv3Fun
/HEB32vU7EicbIJ8I6WQZ+iKJF97CfT496aUQWjWJ99h06bMWe1lNpfXsVRlPuulp+xKI1vB4sU9
Ck/IBOEjxE1Mzv7prsDB8K/cQeb+gy6NdhdAKDDeiq3w2bHye2LxyraDxuhprkdnSh/nYBxqmkl4
tkdm/OxAXfPNJXMdNmwaUR4emgj8MIPiS4vK98QVxFFFIM1/tXo7eiyAAPK3ztPh9r0B34fYwdKy
VGGQacbejBuxwX6Hiy3GduaAwDdcxYLR+N19Y6SPIMdfGxnsflg3YeP99HU7Fi0ceZocAAv3FYp2
UQoZG1VOiTuPXxbZLnwDIdf802ePbu4spmsGjKnm6eCRmmgsM8BDPv4aB2UJ2mpqvTb7alfcvjei
8Q1RbG4Czc2sJqXrHNC8Mo/ZQjHzygT/vbJR4FDafALLsIFcvMtBNlo4md1zyeNUYpuECzd81f+R
+ex4AhMAtg6uH/z12Wf8fb5AyE+tu3gfOFR4gpQiyWtqTJcbZ9KL1/Doqo3FysO6tdrmFKwvhJAS
W9/91tNlIJGlGFa5I8DPoy4SPfNQH3RYMB3qOEfRshM9Bin+ddmttG0r4dP0uruJd7zNI6lCUCAC
ezPD1KXJJy8SbZwBojZpDlt4fKXqAfk7ll86uMz53zE/Ctcr5l/9NAWuw54xRKQf/XBcVQBBwDXr
WM/0/1txniK07l4vzdIr9VUnjPnVdE/F1F9fqwJBzkNNIgutjMKsG87so/gywkmOhv27Rfpmhef+
DAps16nowb1xNtLeK/N0bH29uRXKHt8OPDXPGz9RxxVaMLiO4ouJRZlNGgJ26LzZVwTQpdsRSTIH
ScPc1H8QfxQg0gYR0bkBzZGbTrWx5TQ7Qsg5yEI9x7mmgukl9KHGBsZ+CHccr44bgu+r3lueO6sZ
Fk1ES6QpHPPXM4tUXkJ9IHexTJehpSgf9GfupYwtW1XH/gv5AnT/xIeJXCrvAtJcOQbqvYmAK2ZZ
KAacqnIgx5OqFIK+cbPXrqlcBy/G7jwQcwUoU7DmcXFdzs/LaomDDpcvogFkxwK26M3Xqgpk1VGH
+hVo+5MN0BGTsnvBxZQ+IpCZWDwoPqkuWtwxxIRYNPU1llSHKzJRqqdrq/FRsCJy0Fu05KVOyy59
8FKVLo2EddHMh76Y2oKhysTl39zUQqASXUKCirrlCMjrVKDLxbMs5rJ8Ny6/roJ2vlzw7QcMzeEo
CIzotczo5QRJQaCEoxvsF4pr9W8MTWccNO6A2dYsEMjpYkOxRYPwNqfYkQqryJSBgftmXgVwwHcB
gJiGqPYAnScLUbRykpb1TdMti3s6afu7s+KhCsjG+ZImb75K2ho7KlXoaYPFAvHb+1s=
`pragma protect end_protected

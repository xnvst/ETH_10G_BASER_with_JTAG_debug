// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:19 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PNk1F159WoqRZjutIrl2IYtEswcLxSB9soLcxC/OE1IoA4XJy1scl5ZTCznxtDLM
o1mYi5tW1anJHqFds9kFtPeza0KQJ73I1TFRzFEno1RS4lInh5Xw59OqI2mIwjj4
3jjZ4CztT1NuOGTsxJO4nzQ/X2bVMBjYYdrS3eitetg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16624)
4g97XLA4YZyl2xlajUhmayu0kKiJ+WOAcmrcMIRgzkNxGzv8tEabWNZ9Ikz2B2U7
T0e26+mkOMLfZC890CS2m/kqMHLqTUbYzhm8fW8snmFKcSPYi+R0hv6KTeP9q7DL
fRDsfBiVJlc9YVK/u4wOLpRpg6gWt/F1as+AdQKCbGaeN2a5fZjQhHa4c91uiNpU
vMlwhZtnpN9K7e7+6GwGDSLi/UBcMtdMh736/H2fiyJ454lALYrZpHSkb90uACvd
soNaUkzL3DNvmtWMgq6kS6s+hRFz/8iePMFsDLWpY8tTqL0BHThKCTvfG2UtXHG9
edBirm8x9yxXNDyhK50AGl+iwoJDlF9Aa81YvlYS9/UGj9BanDCsShNrNudv+RhR
3V5Chon27hJPjvtA9i9/TVbDY6e1ZNhJAk66C/Tsz2i8HDCnvsDIzeqR6oKLgIxa
EU+2iEUS2YzJ/1JJiHq+8aDr7VtMqucPjK0ghUsGRg8iJx5knDkytz7fSqqs6WJ1
NDrLjAdZmRjCQmMPAxn6Oq5Dii4VfG1BDx/dGetyY9zFP/t5SUCNqliPadSU6M9L
udGhs9oMCZv2ZKPDcX5s25hdL6u2EW06/kdOYAvFTM7dalNlgyufdotQnR4pU8mM
3fKAfQh6v3HCrguNCGi9Mitbrk0PGY409uUh/0zhnksaDSKFvBr3DDWSU5KvwRUT
sQpuQIVL1T6i8sBbqvLoy2okJSNHSCi6RXG7eVeM43xuppknUO+S0DSRPdU/5Cwb
H7jbmwXGdgpONAoS7OPTEa5wBEXRzPQt1miHDxse/segBcgxPfW3PR848i4BgDe1
m3qXvBC/OfVgWLtszRIxvJBPbkefi9pEqKDJ1J5jt2py9HqyZeJD6FDiJwRH8vm4
c5Igg1JkSN7lXOJ9Es8I82rK2zJLErw2+I6czKEujt5CTlIp1dzt03I2ht8JKA13
cTCzQwpwd5SzpfG/s9pQCvCHt1L4SPIMhSPGwJcg3o3jE7ebbljVzLPg14RFlH46
PYcNFlZs0eq9SIQB1krLhaNiGntVOfiTzpoXyHKeDWHAga1Csr9hIzpYQ2hkHndN
ZnM8TkQiIoiDZyZa+JCuhB+ho7DptZcOyuZl40eY0ILawFOh0f4AH/f7aDVOCv1K
IYJPPnM8g11366n+AoTx/fndE37B+CXO7UarabWHohYnu7QiwMPbp+VC+bpc5q//
NSQu5SD8x3EajNS8VMMyWCp8Dy8Y2MPMcta1mKoejiZeeHqYkGwSNcM54o6wZcVm
tzCg5gUDO0yV8Ng86obKmI2Wz+L+RkAY1g9XDBXY9/hGhjLJocOOMvedyX5O+AUy
L66yuGmfDYCvocJl89vkL5pXkE+pjE+/z2bUm5UHe97XCXlMaPOLvvqTUA93ci51
ahWLqaBqWRVN6UpG3+ALXinKNzCn3qVUPJgXwfenjFACPhjQx41SdA+2MBWoFmP4
fzfmt9cAbbXSkKoeTc74i6jtC/R653zRQiSelkGYx6YaERnKCxl5dntuNJBseHyr
MHlJu4MuC6B+5kwyOAzfr/oKTLs2xMy6XCEieDpf0xkL2yKomcJh/z4xlV5B4LHT
nEpofMwaTBzoP9PSao850PL+KPNPoTXrD5DCwzu8LjESUijqoj/kRBxMWMx2DZB9
RZhTXvY5gaTRn1tH60gL69LW1xomyibyYPeUmKMu5yKnF4uWK8JdPxclXyBduHmA
I534Jiwo+2d1T8lUCD3UgjJUHXKbm7NvJhSgcTbAo3W6DYSsZdKYLquQsNgdMORi
tU2n+4AWAHD4BdNnM6r2l2mCBZHa90VRrUGdP60Mg0861hHm1R/LIdaLjQWZrt0D
2k9XjLCnG8H4mkrVPNZnPLdU8Yoyk4s5ru5exIpBvAxawtIhaU2vw1HCLMLVFrZq
Z1oc5GML6FfJlly33MVDsqrJwBGgsbHLMshufAU0v6j9FIKE4RqTMYi1oLfuGdFz
LTYqzySdNQvKNA3mimDFt5rpXzNOBkljya3amsZXa4j7ZscRE1XuaUp7/x5a0kH8
fLNIvUdAj7wsW2BHfJ9K5ucjMMYCR+7gOPx4q8/3iMY0j7RqL9Fis8bIiscz3J/T
rPj1jDeJaH8N8DF0WPqiftI+6VCTB+rVSCHFup2uiDct/+kTb4BPGbS7NlkDqjb3
OpR8lTQSG9vsTBJYmmRv6RQiJ/bRATxmWC6CFQ+PozSVOI3bXrCWrPQjYgICd0B0
Gd7p4cAbjjG2DcVucD0hPLLWuRP8wpvmJIDAhh1n+eMLCR/h3S6Knje+eS5k3AZc
Xtdn4txCVuXt2D5KeW2TDe73HKl/rowlLRDxm9F37HGsi/F0/Tq3M0AzfCZtKeNb
IjY8rFj+buBcvLJiL+3TX0ppduRayUzfa/fgliZFy0p+6MxZZD495WbfozXHwxOd
8jMrAyKJUhR+pUfTBifFb4C6VRwsS/LmQAK4nPgVhq87UKCnWYeOlGblAVmG113Z
9X432cvGS63FPz473sWUjR3Gwp3kbAisBOmKZWBuW1c+6c0q77HJX/mrk/7WV+AA
P8zBpOoU1GFlGiotPl60nsndQkrcrN62fqAYw0+SCjgB0e/K/c0z8JZsOOUm31J0
ftQbG26TfV3uOce4K+xhAoZ3KiREPELzsQTOeybnTZ3666W217MlXNpBQFrfjKPT
UaLgmQUhFwgFUSdFhjxVPQVzUU1cGW9ugaDWY2whPwHDXoyGlhht8iKTFVNl2wjr
W/MWypea6riguDk1t/9CGnV3twcPde/+QNl89+1KqpYR+oLQalWvjVl+y8N/NFmf
mnUEXZAt8sve5s/oQZ91gYDNyEMoZub7j1YorPy3ZdsNGKG9/phbCGnsGjJSD0pC
xCrqqmTlaSLaYDeKkmikxKUAd12s4fkLDdc3apRj6GJmLJmdm2tyDIED32F+6e84
KZo1RLHV6F1iqE1IBuHnZhO4opLDqEdQRCSi027tpcH+nShSq+otZlzycfTtRp8A
G72MFR+0c+LTaZckBQ3HznVCaEFn+0FHDaGBfS/oaPwjCPdX/Z//jpSe8X4lAT4m
hYd72V8Zjvenf9bIblS4UU2/2tQuCrquJq80W+5f/2CJG+ydqIdfQ/1nMQzFRlTN
Be+NPoL4ecEMUr42stP0I9h6TDeE4IiTFXm2LQMPmaDiDlalV4PFqG/3T9ATxQE2
beOOiHnbHK8QytjR9zo6fczqsGmcQZHgQJNziYLpILptO/5Dn51SGSQCmMivD6qA
C+Cy3EkKsZK6PH20FPtVsFK4pHaKq0J3tpSWOq7aKL0XO6iAkhPe0J/khidt2U7c
AqY+tcgTedKVGChyePC5Wt6qIgwBq9FFdJ6isohrDGqADk1TOeK4v0g1hpidzbu9
7g6mzKaWxnodTCbIrWN4nak9V8+keAXHMqvaYcHdyOjuJQ1Y1xBWtbF1Ji0GNNYi
H5GstPdbuaf589VieKczvBED+hreQCasXLHB6jXblLZQKfZNW7PTLsmcD/vc+Uym
V2s4gbSRI/oP3B/BiovbJC01mKrpnp/yH8w8at4uHRUqFUfGNhW3+g6xVMgjDfYl
1HzuT13jWh+2eGp5DvprJqblATjQ0XANuf4UELt4rVHtnT/lNxGJuiSO3yu8Hqz6
12J7iBQEafDGOcWja6YCvhMDFDvZjytMePnkWSstwcsmy8M1ImdG9O29PV4+7SPc
BJ9WnxVD9hQ28q5ImOmudmvEr9BVpLFC8Ecdgv9bPPo1/DJAZigA3Mtt9rZHFYRb
swkBxvALvZcDx3VGDjoaAElW/c09vE/5GxNlxPJnBe00Bf2dJdGHm3OyFWU6wMsc
hkj8tDqs6u7I03ZqrABkz5skch+8rdydIVcZRxOc+Cac2usVmr4X25xHGgaUADsJ
OX/jhy9Qb+Fi0LP/MLyqdfWwV0vQrsG6mwF506089r+jbpbh3LD830CUgL0oIgCM
vmxXsxfv8e650jiaZyk3HDt0o9A0+H7WwfnkWpYoh3DxZXwJXeNw/qv42cjK69Is
1qPF5kLS+IDGGV/sBZnbBpPVuR10/OIUNLa6J4tqu0qJK2Bi65qvA70wfmGgNBeO
xu6g+JLYK99BJ2HovN1cthRClAp+qX5oF8S6JvTk2iGr8hwkzEFhoQGPX1lXtkJA
b8PwO5QtuNeR3p6U0lrv+FuisqJXd4xo3NZx7+azcsv1t7MIoeGxBQzWcGanY7LY
aiN9v/Jqtz+Bn3RCT7+dCrgFHGQTVKWtlBzSB9I97Z4gue1r9+A/+yLc+S0VA+pK
vLT2kDHNiJoKXTfwV6XJfmV8Cs+qTmaP38byv8Axs5AXl2KQcMnVxOyB3mXQSWoE
UeSIzAfd6qZPRKXpw7UhRN+ifI/EYf5JweoBHaRzJdxYTY/e2kYfhF+gZkraAOoF
6A4NsNmCXK6eNJsobyLArpgaUrZhFpu6/YC1jo8+VN7lgeEwumhxBaB5pvInoY++
AIaJ2q/5qNamqruMjooS/R4cUrrbItX8cbP/vCwVC5RGkhOgL5G9QUH7Hl0t097g
DySTx6fJAo5SmI6McFKcfLylQtgvN+2m9AsXfUC0ZzcGOucTzWTdf59f2Jgt9s2y
aAqYn+Q7KFgk9AZO6BIg8U+dceL2ECJ9L7s4h4KuB8Uq69bsPYNkepmTb2aTfSxy
a02t46nfWlksh2P7hJ1guVPnYuinwBGqSiYtLmmP138zy7SX5fPZQ+LhTGEZWGuG
0S9f34MARsJMszylniTm7Nvg0WM8tAJgddHaGP1B12oLrUGiHxofdC0NsFt+VU7h
GWSvIj5wUyhtIjhEBEJIa73y18taQxIN2LILx33lygA64HwQio4dSoKiIbwUUAmJ
Gdv/Lx3zIXVQpUDILP1Kbsis8BhHDHpAfo8+S0cYXX9Lj0cpoQsIAsy8nvKoQULU
m5ngSLGpboZUfoQFCaMvey3C6l+0LpQoCHXR1AjjR2h0qkf6TYc1yRQM3H1FRLkl
CuStr1u0ZtROKIiT2L/AHKEXLdpRiWIaum8RItuak1naOs8e9iQKqJCLKapNontH
qdmNxM8ApGZ8TMKpSwCBxRv23thTeRThl1C9h3uZ8s8Yv8kG2udX5tw0imGhW+I4
1OpgJM88YRDwTTZ5F+mihWGpUJ4yi1riIJcaroW0tLahmA67CwNA8RhCbxGCBi7q
XhEbWrHTe1s5ZPlpwqRbb/Q1nAzaSvwBF3uh5x/rKNadtdSkYufRHrxvx/elAgMD
1YmAvzyZS6t+xHvRcMVS6XRe6OZFAGdcSxdPmBYGxx9FvnJ8eYJX5EmX2WSJ9Xcx
wVDNZ707SLnwOfgJymYorYnV5z+KKOduufhPD9nPep3FU4ArDgbl4NA6xlcl2D4Z
vnBgfRNVi9jiE4T3A1gqHzY1wshAhvUoZ1ot6oTTDEFKuYaouzRff3TxLYuVKD5g
O74+Zn21BGG8/BMZlvU+CEoGKbog/mn+IC6tL7E2kJkCJ+DK/theEyPLlKsl1GYD
vmYMMb6gBAqIEfCkIuOVY1AUQpfXVomxNestte6+IU8itdnGQdNa7xKGZM03Mwzg
puh9NLlPEo/gRRZfDamdUxd7Yyhw+v2WtUd9Ma5gRCvzWdibBQAudoBS1YoiznQc
vGRwm6s5fV1pRwDDWBpewF5pdo9Vuehg9VZTJCBLVaqvpi0VmKas1jAMVTiSNMDz
G4XtJxzKuEVBri28Tc4buVyIrcDeln1NKN4cYsJPSz9eFzxLWacsyLXlW/zBmg9R
GF1sLJnoU9htStE2Cs6xTfiB4PnNivWh2w/yNSEJXmYoV2XDmmgFNZtxN9ozHI1a
YnBjdmSpdMWeGWsDZJs0jMaffWEwiPLGc4M/VC2Llot6WnG7WoCbCafsQw/RWFHz
NpRGTHG4rmXbLMtf0bNeiSWCGf7aiIUaOzwh38UmZnhcL9ADKFhaG8psANRgd3cI
86/QHUsrkCfNDj0+YKHAO3YimgivcEEIaGpl5q5WFRJkzUakwYDkfFeFis/uFVYO
17Ke7tFnPXNwsyokGY9xa6bANdkPVsRmGNVoG3nYEhBBk+lcKd0KOjEa/0y1GgKx
VOI9e2c7Z6v+RXQVNsw39KyqGpZ3sRpqKMo9rLsoxCXpc/ZKwYoYhmpbXhUlydAz
wFtH5oK7qfzMa2M/mA4eTKukmovmqMtaUlD600WoD5q1ZYfJTgj5Swzakomr7yoP
KNDY/0IeDjcqzHcpeJthjt8xoUcOhPTYzUrxzE7a5ZNNnjEB0qxHjPwIDzrHTdOE
LJP+s/l03YDkBdNMOV5/zGG2HDxxUU0ZPxHkwK7h62kq+6dE1svHAvJqdBMJbgDJ
1axu12dOYKyBycv+RVDo1MW5MDcDlZkVq9fYIzEvTYtKtz1gNKAKgI7HGQwMoy1I
O2rJi5oQXbVgx4LlIZiis047MCwMzpnlnbDAy3tM3IA3oNIrKUnis8zmtub05K0O
JiUqfWCNVNvzW8IK+W+lLsVwe7V/o65K+l0pSpTuGQtyvwVbEazvxL+HoWKLRwlK
7IiwYyBknSB09Z1broMyALkPteiNFmUgj9c5zXNQr0wfu5DkR1NWRaxhlMOrKxDv
cJCYh4HPTY/K5BXC2YZ558T7mdkM3DWDsqaQNFpYK3Uaept+7NyliAOk+lBnFZWA
57UJp/Yf7ZrRrKp1dgJnMwI7iR8Ao5nnt45hoqfevFSuU/FsuzM2u+OpVkZvxRan
cOaemzU1LKRM5DFOrkQzxSD5yl8MInM9OiTr+Dt/VH1O4bgpdP4L04CTlwoceYNI
Fr8xJMmKHunVwwKrDYj2IX66K/wnwmRGo8p5i8N+9dAIYYJ8ZuKCrdII5hFa8oKu
EUwkFW0lRH52hDswMtUv1GxPBo8mFBSaXmQx/+yJceVCgDs6XMJEqbojB/RbWxRp
ggg7r/PoLiMt7f47jtOZeIVITrWa1tSS48ojsEBjDy+lbC2F29OXTB79jBVHN1aY
/cNMymStvUr3sus90GuLkYWD/UAd93gB8l/lYUsADZsunVS8cIVIDVbBNEDlHuz0
MZ1QONXKNCYkuqU7vw0mxTqjh0eDzr4v/bYYxcg5nX05RP4pofIMtzR/dSMTXDh/
NT4kICvw5D7TrtvlFjRWEeir/pySKjPc4B1h9ElQcf7cPLHrVXwT9o9IvpQuhovM
kSSgM4+zkyCUIq8sU+x6YjN2uoZ1B3g+Yw/gdSsT4z8FmXJukgX3NFMcTb9faoSF
tpoiczt68svWGt7jrPN/QYc3mP3nAwuZnJeRWyeMKUZrRPohe0hBoEyxLTKt60de
RlXT2UCZBhLGJWWgWbFIBEv94V+KM3gk9fm8EY8yY+TnELOJf9ZR7WzNEjIbJTfg
SGUzMMRD48PKbbELPiqSW0LqqL8JGuxxZVgv6fK2M3YUmQ3eBCTFbCIOZNcq/QYd
qDfKLnVdsvzk6U9O3ip88pXmi0tkluIjGKVKfKBxatccEJWyHyQscWvyzYkPCTdd
h9flhOW9oLUAWF7MT33qOr+d7p+thMhETLEmsYuxwZ5vnOQVyvX2IdTFGINmhBwD
yHhB+q0KflnqZj6AQtLVQFNS0oJXF5363ZYURMGTmxid3gonFFclabjsvaPV+yJr
CKJ3H+Dey5/CvzlcnCj+BGUSJ9GRurz90luc2sBwKdJfbC1XUOY+gQ7lIJBue05L
SM3Y5DWsnVgzhPmXk7zHHq0gIqYYPGba/jD2QRLJObg2wqZNsbYrplh+wwl779dm
TiB0Yy2jLfCFGfO8+7MXxzRscVV7zZuZfQ3g+XN7krBHcjP9oCRWbuNmsfNLc49G
AglooyVUtTBbYD2tFaao7RQinKWXvWJYnJynxJLoD6CjrzsYA2qAmtAab3szf/o+
vJtv4KFyL5e+LFEN7UlRD/xbmYZsnrLnYFTnNlA6YciAG8XzqlU/iNLNKVXVWkyC
3a3pY5n8M2CnYzjhL+o/p+Wr7cTZi4pox7zNBXe4G1LuzwLgs1XrRf3Xt5284//d
nC1vgmSZgLJD2JeygsikgsHQYsboGq3D+cd/DajIR6WQ07kJbzkZhMp+iKhTUejG
VYO12eUx0ZnhKrb5CeWf8fVjXonWNWjISMpXXN7mmawqtA7WPbgDYi8+xa7+MgF8
sPDD+MZ9Q25yRNTB5cr3wluflH9kLGCjwjIxKdeweLrSSn3T/8wPHv4uFUan1VcN
BGxYB1or/w8Bjs3bhtCogcYVIxFFe5uab6122e6FGO9E8gPXpuAYavDMxbJ193Eu
TrRaoC6z+OSeklFREfmG36xdHrxQxcOlcD4gWANyq+ABbZqEV/Y9qhfg6DrQuj7G
zIv0ql7D8lrEKulhxX+tOHDxilwZKvOxkCL9ABdaOOArASkstVFVXocPgOTgyaRW
IMQhICg0PPuQs+ZqnB/Qrwp55xOWSwhslRnC+vUq3LB3s2pEdYMiRqZ+CDSE55Dq
5XwoB5CAaheP/gvRF0P91Sy3ykv4CwBIL2n2FzeXkCc1uimtMASyLTPH+pi2zix5
rqHhurvLEPFwEByZWiVi2lnB24WNFeMlLNW4G5CQS328SVVBZPRNsBZhziFBnuKu
6vCTdi7bYSb36zzX3M49pBNJVc3v7pt5+UbiI35VpAk0hsCvkJ/bfQ/5CzjiEAdy
OjoU4w/wbYXs0BqrfY95WAcs3/RYn1naO+wiovQOVBdE/wUP6ic7WWxMLTiw7AAJ
0cZ82j3+uOeMIJuH2MD5hCSXWDzflojDJeDOR1aQBCeBCkx9P7TIa1vkceM1/Zdy
hYue3Ay6uvlGBECFfENCQUVil20JUlOrxNFzBxNEtbbw1bXOf0znSZe25LBK0mLR
XPLs1EPeY5OUxGeXqf4jOx560B6C/otmtKt1TUipIZ8vFOYLf1S4EjJWnNhI4OrT
5xpZUVSsLNdFhP+XZ5FDm//3flPZZWRyHio9z9b3WZlVpTZEtO7xbB/0Td6rkmXd
I/NaoyPiJswfY/+Et76Vpdm7uj8BEktMROHaGnljYugiN2dZGwB8fnrS1J7SXrc4
JsGLcQqooRw1t8+zI5gE7l7wHH9oE8g4GzmRanpNBgELxIH5l2+ChdtW4xnAQGRE
H3jmvy4+Udu3mFTXfuUEqHt+e/g59+weB1GGZRzQhJ8evaLJ2wrG68F/MISfIylJ
PgJFTzCATpSn9E6PMyi/Us+KYt9sBJ7BIzmQc0AITc5NRK++MSlbRTso2w6LBECe
112T/eBlZY5egn+7eVJVudUjxiK7ZDyS+gSJ7qhOCaQL46nsSPiq2+cJhB0FNMFG
DRw+cauVkIcdyyOKPxjgQmGieWUIqYcfAoU8VILs+GnJxDbbismFbjaJbcR0prQJ
ts/P0cvTvXgsy8YmNBScbn9LxRECCm27IRSBDE53oS2cWDGKUAKL9BSdBMhuK4Mt
Rct1bYXvLF1NCRH5wXx2ZJKZ9Rs3EnOonloWbFznuX4OzWtauA97FH9iI0QeJjMR
4cIKzy+gPIvAn/8ieVjhosys4OtIN0in63awi/ggof2OU9ZDEeYpQZhBXuxFXIpk
YDoufoqY4KHZXNVo967TZDqcA+qpz9I5D2pNh1BpXEUWUcAUzadfjASIOgd7tTEB
eB71RBOgzggV0IUVMFYFvV1OZ5kMd984RoH5pmbb8Xe5DcKydHa4u2+WhRNlm1Qn
zPUgtZ/hwFuuHoQUvjN9YaCWxa18gfhldLBUCRR8DskY2AejYz0kzPmln+z+zFEz
x2aqnMVfOipADwZMJ7xmp8+lUgb0NhQqjyTcfLStYsaTqzeWW+PgY/Zb9F+z7pcQ
+Zu84PalnSHWDypGyNBBiMo30FW98VfrcEClTR4XPeVCGmWUgr88Js6wZDPyQy85
Md+L4g0/6iho7b8uIayp1vAG1h7A+lnu6yXqkC7ANjXm/yc/+w+PutJmlHNh9k6N
rjTkw4okefRFhSQ1XETY0LjuGETBBIB26qCDE2r9pfhmTCRpSZJeMpxrAZxJj7lK
H33tiGYG7520RXiYGWnOBXSses53ifoLZZ1FLngRgmsuFtYCpwlwQWeBGXBr6JQ+
jJ0AXu6i8taenZEpXeyzXrIMVb7BdJwCtNH8W5jCMOJmxS/n/fSkW0mnvfiuZe5J
Xff2uG9J4Oqu84O3mHQPh/kvF5m41QMRgWqRJ7053/Fn6umH4jomRzW2ZM0uEyCK
jgNmYF3LRDTqkTI7PrQCZkUNxd3+xhC708s9nLZOzsBWo0e9Yi8kGQYeQgKp9tx1
HPtRx+sKEmqvH/tWN6PeCleSFZpxgBzSITSBQm7nkF2YyopDQS5lw+FcAC+FPPm8
IUuyPjVWn25dQ0UCWlSoj6XpJxoJzuhbSqEsS/BUBq6GjkEdFpC+xU+EN/w+hqWY
KxkAFYFoLKecfo2Lzy/uuolTiZnD2l3MAlkL8wxwdRlwZ62t3WBSgxn0eqI8aYLM
T0dgZdRNQYonXwVygOvpYFtLFmpw9HBXFPSxcbtGRYxFo0tRQnoWrKFk9hE1wuF5
BwEcQrzwc6k66XPFmLem2tCm7yOYitkgSrjRodJ5/7ERAT6L26MXotSiPXGK08ru
KOS5NOwlETSJajQXgxrqnswzPTT+HIL3o8R+cjd+lK9fr5wHnFAdDf6/mDPzOr/0
76dj+0FQ3HXoOYRiWzlxg7PAsszF1uBKjXmhpWOl/+NdpKZ7i4LePy1mVvzJqndb
BNTfM+aXWqTJ+QmjnIv6aCXOWciwrDjpCdei5eoP+4g65LBobWeExpfL9rucAJX3
0JHDMKcIEzl2zrL15XqNIcGWCMP6IOlFLpf46FnkLBcfaUQVxrjEQYCmA3xIq5A+
MSPql5NmZ5Xs9yTUnIkLd/2yBBDDJgR0e0548R+AKVgjogSsGRfxRh15c6OirYO7
CNEHE+gM2unhTxXbWVLoYZs1e2pqnbpt+1PDFwQEUMyYEdzcf+X5vUaiqY9OeFXg
zgEUUKW5qxBdiLdjXr8aO7Sdc8CfwliYYY6fD3o4Q6jWtwPrwjBiqoUPj/eZRf86
Wku9jzpvEpoAeA7zVpbkXWghxl6VRPENg0CRymaWZe2fNHlwo7HPAV/smLu4/gtJ
fwkldkPa+hEjxb5a0YZkDYfsgUlubZw4VNuYmfdm8Uh/rzmFu1GXe9MZf19DSRMn
RPHPxM0gHkJ9mMQ46pFcmfJBXeMDcKqiv84J6pBdzDs9nBEKhY+hOJy+kdLUSk5c
3C+DIWrK/pYCkCyawiAB/ENM9A8q+aLpj5W7zOrmv7BQagzLT41C6E2rOi/S+8iR
dw0JLJ7glrTDf/y/vpATgG7FONh8KL9A0TkQXpiAXZEsuBoNEU9tFOtKkkqydvS9
da5Fm2AnbO39+gcugLn9pxQb18yoFZhHs6I65RUsDv1+mB3+GH0zAfZuRBpKsQGx
zdRTgLa/mrbsJq391EBoO15KmlgPOphwqrF4DmgFlcJQayNlOpdy5khbILfPrIhf
GG29DmX6djYWpmzPSVcWewrra5Cz7uYRINGKpRGg2YHUXyEdcIgKDhyssgjSO66j
5PAgd7wRqXlIdv8XM15FtVvWbYjrOG+7uuNmXbUXM7ydf0IE/j6WqUSFrFmvOh5d
lXbnZZly4j3mCe6kWm/uXU4b+XtX8vvIsA5ruSd4M73CT0QIILPjq8zxDhjKrZ15
Ywm8Fn0zwLSaEtOAoi2YaaNEZISx9/5OuTud5DH1YVNIV2aG2dkECS8v3sk5krVK
2HciSkCnzu87u+5mEkSupv06HGg8HLJFSdnF0eJSaGXzKH2gyjiC3HSmrCIGEsoO
XegZx5G5rZ2/Z9GRQ2eXcPkH+oBy64kP4ccwuJqj+bUDC1nFDIFc1hwuS9ATugEd
alKDUMpszIJ+NwVtJJfEVYHKXyR9wPVn4AhmP7ljs1tmjj3ZIVHQPoXL82Iynp2i
VNtd1ZpO9DgunYvDal7JypZp5xtL2Uyqp2J28voXYbWFZyqOXt17DF9k7mo2NBvw
DWAfVYr7zp1lmueHRKKUP2NZBGDcoa/StRxPraNRS2bNt7YmKJhZDnlOz9NKkouF
mJuXyFFmcxOlFO7RZnJcCX481l27rGxl0xlSV6SC07aCEMmMLdkx5SZB8TudFW4o
ziMmFh/D1E601MYxtVUE+PH9Lf+F8kOsPwe618P32NlKp1C29du4p8u3WxdyLup0
wJtVvslXfdD5mIpo8fVI86s4FDpbMG4qAwhpkwbbiAejhmlovvLaM8mMw/gHM8Us
t1xN7oNH4jr1I33ZuxOnm7GH/ivQNnrXQKzOZUJ6e7x/QE5SUs4e4o4cS88KhbDz
MDqEbLdoqTNrSvQ50vsujgfAmv3Jr99Cules9dpXlCQrGuLPegBTxCZoNNv4g/SF
8tGK915/TV15v8Hv2T+2EpBOc4K7fpHiCLTAekM5SUZXEi+D2OVhuBJjuZfRgeGp
Ufy4KX633pXR1O7o16QjRRDB0v32ISljzLhKPRzXyendIY648tO25npZzFkya1RY
+0DFWrFeYEySr9qwG75UosxK9vJwrnDpW83H7ACoog5s8P7KT8USs1Cyd9nQQbxK
5jauc277dIMzmmbnUXHYznU10rNVQPdE5v8FH4fUDu+DmejJd13/s0mzrNDYZfIc
8uZHtgbVj0coE4dCK5X1WIC7JW+5t9rL0WMhNr2HXQTSnqUgADe9HISYATjUyh5z
IkM77DsV3uEY0y0lulACoyFVT2i8rDdEXCR92sHgua0LTcaw3kYgMJdEdu9aJ7vY
ZUnDhoZtdwXmgSU8d4rRWobatZF69zkz04/9P2gcEVaFy90DOAieBAnmGvr29lHu
H5qfBGdJEjYoS6IlcJSqpW+X+ajWMTt1IE/0XzfrMtvuU7fqQdcBrkQTteRIH4tw
lMZT3suUPQjPN+cBa6T9+ygWYVdsGysMUwKOO0/Y9aVYOwD6OycwF/4wyB62vTlt
PiRddBFmQghZYdpvJuGvBtTucbBfpcwHve+wfAUmwC96YR8B3fmx3hsHvsLuoDkD
yMBNLPMgGMc2w4wcdj1hX7KWkuhtJmmfklWkqbEFnvmjkt8bprpKUmMf2FoAFmr9
p5P6JglASrSj5GUxM2sbn9XqBr2EKntSNoNZoDq/4GSOAGvXY5El0wso1wKhr/mL
6P44oVr8e5V7jOrAdz9JDwPyKQWjV2YRZnYpgCdsTp3bu4zGUdQgoS5MnpWSF3bg
XUGWSGEBc+8LTuuiuWPjLVinXAOGz01Oy+TuZQPA0MeeWqB+47YLtMen2WFmPnSA
kKBJ0Y74W5wJtVBQeodRcjrjvJdX0G4y7n9tLKQn7umAoP/f3V8l/e/GfI5Md50P
xALZS9IYE0HqJlMcySnEpN+WPh1LS1j2TG+9jhECU4fv2D9iMXosrUTGFQlsZVnm
ApNRYP0hBovcKL4i+QjG2vK2Mu3Xwh0yVn6p5p7JpE7oHpgQs4KP3KeiXs/gvXWK
cq7lIsEw47Ge5Z6ErDMIQW9T5KCsnww888UwHVKha4UY0mzhrA092cOL60I3p/RL
QmQLLmJZw/tDnL5CrE1Kwkx0OGLcHySkYRY5B5mSNvOm65Tq9AdL/MgNWs+oi1v2
VkYnFopFbV34Q/f6KD+yiDk30O8AQL9FvMPrpOyoDUHD08o20sj79HQ5QUEyc/PT
d4luShcDuWqA96UKwmrgjnxJD56bhUjYKm1Q8KJjn4bruf6erhxQJTdNRJ2W+YHS
u1wN97B42p004HopGSoQga5249GsnHchegmKO+146SgeuN8SbGoP/whEbKmpvPtW
IJdzx6pray0GHdKWFbrYQS6eq7ocMAAOtE4lqOzaY6df/s7QkcdilfXpQvAUR+FH
6NYXFQGBr6IREg0bxsdONoHSCLltNIQau+GL/AMlhzKtaZu8jWIKtUR+NSw8/D3X
THeE5DhDgd1lkoXt9/m08kNeiqOUU1RJUNL4bRkpazCWtNJ9cnzM9mj2AFcg7nts
CZc7H9Qmw+K5752tZJduHIvFu8uKl68V5gLyHRGa8B6ilH4sIZW6TMNlwX+W0pF6
NXraI78I7Of76315SdYQSQ9y+6CXI9wqXXzzn7EmwY0VfyTjbsj74K5EyftYVD7T
KLUh6WcP+mw+h48cVZY8hj2vM47LdgANdw1OKwv4jq+WPchRw0sElvbPMkSCZCrW
EC08fblErPiS//K4S6kUm8RGisMSBGmzXxjJ8tmcx5/Le9MW8pCyFyGpIfglDS5x
Nb+w3CqHPR8xEMqYz/nQkrrbY4+lYclzo82dqTOaDPbTO4GpfdapiDjKVwX7ky/q
gqgirW1YpgbXxlbMrAHySM5GjCWOHrhvSz9uwdzzklawMZpwW6LBE1V4urAEmtm3
eluj7QQrDEIcWETe65qQNkfOvgqDnLVPzHM3o92wTE3VBswXpZtNZRhfaMp1EujH
fuB2SdbCl8fRTgHYT6cdO+1B0vWxLhBVOYd9Jwc+gMPl5DiApGA8kPLFVfnfNX9z
OsgCRept7UuoZ8wcKcwWQRIro0c7xq1u5eUK2Q4SJklV5I3A/H1yBFG68T6oicbu
UE8O3Kjp9eMh49cG3PPitIEOqGYDqiWoriF0L0Wc4WWBR68jsViEudOWRJY5Y2c3
ACD72zd1wGWMKYK4AGlb915m1E3Ztzj7os4xMAOizpJJWBLX1mtm1MFTX5GibrVW
l8yYReteINtCADJYjBryOYNPJg28zoV5xir/1oepcrzNd6qieJ9cC0KvjrS/Zafw
WcafNGi4/++84NuU6JgwZxMhxRIVMNnArUf4sRod4u2AJQt/DCqr3SHkG2rxNqV4
dZjX1vLC4ms35fH1hbsoveLI7PbeZclZsBfw5fbsfQ683l2koGTu0u32jeq59pN8
Vi5SrJcpcotylKgirj3Mp8543FwsMC6CKTdERnfQOBA4Agt5iB47uAOiueoUjIxC
rPm74T/b+2F3qMXgo58LZkZDVlk0IDd8z4rZ4X3Vy45I4Yvrn3Dmg3mAtdQreQHN
VIB09fElwholmMXpf6Q/bpZ2FIU9hiNuM9UdVNxZ5COh5iNGeBD281hlWOkMeXgK
B25oiok37m4pHj/5gK72Y3305JkhijnIK/k14iustYvU0Kdq+56oBvhsZ+pdfGNv
1owYVB4hnwOdDRqngZ9YLKrXOu6pU32z+qpuNx+Yv4wr+EXOh74xGnEYVErThPHx
v/kHKZMdG2bAI49RzLw5eCbJOHHTLjGqizIpHJEqtr0mkq9V2CRlej0qyTIzIjR8
kU6Mi2UYMBLrfuIK9X/X0r38sXH2znsx65FNqBVlH7BmmlYX3Vuz9vGSrexF3U7i
tYwm+19ELHmjjqCGnFeKpWj1iTYu8cW77qbEcDSUXaoeHGUJJOoclixer3lMDBNh
zhclqdsztm86wy5Z223sQNQEZ4C8bOCgH0nFIR0WBwrul/RJJsRdEgdn3+ezn970
0cOI1OTR0e7p0VMolyXi4qhXrMK7nXnPxNFe59vEmz3kO2lfpPF5tbiwn+Fl67IK
jigPZx749dZVNL7alHg29eBviJCn/AANxtG2vn81wDsn4kJ11eJub9/Uo51ugLpR
g1AGBvYGyNpydZpzv+WjderIzlH7wS90Rb+koAavs1GZ00HdJ+3eJzuhvdNh4jLl
CocM0a2rvwVy7QCbOJ0errakXu/DA8M5GK7M8+C30sjAUKK5SoBb5uQDBd7Y3FRF
JPn4cLcm74j8J0pid9CesD0EnyQVLFCkuuIsflUbKVaL/PVyu6SEudTBYN7tElXU
J98LugYlDjl9erwYdwQeq05Aphy3shxP3e0Ep7s3KJfLZBLyf6tRkaN9xj5cmDhI
CIdW8IhgrAjFJfFSdUxRb11uDHwEUGRvJtQqBaDfemxqq6thusiDK1F7KFYjz5pa
4rVjDCVfpf7TaR61zypL5HHmI94VYQiq6SY38Fss0KChi+zCvC9UvEuQ7XVaLIz5
o1mGxNCuIoXIDI57ou7ypt9HJt55eUXf40jVS4Yc48Xr6DonxztYvuo8L/VF3vRs
2LU83tR5e/H3p+GBYD1XoqnqAcWhDxeDHFDgLole7nKZEsK3O5E7LSSnEitB9cVp
eYXmjspqI+2yf+J290Pqm20rdsz5XF0BChVg+GQUK1/Z+Pv21OFaJleRkIFdOUs+
UfIKfByJWVx7Uew0YQ6EYnRG/7FDKYLFPJbanS58Qsj0vgKo73el1LBtUhqd8Tuy
js2Hwv/2APZ3X++WqsHN9Tz90u8p0fk0ZKDgWLj5WdW4MtmfpT2W9bJ4vZhmr9Z0
shgwHKf1dP60n8o+bheoaOSqxRc73scH1UvWBugaSYO0j0+V2l1yNUBplQuykhIw
Kt2zXm7S2cAKE5WzO+vGzcD8MgmcPVrQRtEbpoSCjK8wTsjMYsP0qSmoOBoX1IP9
IpjYdRApoSDqLbLtaMzN06Hth1Pf2eyJ37X92by/bMHmEwXV6dz2hgRpr9d3+WaC
CRrb2sH0CHOjDwHI0yodrJgYjf8vn8E/LSwp3Ya//8Px0ww9UN4PgwfLIZ63AiSP
mzvJ6nAULM7wpA3z4M86yrhJlDMbZezaekQahkax6maHClegVEb7Gi/wClZ34QnU
C7pRLEdkx3OddEEo6oF5rxbeLWoiwuhe9wlGfFa59ETsctzq1q4p3hJx/817WwBQ
LxNDaMMYbwxcxEjXF3ahrym2uAtgWbGZHYbjTOogoxnYw2e2nqFbm71XNkpm820p
l8ji+DYPsNephVRTldJGlf2gLNfkdxWC9P1r8y+FSxVo644h7THGbcOhaot7UVWQ
/WycN4AmIS5pDssB6dhdhzMZCdw4V0vkBEKxOJWeZDp1m7H51Bh4nob49L7ktSOs
xKqHo0Tqghg7xylTtSJr+Yn6HIHjbtsLyqzrXSyQszDluyUrqt1tVe0aWMS8sZUY
/Dv7ii4p0ssKYtsVTVa2vSOyuy4M2mWKz3vdaf0M9UJ8gYY3yv81xFLlKEjTUULc
uLSEI9YchRSsnvGh6YpMwTM2RZnXKwq/8FIBqJkAMkPwA41x6ixmn9CNjSHJvHxh
sL0A8rA6dTWrCbAtNs5D/Wn3EmnOY+7I3u4x1FjhYrtrKqF8AZT2LZRQUR0tl28l
Luva6GnP5QCeb8RKfFMEevijiEtegi6um0kF20oNl/QEQn9QPQAecqIocEPMbToV
5YS5PmofaSJ4uLQwpaXfBs7h7L+yPuL9S4+qf1IZGOI/cxDQ6y0v1JRGgwRNYBPp
ShkWhHYA3ENiV6VPYE39lufQteOUjymupmlYrWdBK8gFSds7PPgFzC8Y5iNHF3xS
82dF0bQIsima7ksQInCBCdxDi3JuiRKb+ZYFOwW5dLLKtMBa8ySHCM4jLOB1MaOB
IeMufULqk93t2ebeO7vuOfLjOqhVqL9cjjTP7PDBCClqImO3LsRt7Y44MWdUMHzJ
joKv11+Nvh7nN8XnyEJX8BenW/ipPki6knrM6Y5gYRXtnPJv1jtIFtvjjpTcQKFN
IIBKZVs4gceqt54Cuj18OviMJ4H+BtCvNyQVrFL13K1lxp9EZ6JX4T3c7nAquUjf
IAJt4dDSqjOOsrDLRbvXP9YTtCMiE1NCZFoqcIkH2nbKTDVIWcuwxrQSUsZWdWg7
0hJnkApAswR0VEFB7bGP2aGVJZTPVu2pgVbHdNXuzwToZZTNETPD91qJ3BjMx6yS
FyUotbEBddFdgDlZrMilYKPQsJ2yhTQGEaU8hugkenvN/oFm1PsVwL06GN456w9f
XM5mFZvZi0kOQEzUKkc+WVAdgetIwVYcntq7yAapP+hHbhUa7BDY86dGCsjom2AC
chKo9BZ6W9KeG/egwlN33Yl/oNhB19W5xlGKl3V3f2loBRqxXDMUoY3Nabnae6ip
FBp2KQRbo83L5bOEMhpbsK3/j2TL8xQTsGZZzjCfE1ikwTd6nNz6cdSqYGElPIjO
sGhgdr5PY3rlf47b4gdRJN1Ww8r/UyAachnj42wdfQGiT2+ZjjMUt2M9hUHL/b6H
T+hdbrpF/7+L9PWqlhiE2/6tz/9YofnvZSo7tCFI5QHO5/9LW1F6F2OlA7CPDclm
Khh2vJE3xImVq18Hbx9ER2OTw3z0U+upxoYRFf4u1c1PmPjjkZ53z7fFlaZD7ngM
vp0ZIbXQ5t0lp/CjRvhiv/7+W5t3NYXCD3XZD5e5G+E5g1+jX3YgiI3Xw9VuCfY9
lJCOr0UHcF5eAB69mmG5qGBr5rznEmL7toznaefRmWgIfNeuCZQLtIpPaJ5MrIIF
qt1frZTrey8GjHqQ2HQW7JkPxLuMIUbH3WlTucuhC42Bwqb1VdYWnPuT3PaU0Kdw
5ZzaBPXUmQ00BaUQWN/KWFWwkmViK+MONP3B+0dbuhD+NtV9qxOTVITaraouNVOf
HxfcHvo/UyfF071L5GslbYtaxYg4q3mVUq1INkIZwGJLl3noPOY5wRwv9m1kaM8X
1G8kquAIGH63eLmptzvUoJzsiXSEJItvWmGaWA71ptgNibnD1NL/xKCkGzC8sMzl
I1PbzXW+PcdGrT9ZcWfo6hg581x4IjoGyJiKorBCjT18k8BFb+9zrMxukIOo2BAE
O5GA0XoMzkLAliWDbsERffsi9FhsetPwkhDTPwfYJRLYf41IYnkYov6HzAsIYmG1
Ei7kUQVlna7cFjoeeg3rTf9vvU/yBSP+8YK/oDh7Wm8a6ZXwcdfAV8YYbI6IhP7m
uqkuqf5wKHWgA5aToeXc1WJmdXg5IAmKgWvdAR5dbxR3fdjidhr3M0sMAgi0eBws
x1CXQa7aPTVnGr8cpPxgeJ/jiTNR8K5pVuevrXbJFhb5ZKFXoiyrYeOKnxjg1sfX
2zb/oGjEupcfGK6oWcV97mBKhrIYl0hn/CFbLx7556u/Cd6r9gpl2cwxZMM9GIdC
50y5enj3pRGBH7XyXHGm7BjQRQo7U/LU3nFQroa5YRSfwhYU5RtZ42w/Rau+8J6D
45ruSj5xXV7H7/g54u03l0vMTGe6AA7CFtfuHB3P0pfL8lyCXxL8li4Qm0VFr3yG
Pkh3jemSXVh1tXBE4MlKXsgjWOQTwjVr2S7ZT3eC9e0z4bwNnGmk5W/l3DsSzg5g
VoHeQTuqbK6EASn9rEAUDhdbrR3MUBqhqSu4QBYGzkHmkVpgj6GdUJzS0dajPF86
RGOS563dKX++58vL3dKMd4VXX+g5be4t4DchM+EJbOJQbDpj0PGnLNWpbPA5raDq
sv2TvYj+qs6cI9tj8xvs1ePIUcGBlx+7V+Ap28cOSS5DFIq3EAvbqsgNugypS4rs
mw6g+i/7tPmqEyyCwRWbSMBiTpH5LzD47lozv1a/Ftk1D/tmDvpVnDTiHvfQqs07
5jxV9U8/pilzSWbSbujhYQ2wqxK54hD3p7FzfR8gRgYbFJB0yiB/Fc8soR+CNhgn
lOVOoy8nkZFa7pWlz30Jkv29UkKzV79Fe5uK5J7DKa+fjp6TS7E/vfkmaugePWsH
8X06EIQ6rP05K5VbwQOTEHqlSsuxLIIgVcRyMOKFP/NCbmHnEI+E+gOo7vsgAZOo
xyHmEzSCoVn6aYMKEd/yRAo7WE4D/smg09Tjq/HIq7mYfY801iYo5vMZnO1drHQo
HUZhPQUwEdHjQF91/Jk1qfmzFoRYq2WcucrnJy0uC4lKeOfqTKkaNwa0mJq9LrfM
RLUEbLFONtfVLr9FGTagTd+2ahKiOeaZbLyXxbLeq+b6fLAlHVWU32T/7QdTx17y
+nV9B0a6QLtjZWEo2MliDTUc4OS+Ro9fMuRj74kzix3nl0UlBOPgCjN/T73OqElP
7t2B6H75L3S6MQrWtunRjM50O3DJXp8VsjbUJrQCvRMMExST5+Zfqf7s2w/KhR/o
UwYC02zQJbAq91/yzP2feFHdRO7VJnZmJW14ooyok44CIHQYseTndphs0bphhX3v
lJU8N5KQd7YC9+olBNuM9F/fSLF0jq3eP/eaCGAXZtI3MZzBXdQmdhds9bZmghIz
Hb0Opm6txqQRlv+qtkROj18ge8cmtnEkaLrv+ud6bx9dNJ8u4Q8rTn4nmjvtnbUq
ufRIS4bou/Lo+6BhcV3BKENm9IIuEp+fF+K/8iuaL+lxwqq9+kltFmJ6ySXwOZFu
Oquir1ek0Nsa4INEuTUrQg9j+oiHSMZSxYZBaQUspQrpfUCUVEI4HeC5zQh1R8R2
2WvK19wgVF1gWEVs1dYrKdu6EmjAAW+P7YeUmzldm6mZItq9u+droaedOuO1/IT4
evX+rzqOgAeSvgERNjekhkP+qTlAiD5LznfZimVcJu2Xrjl8qV+TRiYzt41Ar6Q+
2GqEO2EnEAbziN7Nx6QWyjBTtJ0gyn7xTPDLdnitt8OjBaGbLxgjyC3bk4Wi8tlo
9ptdy3thuo2fUbjo5DaQdZg67oetlIjJyDp/f/ctdElSspxcRvHVFHiFnyDA/6rE
+Ax0HwQYC/KGXV4377hl8qT31toyFZlbv9CUiXllvOya+GnQ52IGFTezObPvNy7h
vaZ3C38aZpBw+wa/GKDu0NYLp3IGAGsGCKkCUW3Nec9GnWc3PrRlZvLbzbUKk1Sd
eRfwbtRxMxiohCSWnPvWfM7SukIHnd5uknsfxVO5e6EhtvdWCS9PI4DuSCXKrOoa
UYvNEAKxoVUgHWc3fzwRzSOKS5miwwmtllZirmMewtac3MdOPb6tlIe+HRrsP8JQ
wafMMtLYQSQn+CG2nVOb70qCeNmN0goe9LAfquWCkNaFrRGl9V2rccMdncuyut/o
R7QLw8JhsdPteEj+NruSW+qAAp3bHW1uZ/9iltY2o4Dx2jRz07GjDNlyr0+YM0nL
ViiMGSnc2nVFFTbUiOhDC5qK2XSustmV5Kp3RwfH+vnAQz2MFByrValhvn8scb5s
HVwZeKaFhc+YzrIiTd0P5LYDtvPxc8ujtFfdv01HXsD26EvyEJX+ePd999C6+EsU
WLn8u3wbfl/U9KPmIYy+AhaQCC7sucW0vX6E5FWuBzbsBM1euadlGssAWZ7OQISk
8BeXBZmzSCFkHNoi0SAf8MCtfzau0ibKG3ZisYnEkXnYOflyRpCslDa1ud71rdNf
rlFGbFTZ6wiNMpqBCBi8BcE53RC18kpVqO3rSGdYrLwmxLaSvbZzs3GRB4JdpXqo
dtb2CTfS9ekAspfpVBTWtfYnMdub34Pn6BUBiilggL7FBL6DfFT2MNLPKoUrA/9o
dKHlQweRVExVtZdZspZBqO9bYJHDo9nsKOKQJTrsxu2nbCE6+iB2IgKlNIWGxera
JY1Q+FD5PXP9S6iaIMb2fTDhql9zLJXOx4YRs93jhPtvh3ivjP9XRS10XXvfuTHN
CxHEcuEKr0eUmrne7eCHL+ET0AiWUQwOaMqE5GUioWd4cpMT0gvfWAa48CGFicMJ
mqFyj+aFif53tNlUJezJBHDIodmVqA7Ah8lV+enHV0OAnAHajKj25siTkJfi5/SE
GRSoctlNFTy6vwMasKdS9gVKrlmBQozX7dvJQsknMPFMHPBPQESSvmM63iOePK8f
VoCAcxScb6i/Bjnuk60SRrHQ09XkJcnArf7NjaRMuZAk33ElcrRe9nAaVrwLYSue
XxJSkKd2HaUoAH3A6RPfy41Hh5u20BezGjN3bwMCS7p4N8h9Zo4dYbXQniH8rGJH
TudKL2R3VRdjNHjPIwSWTrzZlYOFuPU7amUSrf3sWTV/Ix5FgKwzSWIiREAAzwUb
8IXAiiB3oXugbT8CzdJY9YiFz0PHzqqz/IgmF+556XYroixsVw3I5D+UYFvvBwCo
rtle2DsxRvpcxJdZNf+/eQ1xmCC6BSlN4qOAletWMNZFIodCupIvjHmaeK99t4Ti
YCGgYzIxHeudcfioHJxgQpRL0C/mOl6/9IVZsxKukMUPE6sKNekxduFFjNMCWxUX
D79MsYhVSSwMliSgMnoR+n7f/IWhWGuF0y0LJshvgjFE6IC3Zi3f5d7/aZSFGFxP
2ygDrg//dOp7edgBBbRUDYFZDr+lbsZDbqyEmYh0KalEdOehgrlAjwTS6RZyMWP4
bAbdLJ7JxkCREfKggLofpEPu/nOx8UMCd7X+3XkEtynazgViWGZ71IhbOb4n2mZ4
jpwZpM7QPdwEETjhH9jXe5OauHSfC1rC/5p3/KPsHbbm6lWIvb2S/vgw2iydo01n
BdlBVlX6AQj+8oG3V+ic8w==
`pragma protect end_protected

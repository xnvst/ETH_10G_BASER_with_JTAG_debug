// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:22:32 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WY/dicajalA7rggQsRWjwtK3MyN1eD7kh5eLAIjLmWsLpZJCgEheWiDD024qdZBc
v6WRPjlZgZC//myOWyQ2dqn6rsFekaEI4ZUwsA42ejpLk0SI2UpC0jl+5aGLW1T1
yhvJDh8mwo6Qvt2fNU1sgoKdQoH3xFLdTPHDiLD2UZg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5920)
NVIAmhVCGorV5H9wq317tIJ3nFKZ87hMCpvucX/eDD14PnfzYMRmT/v8enPOxDX1
pv2rVey0u4gWYPTImMLT671RrqEXJpii5bW53j/DnNIbKKJjeO6vDZa0VGoNgRNB
B/Jj69Acyk9qnl9I+JMdNyQvci+mXGK/PEoSgQ/7UZkCU7cfNrlwbArhTqLJQMrp
gcRHdhnKftHAt1PYzRVMJAWSPZt5mYibhT+bXa+AGBrc8vEJDAyBEzoIcng77SS7
q21+eewoo8tAnhe7pb/HEwfXzjneks+4Ncb/6szrpv66G6BU0Sc6rCSkU+1jMVzx
HLY3c428vlzTDfvvt7JwDb6l3BK4NRiHvusH9mD+kS9Si2JGugHI8uGfBTRx2lEN
eLTJbhHBxKZHiqO8TUO5rWPKiiFeR41dl45aYY+QmbzKFOkZ0WNOGFwl44QNzbjg
buLqbwCVutLsFF5vjSbOv6hisfk2E64zxSSPeXuzuD7XrGkj5tplymyJMgphjvz0
vFM/RuN5OkncOqMKMa2cdj6Tw+CpPaFW2csTHXNgOQodRsuZKLdf966kTa3Qgzcj
z8VhudthfaL84eO8R/QXV+EVlN8fO0VAj1Jw4yd+ep8N/rX2M3zzGFdfRRjiTduP
AYiRTlfdIGySdZ5N/2GxUyomSoZQA2bqYK77rm1D2J/4Bfjhx0A47KwviGrxf0wv
MIY0tvkZt82rqfRFYVUzS9srv6wPI1HtH+Zkwdqf0NGrhijL9NInxiCu1OtxhRNQ
WLNNyQG6PrDslspkJHSb3qY7EpoQGcM1iHp5yJR/e5wSpe+nccdrArm6jkitzclm
RhaoZh/v8MhUPO18SfyVDCsMKIcZ/se4rNrUc/MhSSXLT/J7JVyPrZql7G5i4BCg
HwFOV157mkJlA+ju9ED3pofh4uYMZ+06DSm7WGCr8XOVN/fCKsxc3OR0zxXf4z3p
Wf+mzQN/UCF12ulSSzSZ+6Lf5tAztkiYsimNdmLGXfIIZIYecOG4pWn1Zi3jSOKA
NSogTKVZFAEeOKzof35CBEwM/8iyDxAjI2owtXEUeeNIFKdm5UpFgs16w9lOI5o3
qcClcu8puQ+sOftrkt6LnuIn2nBT/bA2Qt1eNcmbYZl8glGrZOqtUkpCceAQ1zyQ
dT/qFEKpjJnKWrhzqKC8fRBRQ+XYvB9h8XbbvAqASmJr5EAdN+ruicG2C9dCpM57
Vr2n8JUtF45GgjhCU4yfcxvxE8mjnUAVbw8h4Ip5QT72C9pkfP/BL+4uhZ9ao9b1
f7UNC4SwVQ+NVkxuXIncspx8RLkkfSc+Y8aZHad07K2IINqkQjjwNFw67jOM/TOP
jNVqwqLqK8iM1OBVaHrsVKgqtINIsNC2qB9dqmkHs97YW2Dj/IJSXkFZUU4Kq/WR
ww6YEe+PznucukrhNmlsZtCrmpk2/Yv8iZM7/TpNo/+koGtW2arb2yRtBb3g3MHe
ekUSpxCxl950e7uOjxYIIkUy9zgHdcLlxZvcDCI2yNYuHsvxKS19SnIk7XOv/Wof
3cLPBaYdnO36x2aQBA2rvo43kjgj8gEAd33/gQtm3HgsauINzbCdSxz1b8sv85fT
pIZ8gcqs+SV1YbKSwpV7kRDc+/1mWI0fOu6uoGs4y/0wc+pOH1pBWerKSG49812l
I1NuJ0mOAXnLsrobIdZhlmepfiXJdAlhOuz4wF9BMr4xK2dU2L39pxz/YhMPzV8f
ixtObwg49tTUx7R9Av44Ly/XePT5uKvOO2KjuCQUMcsnS0xJ7Xu1xLgX8Hyiz9b4
wtYEWQToKt+APDi/P+3CCUmxADi8GKIBCU54DMX7dZAiwjMe9HkgFDUKlXTF5QUY
0bXzzerJQ49E96ovzqxxyxF54zBJj6erTsUJtcLnr/2tkAWhyi9HlyKRVx1/j7I2
vQ0zdT/udwGocxS6P8H7m+K+CY9QbCqDiMTwKajr2/+cqZbypqM1qxWRG3gWKBTH
N4fa9XSyHfNakDJ1HFGdcQXqtUB404IS4/ftz9Sq/8FuIEgqYMnY29A/eQA0oSrM
b936cP64PyS6DfR5UucaetOxF4sZLLilNVdqS43K7AGsPyWlPDwufT9i40rIgWIl
2jWQIHoFIskH0hfvLn6XDa/3mn5PzSW367bNlObU6Gia87Ar8VMKA8f0mwjI4Dqd
baVtW1e0N9NqeZjT9/Y4bVs9PQncGWpMErIAN6/zL+1JzOv+gTMa2CjPNBWP/y1F
1rksalJsOmpfLBh92I6/L86Qmbn57NbZ+tvseu2NDn3l0rBwbQAMIBvY0OHn0IDA
7rvpCWNyvuipr0QGAJL3dhzA80fl0RcX89uLdIulqo3sS/rQLZFRyocRAApP5k68
NuREt/gzadnQpHtQTMB0pEpWT9Xf2tYqSfZEwd/zZfNHMBSpWxQajzymGdFv594l
jtqU9juxPI5yYeYbleMd5yg6nL1h38m5FHNfRP9p0xgl9Glasfs/bPAIv1Ql8H+p
Ttj6B1Vq302KLo/WvrB68tNJVAfff7W/sAzLu8f8YP337I1O7opjpweNIF3AXxca
RHkMGfXEODpOLprHe50buuZTmKUkUjyYrFY1M73oDhGX3mgM0ay49jd5xtV4EaCX
kFJQPpRYh9BWJ06MBlBEwDUsG8pIBYvf6iGBEVHI+n6eqVb5xnuuW+sicXAhBEeY
T8YyZOLMPs3wMJbfj65n0xeUj6zGUmmZW2R3VdWJZJt6UV1xfgeOWQIHGt5lErtc
Fdqx5TL6Xt/gYqqGI/BsnCM03dRltEkdH4dDHVtmMOegd2HgT6+1EW41jyGULj5A
ETu0n7qTzSGwKMiv5qqI0NSCkhSq/HH5GUXCArU8swTdRqdAsEIzRNKzIluGsf2Q
0JqtVSorEuOzudl6SixN17F06E2aeDWRpQ4B/SzIf2SjCBMdLOeQD2C35irX+b7u
V7Xp3KFe37z6gXA2aLtEPzXXVDd52JJfZawbniRTJsrYBAvbc4uMCyADdfBSCfSD
QYopLIwMYEVuV/u5NrmW/SMFGDZKGdnh2uRnBrJI2Twe3E9a0M7Se6cZUYwItDIM
vIFKcjC4OXG8czdS+x2I4eO3urwBwHRGP0hvwenpoZlivVtVYlf3Dn5ITYcmEFGF
KuIpbJR3i75NAcY332CaWqdYOfFwlBgfxVcAEtuG5OKPn59Yxuq5q/Muhq4vvp3V
7cOSIBpMoSLpuX1HtGIpyGF9bes5GicMLUbIxsnrP+LAVCO/lYi0ZEYjnxnZi/gG
FR0YRPGCMqwLDgFmzyfqgx7rEOIpwV8N0m9YjRjzqVTSumiTZDUnQFIb7WNPwTic
hxtlWrxXaX1GhJjaWd12a3CngehH9IaQhk412Xq1E+3U3DUKNIifUo6sDFoT/6Pv
Dp92y/uWtOgsRJHDr7dq7/TG60VjfJRGb/AFMgEUZq1OYsdQbHOfGBb6MxUqQCwz
Tzf1ei2BZm79wYTwGwlpOBBGSrgWfmbqOFSZTVMQfbfnrSOu0BgHOL2ymujSaS6r
jaOB2UZfKV5bz58rGVECHrWZ5SmNUkH0gulTf98sVNgLK7GXtZj8AYzGQEkgvoP1
FwXOt2iOBVJqCqa9qRdWcHvycQWB7mM9UqytM9wTpDOisTOd70zln72i+Pi7dwab
UO8lvPOexu+0F/L+fjCqMkwoY43MhjPMb6Rj2QFivmOf9kc/B+Ai4BZ1pg7d6AUm
EE455GNfl9EhLbxOXCECDeYwLVNQOAg9ry0nTBq4uyG8jzKQIQeztiKm1zcWn13+
qWY3YarR49mflEhYz9zZml+wsjQ3BRdPCdVLLAG00X7oFj4A1FMr/30vvUGKKr9l
jjHkw3oIY9VORpjiMzGWntuxSsMnLRfO0zPD1p5CtgWq+11ytm2RJXQMb+mBIwcL
dOrhBvVK+vR+R0xxarzA5ewMRLkK9BJxziUqBSU1gj70/NwTgMVH8kdtH0nbulut
kDfaCMzKwEYK368VRXsPwbVYrkRhzHGeo/ABI81FiNSzDMaNm/28pU911eRXsAXD
NZkQid1WWr2dglwM7Kb4Tn7RFi/J0g/LfpwMBH/qQt6BlE4gMPfNjL7m8UoIXh54
fk67aLIy0LxCOQsBMsd7rV871/yUMT3chnfvk+BYck8vIGqwD0D5NoGRFqP9Ssru
TFuZOybpEYtv62lpIhSO2BB4Bjehjz3jwn1TC+vgTtPcYo07zf7oCS0MLDoQEXUQ
1LfNtg1L/FZ67k+6py/VvSyD+Udv1ZvePsX/sHJ3z9hX7oa9aMga5lsyA2qDogBD
iIc3mMsKlAXZ/kq1VTNZGRHTjdssMRAWN+3r0mnoJeDPFaOTKaE1Jy8j1YE3zWAL
+yjhrPhxbww+fyntxKFRLujVwkIquupEIHmEg0rk/kPjwd7ETWeIIUfXm+V30LzH
ycNUeeVWu+Vom9eZTU6ij/t+GsifKV1tUdWHwQjFFMuG9G727D5kHFwL2AfvRd7r
F0VEciRLcqIl9JDc9mGzAia2ASoORanR8BAb805biEoxcZy3JMlr43WUth6S4So1
c9tjLMMkVA+R9du3myKypJ2/Rj6szlwQjkpLoe7V9PacBWCdPcLCeBWmgkELf9f/
/QIxbqyh4NZd+UKY1y8DE35iYRMZMB9ffvF11qM27JjRVdAP4Jne0TVUJXODToFB
hl1SXROURZXRpOqvNMnoI3stgnw5Ejm83SyIXpq//0qlqgzeqM3BWe1AN2HqdB3g
mIklf9NAu2Z7FJ4IyegccF2JWDind+559O+tKZmaJG1Z5dJP9y78MddKN+3Vu9U3
ObpaPrWdgM33QCM+0/uPfGn1kIYNX8JO0A9LjFx5CyRjDzEZfnHEfXCo4fZ5ANAU
nrzaItVvHCltew+IvI8QsXzoKynBhyCp56Zd1bb9G1KAaP2ru5Iq6Y0/yB8EeZf7
jCJEwvQGyYVJqfKyIdtnhKmEV3mIgejG/Bb//E/9FMSJOp1KN5alQCCw4N2uLSxu
6D/240jFcGcEp4HRXcyQPDPx7waqMzBXGkvvihMCjJpv3ZyfZdI9Pv++rQ/PkNoP
+I/ZgxRDnnOy8/hgt6jkiuyyL1DcQ4LFxNMW3HrlE6jy0E8w9aBjLV0R0GsCLlC/
/bQ7V3bWaGAPZS6E8iPAV2YYUJM6YOA3zaKgQtkadw18dcaCT5pdRTEohHU5FdVt
QfjmlyQ/GBDUfSNg5gB0rfOoxf8WLcCvu0XBgKTSGlBMe4B60HT0mJXn8upLXZPP
4uWHWWTw0Vlpll3yS380zyvLc5Ub1Ern0QTCD82jzDyoVXPzp8aKKls2wWql4ket
0qYlvQ8HYzyH98zGzDPzlPGnYmZmwTIOjkjnLM9XbBmyRREfiXVj8lZmxLXRGiHp
DHXuavQBYOFYI2NbS7r0jNNobiKLut35qFVZlsj8480ukckd3Tkwy/MyfzmUgBjm
/aPCQrIfp2fkJfXTkgRvs2mzCm6hyAn4cBC2OW5hzKWZYs2WxUGkK+Zie5YcvLSv
ZQIWjkFDgbP3QDgFpQ+acLKpwTmGQoXU6ggUXLTlxCzFa1kaJhdrBrMNo3DbmrOc
t9wMhfcyacRl4+2qADHt++GN6iy14S2i6fv7i33SLZGuaLg9g4DktPl3s2/Ddj7u
eQ9KUjcYBLO/g8PxX5sOClqupjnw1gBY2uiiRWNQfpQmOU4NY1zaFbduXeJiXJaA
mpSnIFA2eif7hvVynw4x+OAiVqN3A0sGg7thTgE9D+7f9ym6RPs6oyYNz+pagjpD
M8mZTK0pZi+qTjWeJx6BGBiqrMF6H1w4ENsAxABNg605B2PhsQxF/X0AGF13PBMG
oc7SHQT8CRPzJC8JtTihKawrhzjovIslJg7dSgmq0KKWKb41tk2AQzVYLop2jhBA
nhbVvCcCXKoqTFQZcL/C2ReYmEvdjlGFuqQ/+xdGLkZLyXZIR0oCdURTlEX46v8r
lKw7aLX5GyI3jR7it//oK8TN5YrDFRO0kBJVjPU6AhROX7Ml9bM751R/k2Y8GHgU
3eieP6tBBmhoufTYRMvJ6IAZiCmcACiB6gn5d60yDAcT/KRgIqTR0piDGAzMsb3R
YuE8Dsd9L5/sRK+r8ex0LFMi7c46EW9Pey3XFLoPISytVqBo7zaqj+07jO/JFiOa
06jGcH5vr+lSjjGgytXTaAUxyabX7irJJZXK389+UrWVDcAHmorqPMtGV/m6pvm8
jug1NZWjhIRpv4kJbDdBR+MB3auBR7s4pEmBQMWVWZWR3H9yEzQKTtzHfqvm8RAw
PzXtFQdsIaqwUY1qDhEMew2ThU6ruSBA0o6x48ux+UXmod0dPpId9ytszkxFTF4n
N9Jjl6zg+JDzq5tZDOBGaVnQ68T8oUDEnF5S0VMEu1JFZrZpgws8dq6FkAEQI9E6
3vEA0CkgIKpaxM4g/Q/+f1VtfS5FX770dSm6P8Pw9MJG1R5sY7cuYnsltNYtEN7e
hk+HIadRfLU1hBLsbR3DuQyQkCTPfo58hYY5YyOvf1TUYkWnRJpUY7ezzUI3bfoj
XEhhN0ZAnrEzShrmPo3NZN5UssxgGQV33ncYWut9SN1dFi87u7Ie+8Oz2U++7ptO
d8Wa/mZltLT8DH5zXAhzCF6nLvwlR+v5Jds7hx00E2E0LnjG9PayFR+YIzEAW51W
jo7K9ZFU7p/YEYOZ9fhjhBaxu1C7Uzk1s3wXJfCqzLkhR+Cqcjc5nILcwYfyr6Ac
8CKD2xSnKVYzP0+DWvLD8Pf7+cz9K+KBHvEiuBa8gOlj7Sclbq/yBlnt3oSy1ppN
ZY2Ule3v1qr0Tc4LDBDXu3xQhtKowHaY4m+uok142TlBhHCGzL6TP+SQfo6vbLEt
0HujTHxPZveUvK48AwvKBfjey6drY9efF/rkyUCLb13YVkqZOQ5pSAKolTHvHUDD
uvPxaM2QxjOzywbAd0HMYmgxz9bJUbSbqiT/+mJL8sw7t6hqoZmHYYWXYvmLFy+p
f4tthAQMksz42+GADG3u1RUnPH3cUq9E9cOHfLiL50SSYddsXoqQ18jtkV00Q52y
PDlfGmc9sSdYclapXbPoHwneEipyeo97D8blMTWTrMyZHULf5MdijeVJEC6pkTvC
icq/j1WTxovHayxtPOgjrH+wl9dqlLOCzvbTY+EqgLWi8LvMb0bwwYTFSbxp4M8c
L7IENZ1sx/rkMVjsgE1IgyrNGEYXGk5YggP37LWLjHX6pu7RlhEHUhAAfziJqK+f
IvHfSMIM84L0UwCBoJWxGSq+gHlyG6njrEXF4O0X0rB83MT77TaJmdSZBfpaOT8E
yFdJ53D65rqV4KCZWpARIbC95HAj1BioLX0eEvih98KeZzICJhD4N/APY2PnT7SS
Z52ztOuZda1TwllkUIUIAb+dqCAWKauoXQMokZxJQ8aN9KWiTrCbzHyRgv1UFO3c
nNA7P32k004IA2llj/ObQcxr1Y4vJXg/NQyMMYxAxPfLyjTcBYJdLHS4IuXaesII
exKVa8va/44oVWj40Y7UQHTmPxosbhBUSr95w9/d4/LqYa9sml56DsHICIg3jAmk
I6o/Gom1dl1LEVDtStndpI5lKynbaiOjTP/yCsl/yjXC54v4gKsadc0P9Uk1XI6J
XSAIrxwnLLB6RLP2qX1xunVLA5koW9uMl2guMAhw7FW8/z77W49ipFjHwTTolwDn
4SQEljx22kYjVutP/LO2kFwJpvjdn2nEET9FGRpEhNStildmQ6X4jVmiB295d6eo
yFGxFAX6paySSF0c0070K46fZ2Hl9VB/TYx2sNg6faLtV0FbFWyll9np0e6XkaN6
DAO5Ao+yr87CHq9fIwZou9PxI0vOy6OqufQNk5dMs3dRknLPNwZdjqarCcgJlwZK
y++PbSKvqPKqrhBbunAIYw==
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:23:15 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WO3pnkHWkm61Bw5fbLo4jjO7PYCU4fZjdVuLrl3/G8YrupgTRp+7CzYeiE0d9i4U
7KbYx1uw68VpvirDR038p/h3w+VMRa6kppnxYEAOYTT3iwBBBrd3nCYVbOa6ejww
fnbWov8D5VXI5cH34cQT9EiJODENnw+UbMo+EPCA96E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
ZensGgjokyweuiBZuxaodYoTARl/f1i+yq8mznMqnEDov9QxrZuYGkNmaDu8jRt8
FW8B1/GbV3W8zGtMaXrNCi6zxQrMPRQ6gdKW+vgb21RkvRwGxzWq+mfeRlZ3Id9v
H6ottgWGcJeqONMIYy6X0f1TrCO+HZwib90Mh3Tb2oCEGxEU2Kn9ezBRXe9I+Z5V
1wZKkGqIJHEJ6NoKnGSnK4L0JdSeRUf+TjEwx8y69Ne8fDEHyn+8YhYit4uQyvyb
GuG4OKULpK95XVc5jN38bH15aMGuNPsIAK+1uJAmkNHmzp5yReCOKWbNy/E6GxUw
Wpf/bcz6lyN4GVI+tb40zt8GMZSH1ag03GHbWp2VhStEh7/kdDeDF0KML3RuNALi
KgyG1bAN2JJU2p72o0U5pY9+d52RvA1/NE7XX/eFru6OiaLVXqEJ4ovBsELvftGY
QquZXz5CUYFmnK5kN/LEQvTtQAgSrWJTtCsrenDIfHEiMDxREWtmu1U9DA4RXURv
BqVPqlrArMSVaWNwV8ZPVGJgjPzPO3xQyEqtjRz6Nho7c0skV0PuXTqFbyqvB4iF
TLvJU9HgBwZKwbro0tzapVGRd8P4UN25QO2aU1QkGdXmVYS+GBOyaM/xye8uaeLX
scJdADMqvTcETcpAg9ruQqeJ3TDosT5Jiq6g6MByFY1+606xYr0BJNOHfXrWuy4m
gc1L5VWqcuTif3HJix0jPYwxq6i5zDHFo0LPlFKJee5w5/8Axvdbf9cw+hI4/fON
4DBLsf40CryJbazF9ofaVCWHS/tVyBKYguR2VgweTnsNUNIaEolCJvBmLVN1QUgO
KYOEcQJynylz/3zXsHKTJBUE91FnYWrLhPNexBx+91TsBzJ86cD2TG+OnYed1QW4
6UK9oS5hiWLrO5+ZjMg/DPZ9YB+rsineSGX7hggeSv+/4DyLD44Un6YfBSy832VP
HM9eayN4m13QH4U9Zzc6ito1mRMixGml3vJ4AMDxIweYhe2kLkDuUd4wxeOcpDLG
fKt+MHj2RJXq9gCgm4FRLPZH7bFWitiSoGob2I+PCYBLsIW4C6JiHtAFZHpoGyuP
yrjUOUIBtWM0uqRu4s6fKDfVzcqJInKUefukI6UBfIy7m+wHFB8niLmztu7++tZ0
REEzFd21FQh3nGk5W0SmvRQbScEvE8SCQBprIPXwPDKMcQAmqMVRtW4N3MZRS0gE
SUi2zb1k+RkOrgqBokKMLcVNsxL6lrQO0j7xkPU/rZrYp2sOhZSnZeyLWbkW6pGj
axGk+jzTFv0bTJbotAduTJLn392+QmK+OkwM/1OZo6XS1Hqj+bWGiWgs1b1DHz4h
i/dcE9Sc+bTjN4TjftmHl/Z/pTdxwxnCUxhyMkPmZ2abB0SpMcUbivND9XT7losz
tYv5H3gTDro6r4/gDDwIho1xOyUpXw1jy2Kxdbf7/kH0234QN8Enz6aAmbnXDWGk
NKu1eji7otV0U0ZM8pYfONQx+NA5CMeAT8ISFSjesDDktKxjkQ9exhU/5dZ7dgzE
7stKYr7KPEhdAzvJv7U0Xf3+iy5ugg43iiVqoMrdiF3g7ijfrBdxmVJ6oth3CXdX
3p9N9MldZ2Q1GCrAPLcCIqNNK9MVSox0no1ecJXdW5zSCxYFeDz6t/BczbvpYCPA
fE1EUxxqoZPF57jylx7d5oO/qTtewZ/rIRQv4oJ+ea0xqt3EM9yZoJe9mnHK+Fkl
jAvF+VzeGnKDV8KJNMf7Vi4wcGkR1Qvn46bkHhGt2THFu+iChAWl+09OjEMh7oWR
FNLplEycLkilge/mrUBLeKbuBCl2pKaBX5QaQv0qXuG9TfxdnTOrNBwYrsQwSwj9
XgMBJJm/BUOy66hVr/JN1XR5bMUAO7WkWlnxLkLX/hyRIVon3JRNklfO4AT5eohi
Qe9hhG8haVdInaHJUeBUVR+NBzYtUr6NCGUb3ITO/S11o/Zs0T7oSkw0Fp6rE1hA
a023bCHxyW5ZknQR0LNoNW9tzME3mFpMiVKdMvpm1C2KfiImuK3XU3OJoBjGIVJ8
Qwrxn4OPSfgnhMJFMaupeTgzB0RaRFDvApPauNpH/LbbA5FJLifC4wRJ77O/hiHn
wpaqQs+LJtS415aYrYrKTAkjaZVZXqBjywY8LdL8E3Axjcr/JjFLe2L8d/T02BHk
ErGNWQd8yWdJhaI1zTTWf/HzkbU1zROwT+e8ngBd+HOeecx2XD/XeCXkp15kDBsQ
DIhYEvkZoOJYZBqS5KkJg3unn0NdhANQis/fhGjXygNc2RbdfKup0lQrhJRlhlQq
8czfcJe2SBdTPDs7OXj+kr+cdf0AtqzHWTE7FtMAUCgLqQiuwJDq6DHAVPcQVDre
Oe/GiKTKFb8B3JRttqUDZgr7q38vWWRFQldSBMGrHbJmf6M5bVlLM71NCePsl1qM
zqnXYFzr+NjjjnCEzq/iJ0zcaPbj+DB/pGcRgz8YtdhfCyG1OvOKzAmhJMTcc/hD
20JuGfnADDVhyN8N1xXgL9qtn6xxAGiRbliwfp0I5ZUv9CbU9J4zvsBvQA3EVOGd
7Z7Vpl/XrDC3CRaopMRd0En7W44m41bmUZ6aQZLmzN+OgQx6qwBTQwOhTMFI1agr
V2MVSbuVfacXJuorF3NiKGQOtTCqGdIE9s6kaEvPjsmmja9mEyCp/u0JIXCUMKEQ
bwbWEU6VTq1U7AGZ8BmFZ8Bu9+ikB2iVtWTioBQihoBupJ5ICxscdGeq9ek6EpwV
p8HbXqz4wuUc/EJlTgeO59UnbuuYJfIe3b5ZvUbzgNHAlAmddAoK2ZTfR0XHJW7q
VdfORNdjdikvf6uHERABX3xP2E/jTjXlKU+XD/1Fx5GMyE6MYXO4HUOuTfyQCRbQ
/ewETWfRjVhw2Sx2HJkcL71i4SA4A2e5zQ+l8R2qk1/MTZZkfZVNmKRm91BHlOKf
HQfcuzylBMWuvKBRo6QBOECc1fi+UGBivR3j86pilH34wnjLanUkAz/ytDXJKJc4
Vt2a2h5TemM2J1Yp0njMDgBSEqI5STUl7lJzU1aHWaqyzJM7VCDIjH1nA2qcg/7D
mtQfNS4TLhsHI1YbXTG+266i0AAE29VRUjUBcHs/vxltlR83LIKH1mYw0F6MHrgz
8Dpwg62wUyms127710Jwu6P575n4Pmd4/eR5SL2sxHtN9P5oVTRZwa2w0dlXQ2xW
44cz9ZXwPYq9ccL5U1f4RWysYGrYC3Q6y58ulRMC1GGg6QxdKzQ4cBhvPbT4OWNE
rdDos+TqfqriwqHoJLcAmxHy5P4nGwxmcW7SOkf9/lobrAhlV6i38Oxs1tfg4aaM
bS6cpsgWC/cZ7nCCQYU9HN40pybnJnGuBV1hiNYw4z589iqnER3xPhwaq9C12KQb
bdA+0KP4E6NM4WvsbCxlDcN0AoolwpXdLdxw2XEBLdyaZR9MBPw7tk+TvjMl2rX1
aS9F/4Rwo7pNcFf1SIu16kyr7jpe4f2qXmeypmM4ZnwOExkgZcV4TUQ13g5u8K3B
NluGPHGlndqomI1nUFtylF0meu2CZGtpd3cUKCSrCa8W0m3my3cXHf+S4BZVqMgB
9Fj/iE9QvnxYB2ZTSg2wmMuX5rBbZMZgtaqbFzZfaJ4LVrE0EtvW0W0tLvLcT9Do
PkYPN48O5zKCyjR5UcEoa6l7ViwWk+58Oe87vq4oHFfI0+IyD025RXXCl2wsGmNF
uDRLH/ve46QYjyB2OAiV0lLSs0tRlpK+j1BtekInYl3a1bg1GzL6m5ll1AoW1Gpv
mYkbYVLVU+YkwdbP079+levC6AtNWe+Ak2E25SRBCfV7SHv5PEaLJY4b8u3Z0Sf+
JVNPynhFooFbeQ2srOIZJzl+T4shdIGrfPz3d43QsvOtL4Yv7mVVsT8JuDSPihYr
z/dmjpbVEjKtL3bdGDGLGFpLQs3nVoNNh73n6dtgdx7YkPg0XefhV4ExVUeCBHcT
AvWg8B09aE3+rTpxJ3uYkTMsst8o9fT0iYQQa9QYWWmvMpBRusuSAvHDOuBS6haE
nql3BI4k0OdZIYBECXTyfZtGeztAG8Lc350Kw1fs25PqBjMJuWIF8GDBuqM8lwGD
oKKKOwc5chy2FuLxibXOuieYUGKQ8dahQwJwe1jSL9PuJZ9nsptV78DTQ4DlYain
IaK/h2ZcxvpViNmPc3BTMyAHsHbBp9pTec0xnxQssmdZ7fQ4Q7YT6dTnIKWW5lRM
BuMM862OAiEB7dml9cc0tlnKeHHidSBa4RlwqMs28thWaToDdusbXc644YA7AQ4F
zUvdTO9jt8KtjUkMz/Tf/oh8DN93Mvpfok/sLPC9ME0JfyP1K2pyI0TAjQyhzQ48
tl2Nw+qNnIzvKdvWbzATvah3WiTHwdmuX9BebDV+gl7dFDZTEC/xAA+FSbYeNV6Z
7adgBOeVdNDRQ/qBvUtGL7WEppo5L5ZLJt5WgizRKwL9dKbP5Smr1tnfKCVMmTf+
8hqA5fSjhFlmEpD6LoWmiGCsuv0oeuDM5k5PT9P9mSqKMydJbIgzY9ldIrPV7BLz
v+pi1RIog1U2OYzZ/VIwCQ08tAjw9fwkwX4b6Ch2JdOV6M648yz8H52UHyoXXJoo
3lpUqa3zr7CkMbZYppKtYNGEMqIfONflmasfWwR8CdeGYUtZGCAaD4tNKQW4Ir7P
1SpQEBSfTAMlC53hFbJoj3MaWky1Mw/FjJ3oPX1p1bRkRLziQ61fzcVojzudx8+k
w+/KffqcorM2JWYggNFQNhdVlYeWzdQinYd1lVhl03c4u3qr1v+xEd0djbfIdZBO
kLXxz4Qyj1UtQLcGC1XDyQy/KpsDNbDIGMjRDF/w0biZ8xuFHK7HvPmkzS/Xef9c
WcpOkaicIQjpDiHuyst/MuLG2AF8d/uG4XQ6aaiafEUlchiGHuNPsvIy+92weQjh
k7MHlrR+Kf/96iXjUt2q4aBtCQkLPP/bbB/z6wMVdIl2RNrzWoueg0iXuPIBFWmP
5p7kR5H7Akl+wvW9v/dgBorCb6zwvQacV7r0GHOECFQIPXmqIcYG/F+7O/zEZb/E
o5XxWMph7ES5opCTjR+JBfNx4AKTAFrGkakhsCzSySFz6x4b7HasYUj22iHiuIT+
Za4opUDgVnxTBvVJs04+S62Mu8T/hTO9lNcChU7tjpGXARRBw6lOZUz1dp3WgjWp
pC8h5OzlIQDgl/OjoxXqrCWdCJSkWG+dl6GPgZAEMVwEwhfKhA21J7hJP1LFrGLP
HrYrsuRLdglt3v0kwZRswFBdc27Q/qFaS7D9bcgtMlFHAEw+bKQVdaFDmCJYGJJO
7Bgvz4eAa3/jxLp1/dsTGxqrJxN7j33GGyyxMew/GmJR3BDLsZo5kfrJjKlaczMr
74kuD4fZqv6mOngWe/s1VV5/WfzqPw6zY9k4vl0lb5SytD5+mccN40tDZsVcbVXt
NCtJm1JjNDd8CF3+Ds0gK/drSK2333d09Apa0fy0duL4wXu5Hka1MGhF2D4tArzy
3kSVi1itEAxrl166lLVFS9mCgvVyVrEfixH+e/BDJ0wHjDQc7QZgApZBYMynoQnh
CaH+hFvT2H4CH/JHNU6TDb48eiS3OFzeMD9bzgEGP78bHYXpi8LFGKnMD/IQaT+U
+4PQYAbudV5WXqtKYM2i+OLoc0e6filkEdx/yTqEDzzatm1HSh5NYgSr5QIteAsI
iNful08TF2KWo9ZXIce1z7OjktgtnTjeCH+C7n09pBR5ovAkMuQAC5r9L9jdpEj/
xGLviY5hAm6mcXXHRnjddgqrVsrkhzppinjPGld/P1Wn4XjDuDDanbaSlBGRw1bj
OT7dZtynMTaC8edmKCxdZ/NjccFXkMyo9ytC0+ars9SVqgLbSxIVC4Tc6DiYRYUx
nML8kZR8H9YfGIAjZ1xbbYJ4cn/yilEvCISVkkIeDXiyiGv94zqebQj+CreTSTAb
ZfDm6NgI2IHxxKT7A1DrFF13IIqDFhvry2ds5biwVztGfuXbeXov1SJP2fX86UHC
uhoa0vUSWo3qACU7GLLLF1EKd65/ZGHKb3ds/QEL/jnEpdy3ksHYSBuVaK4Z4aNJ
9W1IJFRjPHmbYYFyfpLuEPKkn6FQB8p4ZCtlP798Q6g89bAnyJ+iJJfXRvxIOaxm
OZS3fXJxE2ajpePz4RD5QGArlxza4riqYQic+tnRyqdkMRQf96B4gI9bHw2UCPsK
3M6P1r8DuDLbb6hPKWgutj1J2V81eSjriHWjCaueZr47HNBkm5axefjQzzNyzFOg
II9yIr4fWg2NQc2ILwqKRG+/7qqMSEALtcyQDYjDz/KnCCL61goc/pAC4Jvx+EwC
NyN59nBfo2i+7Kjaxinqvmhfwpfu+RbV0yRb2hYNcmMRZ4kgSIjEcUWIcNeOBp4O
9WaSzOjxsd4IJYXp2CznTaRA2TNWv2+eVuaw8enShrURcR3gNZNrIp/YqTRjsv9x
Pd4oiQHqPR05i4VISFJVOuvb82UuVnpfHLnGGdGBxWZJrEFwDjWuXqEoYL2iDTYS
JXgZc1QcFIDupZaiHBdPKBZVfuul9E2ShgDi8K9vVYF7rnFY4BeUeG7Wne2NwpL0
8pr9hMsR45XYvT+vNOtV1IcCbaprHg6HawX9KSOfPzAvY3C3WFIn6xqWKtu8fN1x
T6RxXn4lqniwtwDTLOVrKCtYEAbYyYOd1znD2yYt2PH+l9IZ6htbxh+Lawg0PLlE
rjOJt9T0EodlSQn/G26npXIAmT2ExG6rrU6nBCocPDc5Y9TToueFYgC605yCj9ZE
lymnOPl6Cu3dsmUaMbQHWgD9qE8YgmcXCfl5fLsDJBOE5B0L33B53oUoQwfBNvha
hCPC1tYdSyuboCIcCs4cPujE71WWxddjprebaZ163UURYLdpoaJ5jtbXDnpoA05t
8sW2iWC+hRXn5xii9zj5DLtkOOE4nhEXYLi24Zu3QDHS66c9q0t1q03+hTEAm5+F
JM12UtAZx3Nl7zuoIF5Cmx3WbjOEao1H+c74KujMQKtuX6FfJQx5VeMGKOReakL2
mZH1zpu57b5wA/O7doKtI7b8+xoCCGk4RB9f7Os45GFZxybqcWcaNU6MJAgiiRb7
PCl2oI5WRDPYZqTqcCMccaDNIffhzXzHzFziCZAvgmOVA3h0JPKZyT1oMfh/Mn05
rJF9tXzHIwpA5CyADm9TzKgD29Ose/phIgzcAGpVxH73X/wRVf4jiC4FmP2ACGPo
2yZFEI9vMU571e0XvXm/vYhGhAuHh3jh3/cmw0IJW+pVogunbuUt982rVmQNtSaG
1Nblos6RbDeoiQBFkaP8LVOZhaq3E6keIMC266hDKuywXUkE9W9eUL/2iKLLbKAL
sgt5W5u64It6vLDMBTE1iVabjhVY4Zhao3jNYKXqxVcqu5dVEkQHv+hREBCv7boO
lYwiXzFr47DG6NrKjJmCaMKDIzUhtfAj5KPjVxXfiS1IbApuDyAfIdz6+i6NRtoh
w7jVdwYessspmmxi4Jauq6lIrwRGDGzW2sQjauh1LdnQIWIVhXMJQZFHQUyuDy/9
5pszvDOyQsIMuYlYercQm7KSSSraA6gvbzMIjsx79Zw=
`pragma protect end_protected

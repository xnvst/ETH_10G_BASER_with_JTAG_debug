��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO���(�
!�ܺ�Y`�4�N�;M�d�a�B�d~��xQy�Ө8Q=m
��f�u~��h9���.s�8u�x}Rm;�9o���X9 �T���燷ݠsj��U�����.�應�Cq3]2<�]43� ��^q��5~X�Y�3��m �6�yە<⮣��œ �Cg��V�|Z�f��6`����Wg��D�,e�u;�u[�4�i��r�i&t����*��(�Ի����d��Γ��E��c��)t�����}��:�f�I�iΉ��:-��L�3��:bF��\*���Ce9JK����(��*�1m�\��~�T7Ɨ�s�x���kco5ɠ�Ë~V�e���l0>�PE�ҭ��a��lT�>T*a��ܩW�G�L�l�E��l�y�;V*����?¬=]�}��N�X6����=/M��sy��ȟK�kB�X�75�~���)�b�����Ud��〹t�9��JiǕJ���X���A��T��!���8񒤉'�p��w�a����N����3���f���ͦPJ��E�	P��'\bb�a:>muٰѬ)4���/x+�%�OO�zV� �_��VE�j9�,�\^69���Y�%Y���B�ϤT�(�!L�6�����D9sVE���=]wƎ�����?���!����ha��sn���3�ih�a�\��[+�4Fk�$��t)Q��q��TR̴���@M_^�s��_>�*�u7,�B#�#ΰ��)T��{c߬�T�U����)a<ۻ��yC�(@�AѢVP,��0�Ԅw�c*�W|zyk�q�D��G�6�BRہ�|M��;�P+�X۸S�K�:�v���D�;}[�ϣ���(P�\�Și���998���L���>:
)(���<,*-qkU��M�2�J��#�;rŚ(�`|/����W�I�V���D�Lo�խu�s�6���E"�5y���8���鳽��+�5�-c�O g]���Dp:HJ��+6��_����v$�a�߬}�n��6�F����$h8Q]Jxrq�˪����ܴl2%���H�?�,�0��.O�eǈ�ar
,��3l���6� e��7�����e︭�F١�^����_WG�Ʋɿ���U�ڕ7}ۮ�M6[��0C�?�Ee`�wе�@��m:�>��ot�`���C9SXR'�%�;�R��rd�c٢Tj{-Pv
�����\\�N3��ky:���e���|���h���}d�H%����Er�J���my[�Ǜ�P=ͽ�}V�5������Tՙ��K���l� ~�oa� �.Z���4t��5�"@R]�v,���%{K�,GF�
�ߴ��`H觭i�U�~��43�|h�p<��WF��vђ�Qw�����g�i&��0T���ȿ�%�0Z`]��L���8k�{������T���3�?��͐���;� h�	Ǭ���GjX���<#����JTR{N�!]~�����b%�0��
$)CD\>�����;*�W�M�����(��$7&|/gJ��*h����.<o�t�J��[ߙ��u�~���1N�#Gm��զ�ӡ�ni8���,�N;P����t:��[U�z�[���"a��qaW{��=M������-(��p^��0F��j"��y��ۘTF�������G�;�Jc'�K�(�`�Y�NV่Z�!�ȶ�� ���Xȑ	K1�fy��<���Eϩ�O<n8[/�֘�*�^�` 쏸F*� ���]Z��/�'��Z�D�?�.�y(	=�����C���B�Ep�9�R;�/TZ�L��ZwJ���hfR@!�M�T��((�1�RjN��F��o��Ue{��.X��#4l�5�ܵ�"�i��������ްY!CF?
�o�@�d?�04�Y~!nШ��~�R�M��6	����j��]r`C8���7qӸ�M��_��~�2��D��h��C��5�ΘZ�k�yj4��u��͖�:/��,�eȁ��,C)�aY�)���"Z�uL�{�=*@���x��3'���❨��#�7�l����ޱ?�ې8�xV)~;���uNE)i����_�V�ke��ML�U����>V�8���J�1�&�W,�S[�0P+���v�LE����n��X�H�s��0�ߏ~/4�ĕ�|)�H�T���i^��$0�c�(�W����͌M���J:�DI	��D��SR��5P2���q�qs${���dR�).ٓ���B�La+7�D��w=�ހ@,JGuj��#��bS�7�5x"��L��H��ϒp���I�[�)��N���8K�F����Zj�`�)ڷ�) b��9�hqI2Ь>pw�W�^'$`ؚ�1q�>�i0^<�.1��B���[� $��}}a�����m��+�����m��P�23
��C�����g��^�O��+��/LI�k�7���s�v�U�:�A�y�p+�w�/�ٱ���#�s�i�tG�G2����n�_�B>׆4a�w�^���c\޵�~�g���F�pZu�t�A�?�_ ��p�/˨8�1���W���y�ZR��c�D���jJ�5����>R9���?�*����V1��@엧�I䯦wp���n�r}����˂����P7���ã����4e_�f�-l)Ԕ%`ϟt';{&ߛ;����^zl��N��4[f���*g�U'�%D+V�
�%���I���$��ۗH�BG�lv�C����r���L�=u,��ՊQ3Dr�#K^�
��Y��L-���{6��,+9��������U8���.l�@��ǢP��<J+W8��ej��_&!?�5�E���5��ę���4x���
U2W�w�R�9[*�u����@C��.�4|PEفp��Z���ɓ�n@��LÈ�r�c���{s�+EN�k3�ؕ#J	�Kp`ZIS�H:���u���&�d�e�wrPR�s�w5
S�O��	kUE�o|,�-��;�!��&��f�܄=Zh"�%�7�F2�S;�p��+n��B��⿻�Ӆ��7-3�/u�����
�c+�m�&�������f�5'�l d-�H��w#�xZ��1��uP*:��T؞T:���XT䩉���]�if����K�<~��"�k�Ș��#	�C+��C}4Iv�S��*�?r�Na��O��O�0��!l��2��-��z�hJ����o��rZ��cA�.��\�_�u�r�*�|���ʚ�oz�=����������w!.o
���oCO�R`+���:���Iz�����qF�P ���� �t0�g��jꌷ�+�a���ac�[�8z*cNR����U=}PF� ��Y�3�Ϧ�L���b-%����v�w'�E�E	��d"��i(p��)�|�]���&&cE��m I[���ug��ƟS�|� wم[吙/e`�Ύ9&W����m@"[`���(}~�駐�!�v��	��ʩ6ٰ0���r�
�h�+�3�����R8�f�!�͟X�Z�vd\e$�8����'��`Э���d��!�����b����3�㶩�:�Q�j9#?��
�$���fN,��5��,)�Rc`�C�s�>V�P$S@R��a�v� �p�	s�,۪�3�Gwm�qg�Zy������j!Z��C�������Q%�a��"�a��.7�Sӱ��F���B�%�5#�IgU��]�^+�-��t,:TZ�p�=���~����4����A��^[�R���5�J/�F���-10�O�&)7�A�$�r�暾�k�]���^�@u@����.?�� �;� @��wM�S�Vr��K�
��X�M=��cC�^�؜.D�s����_tQW�1���J_Ͼ�n���!}�6Ҷ��[�/{3������)߉�J��3��Σ?=����7<41�A��u+��eH����ʋɑB{�j�SJ��{`��iQ�<%f�њ��4���V��Y��vr;�!�4�����ۏ���vQz;�ҽ�Ck��7�
��,�[�C�k�Q$��Ä�ߛb���x�g_k��DB��R{X�Z������K�w!�G�^���Q%����#��-NIʅzB�.m��5��ྺ3<�R�!P,��9t�'�W�U�"XH�b@�-ޜv���b��xuФiMI���Y�����CDg����#R��G�D�F�`@�8������_lXT���Y��Q�%)����q�,�$lye���ߕ�f��S=}Yy����l�4
��!�|Y��*�s�%NBq.o��t-�Mw�
7�Od�J/��C7�_�m��z��ۿv&p��bBz���sq(|37��/R�x�u���@�x��&B׺L�8yQR,��\ݡ ��Ǽ��=7�@�P�^U�7`�kG��+Ak�� g��v��W�����F���"x/��Q�=4��1m$����'$t��[�x�Rn��;�g��b�E���B&��E��A���[�N��P�\�}��Q�������jO���ԙX��rT����(4�Ƴ��
���2� ͦ���7͞+����L���`�qmE�j��u�l�5`s����/R��Xۭto�H�nD�f�������_oe���	�pn���#׎��<����ON�u>�����
pmƷ��K.hRd9��g�C.=�8��k�J3d=>D'�	J���+��Gu�p��&�p��m�����a���:�d����H?����c�̧ƈ=�=F	�"eR����U���&۞�B@�ba#΃ؠ}5�M�dg��O4f��"?"Evx��Ld��Ֆ֋>g�t���1��|8�;��﷋����Ӡ|�&��(=6��x$}�����?ǋ�[���|_ta��j��D��j�B�+�}�I��-+�#Β�&y�̷�^��<(��!P�RC`�Dnc��z*�X<C<E����6iƚc_��ˣ��j��Ͻm�����Vʳ��j�1?H���k�O��]������R�85V0�cI����f���D@�����'��YR�w�9Q���I�(8�j��"�F�9A���g�?5��Eeb��3G_@��������;�Wh����~��Z<GV��ZMgE�Ú�S��Y['[��}ǘ�=�d��T��LYn���u�Q��?��y�_�X��f�e���
(g黟�Zhm*5���M�.B�ݩd �R��`���Q~Α���=v�_b�Dd9B�I��#��O+�2��*��Y0��h5�sw��jp`�5��V�X���c��2�5[�Gi��R���)03�, �~"��T���ոÓ% zJ�r������~��%�)������8x�����YX�9�7�끨���W��������m_\M�>HrH��q�\�̞)�%>k� ,��B�t;��Y7�r2�.�>CGIkp�<�0̀�-���P�1	��D�KU��Q)l� gd�I�Rs�g����9u�������i�
�-ڗ-��8�~	�"Q@���M���z".���_Fx��w�K�,�䏝�PG���k��6[էZIlA'񯴦��7F��~?4� ��{�Pwwv7��݉&G�B��ՙ�f`�t�3ID6�~�<���Uz�8=/_�ܩf)_��t4��/flʩ�*U���BKJ�H����C��A��ֱXݤVd�9י�7}q���Ze�gsAY�f{2(ם^��?�;3M�X�Dy���Ԍ��j�����cg�:ho;{�#�&a��2�ʼ�!JO��F��W���l<�~'��2R(�s�F��h��Cb�5)a(r��jn@�������ʈ2����Y�| Lrp����A������~�:�=Y�{�����{�����
�8�Б�J�6��9�sA��4<|�)�6�C0�mܶEDF^"��'�oW�5-<;uܣ�6N:`k1�j�Ou��NB*���ܑ,V(����f���8����I�H�Ա��/�"<|�������7�O�%�I�}� M���I�JEܼ�ۧ}b��E����!��h�≓=��Z�CW��~�2��(u��y��<Vcz�ӂo�9)'�u���N��4<WS���v���J��e�K�_
�dci
�<��6�EZ1��3͘� �1��� ���۴�sȉ��sr��|Yt�Y8
9�F��^�o�^I�x�K�!�����N��bGd��U��؅�IM�ۃ��鼁F��}W����1 ��W�c[�Y��ό~Օ�5yER���ܼu�e����+w=���2w�UN�p�`r#1��C�u�3)�X<D��+��1��d,"U��<'Ys.CR)-�T�,2���hi�_�����a�;��fP�
9���~|\#��b(��
�����S��G��*���j"����?S58m�W��m�{]��!<G-u��fy�g�`D�^e�0�Y@��͔y
,�t
$�=�Їj2!*R��&���N#����QnF5���_�T��������g���c�=��lw#���X�I��P�v��ǜTh{1����]���X�R<�$}R@���?��=���&�8u�� �l[�TjY����t���/�AbFZC�Y��j�7�%\2�yâ��t�;� [�p �� =�8�8��hF�Z�Z�{� Im�"�/��+�UQ�	���<��C���O9#㯷�1��}� �$R�U�{
֠�:\��{�"�lx�5-m��B� Z"��K/	���:}����c�K���C��-a�T�_���^���S��џ�.^�|ٖO6q��RK�	Nt��h���ɄL��aLu� ���C�Q��s���=8}��u�)G����ɅǛ�py�[ W�p��>H�$'��n��pnѨk�mZN�� �Gµa<�T	����?O���K3jU�w�~	�j�~�C���O9U牟�r
�{U�s.GQx�ǯ�/0('��|\X��2�����U�Țb�a	���h;�`>ZV����M��5�z^��U�h���1���j��� I~�󉞗�/�_�LWCkSN�����`!���cI�L{P�r;$ti�׃�-�>�3h���N0�kUv?�8/B�f��/�Ƥ>W�C�,��1�P�ӌ>$��`�$��v%a�#�ŗ0�6I�D�'�je;�n�y��f���*|�;*}�L@�UY"#��(�cZ}�7�N5}kz��۱���R"�����ӫ۪Ex�e��7�r�Yē���������i�	�A��ʥ��VS/�-WX��k�/����e3#��)ԁ5ì3	�Q�nE����|XB�`����> B��d8��K�ܰ�/���Nx�����،�5�w�̵����+6�ɖ�����M�3���!��q��e����q�qtI��/���Pm��� ���#��b;F[�A�BP��>s��n�Ua�kk;Sn�?�ݻ�;�6��/������:Eyb;���u|����,�������̤��BU� x���-W��`x˘�
擃���R�f�k�W<�E_:E�gAX�-yx�S�[4��v����]tm�&����Q7U�Gu�Q3-=���3������m���U󦜙$���C^"�ws�?�L��F��b�O�Le���C<��.M�ܳ�"KК�"j� ��aJv����m�ɧ]��2�c�V�=u�7�&<@�e!�g�Wz�f�P�^@j�S}�P����B?b,�cy����2�[��j��i����:}>� ��u��$M��;��tYd;� z�����$�K�i�6}@}������~V��[ ��F@��w�}t{3���mao"^�*��/��RӀ��4s<��_�;P��?�VΞ�D��w���J$�Cg����������L��R�-�#��>���arx·EwkMo�U˾���>�g��I7�:�¿L��ݤ������FEz���R�ʱo�	_A�0.�h�G\=Ӡv9ˤ�����&V�*o(aT \�*��Kź�� I��^�p�.���ԦY���,	�� �:MK�3��*m��U�%��]y����i������3ҤU�g>p��B�פ�#�(�g ���yOHLE��!{���#h��~)EG3�@�M�u�ލ�3�n���Q�%L�i�Jw�r�/�t~�E����r��G�Q���IҪ[4E��T.�������E7�=�݅{��u�_u%
;�5�H	j���L�eó@)�ٹ����nWC��O1p�O�1<��'48=A+�00�� 3����-!"Cw�]��FR$	|H����m%�4�$�"�*N���h�-����W=�n��)���C��t6��'�.\jjg���(�\ey�Sr壦�ی��DDqd��6x�m�8�2�2K�Y җ�t�s�@�Ա��L�gM�b����I���i�J��`N�~�jM�@�Z�E�M���ʮ`��f��'����q�	���?�=��a�$���o<����Zn}F�_�>Kq3�բXm�w��я�E3���К��dg�~���;��0�6c�r���EC����_l��̖J��盀1�Dʸ���ݪ�G��qc�յ�\;���Fh��E��:��񔨁��G6;A����@���g���灋��u�%�vD¤�,鏦T����f�N�M���m%(���ٿ��Q�nG�!2��y:�z��A���7ؒ�K���^�j�P�sm%u4�� C��*��ɓ}�����ANNN�ϼ����7�T�u�ur�Z�2�ѡKb@:ԝ7��u �Ԉ_A�W����-8��`P��ʫ���0}�=���A�w��Lw�:y�����P4�ht5�u�W.��c�՞�A��]�-����|���`.IΛ@j��'�UV�-��"����d0;��\|bܲ>�7��+"?��ƍ�n�{�W�H��Wr��e��!ȹ����m#�]�V����� ߸.-ğXӃ8�<�7�@!2Vs�˥�V�OE��M:����狂��.��<������$Zw��QH1ʇ {Pz]u[^^8�}��b6�pG��P��d�d�
�������Ƴ��c�����8m�����$�k�@٣�}�r��w�d Ar��7�Bqx<ת�(��X�Dc�!���?��0c|:/�Jk��	r�����]Wc�gJd�L_D4g��F�2q���8c�E��ڹ[�Gu���!�Y�P�l�S�p��1�'�Ls�=�F��_o0�K��TC.n�W�ԀT��WEQ�aV��R�K8ů�?��t�SW�v�p%��@=6T	�&�!��5'��N�n�&B�g si���b��ft��.|w΃Z\	���Un��Z�G����&}¿_�r�,�8|�3�"��)����Q�]ݭ�OG��B�=�V���!�t��0 ɱ��ή��W�~���D��r�b^�����|ϡ�
�8��p8zDM@��>���if�b�i�Ј�
�����oO�%�v�$��AI[X�X��xNjh}��<���մ?|���g�l����LN?��Rv";�b��Ҹf�]���M�>e�x�Sj��`ORÞٻ���<���N���H�X@�1��>O�E�PDU���?y��'����*躍hiB{܅��$���)��܂?RN=T��p�3�@��q} +ݯO3�l�LcZ�C���C}s��G���|�ng!p���G�Am��~t�V��o 6n%�������6�j[3�$�ߠ�:fԻ�<�����z2V�A�Y���Ub�e*����\�2�q�n��*+	-�D$�a�]S��ъ����8�����'x�7�g �1R�]���֟w����T	4|�^���l�r ���.��<�;��u���Mx�Z�T��x�hճd��?|��.�).���q�I�u)�ƒ����I�xk�� �������h�%]-�����0�&����W	9,�������3�M���˚�JB�cB�n>���`�|��ο����K����8�]����r?���^)z���{���O�Ld/���������=:u�{VmRG�3I�e��ӿ鐅��҄�l#wf��<g���C�lÙ�m��hu�Ђ�G�_W�T^6L�[�yQ ��^+L�<l9Q r�%
<��.Rd{�Ç�g��.@'�Ȼ]0'�٢v����
֜0��YZ��f�}O��� ���N��Y��KL|7�J������~�16�k$2!�%~H|Z��x��_(�0-Z��mnz5�5z��M�H�FF�u%Pk�� �W���D�QGhH۫�~jFIG˦ Z��8v^�h�B���џ�f>k�N�oёVuU&{~=B��;(hyl�+]�h�&a[8h܎���S��7]��D�ȝ�!)b�iO��"H���b�a���k���̠���3@���G��%�dGB/E�	]�M?I���0y��ۀ}�gs�$�Uߙ�{>tQfE��3ke�R�d���!�f�iK|z9Z� [���1J�
z��Ӵ�l��wO(�yNg�ν�b����>�S��7X�����J�`��ƣCP���Rl*{����p�/2?Q�lT����XV���N��:o	�V�C����M���]<�"xl��!�z.���_�C�mlV/M�G{`���_���s�ԗbD�LU�� t�����H�:�#GU6�O>z��X���P��� ��\���w�}ݖA���#8�|�GI�,����N�ܹX���&� ڂ���Ѓ�=�Ĳ��IS��c��_ 2a
,j-��p+=o^�'L����'���&�/��Cx=����������u��e��� B�ܕ����}z��b��I�-��1�xSk6����;�x�rÀ0SV�4ni�=VN�^v��_��6��^֬�0er�QԐ3�1N"`o�33�C4�@`O�+$�7� �|tv:��Y�w[駁좱c�d>0<��eM��Ɵ٥?r?O Ya�� ����ƣ������Dg�+Y_���3e��?A�-Qa��BL6,�C&��TJ �	@Z�kywPs�5P� �����u�"䆹TP۰�m�=!��'KF�9 
�86����]ǉ�]�,���J��`�i�����/r����c�b"��8�Ļm�K���^g�R�"�ߙ�Y����yX`�^�@6b+���=�{��Q���%������p�ZdZS�K���3�e4Ѫٱ=/Y�S�C_ə<]#oA����	NQ�7D�)i�1��'�R)�R9�T�{��zyg���G�*tU�G�_�-�Xօ4�ְ�Pe�P�ѶNʄ���\�p�C��'ʺ�C.�`�� g�a�
��t��75�lk���B�}����6�|�s8����<���c�= �pҠ�l��"lr�9�*���N��!ɢ�s�N9܉5]��W�U{4�Bk�d��\?.�})�9LC��d�sU��p�M�,˒��h��]��4�pח�3����f��@�xR:��.=�p�3Չ�Q�&� �hŻ?���y��^@�H�Y��1y�8V�!,7�0���R�Wƛ���)���A3qB"$.uw���0�r]66�����`�1�r0�[e����(T+~|4ɥs����Y52��
���G���ݍYL���-FĢ���>#^�<�����}��1"h&��B��㻑;#��÷w�e܌�T^="g�`����T�`�2����s�sXt|��(b ��T!TX�wq��";�Ld""��+��1ڸS�0�����zd9 /�$��;��\���Y�/&���1O"����_�[X`v��q.7	*m�nfn�}:b�\�R�(��Dվ���c1}֙&o��eĨy)qӢ�A�h��v�rR0�5���q��h<[�\RW1f^�i����ՁQ��D��=��!s���8�,$�{���!�ˆ�I�f���(��"L%�	Ӟ�f�Y�� �����.�d�۩ڞVl^JG���G��3tE�v���c��M3-���х�Q[���>1��؋��|z����n�Uq�HZ�aĐ�rI~@�g둘�d鼩�}�3O�hq:� �������H���#��g|�����
�N�l�{=m���N�*,��h�v]��1u�۠����Q^96��FC�7��T+��+̽&��[�*�˓�m)\�����Gи�aX�J%c܎��������6��= TL�'dI��f�l�57-ڒ,�م���)������;!�YZ�]X�%M�mb��(ꜫȯ�,=�P�} �Sµ���l�"�����,~_�=�-D�/�������k�M���t��F�&z����1��`�ޤ�u��H�%���@fV)̢�T0lc	մ'P��="б�xO\Do�m�m��/j<��_ǂܵg���+�L�Qh˥�O����P�)ix�>h4z[7���^�ߪ�`���9D	�ْ�l�⡏�'}�h ���T��	R�jG �B��r�y���p����౬7���̣ ����/.������$�2 ub�,�&ə��7\���	J�����4v��eҲ=��x��#�yd��H�������#�tr;n�b�,��bdt��>�L	�������vh�������	8	�q0�2;/�J�"��姪iEB�v�Ѓ��*�-`�V6�K0�O�6�~��4����ry�9J���`s��06���C�&xI�=N"xsy������V��wZ{q��{�%��������q���i���m�Ja���ab�A�!B�	�$"�"�Q�4��6<oO-�G�
ŠzX�w ޓS�&����xmeC>��Lޣ�CR�v��lQ�h\����{!��<2����������`��@���a����VVS��x�|���Sy�Db��#�gb�<�{
@����.�IU�D���z��:6?hQv'�ԝ���g�K�v�ׄG��V˾E�-��U1n`ٿ����Bϔ-	
��LK���� ���H����Q$�Y�l�b����:�M�����_Hj���7�K���id��n��\��7��Ę�������D ��*r%�pF�	ֶ�c:I��OCa��iM|DP��x�Z#��YFxbH��U��o1�{�<җ/
��f���%�bo.�S�����&	���OXlk��˦��Ď�ӱ_�I8n R]'� ȿ�$Kf/v+��+���ĀZg�z��v������%7����_I��j�c-[����t�L�N1�ﵩ���τ������+p[�����73}����(P]T	�q�K�W|��MQ!].s㨻"w����Eb�7+���L
�7����הp��W|�-$�a��\:7��566�g>T�6[|/Ǉ��P��%Ca����1����
ŋ��>�,�� EH���9b��WgK������$|L���T�ۆw8���:�a�W(R�V 2��$0ʖF�a���L3G�N���D���@�2��ͱ�����y0\�L�v"�V?�oIBİ H�1Z�c��I~��ۘ�9Ww'��o���px���^0@�����&v�D=Ō(p�(��o@��d��hCK�2꙳H�4,ҕSE��k��JR�X)�)�����((�fg���c�ȓ�
��f)QX��AP#�:�(�GL\�e@:4k�t\�܀O>�ҥ�̡Ĳj�2<������8��)�����lK��W�&+�#��:z�Q)+X�H#�t�Q?A_�?�j��c�6��>�P�t8R�8���
�i�D�(��@��06�:
K�������3�	��J���N\�[��I0��Th�`O�}L��"�A��}4{M��&Q�+�x	�^��ν6"�Vs"��6#E�����먆o�=_d��2.�by�����p[E:S��[2��-��)�ljL�ؿ��
�
�$Ue�.��Z��\�Y`�,N����L��6�(�%Z�Y��0�f���,[�E�7���+�ăt��w��9�O$?�A�u��4���^@�t���M��@��[�@���2'�����ɋۮ��7q(�?@�������G�-�+��������<�3���䛇;�!PnO<� �!��Y�H��7�45�$<�?ĘFŦ�ek���]��Mb�u:�Y���Hs�>�Z��!�����g�x�_�	r��7A�~D�]*뚌st��Xg����*�4Q%Íˀ��RR��@J+|C#۵�h�<6�WP0�Z�LW���[0��:���H�ux�X��y��b���ڢE�I�i�� d��%JNb�J���Mi�=k$V�A7�>&!�H�"��A��� D�����$�"�0�y�w%Cr�C�K%��� �@�di���r�P��}R��Z��ck≣����%�ty%�:�b����z��������g�	;N/벁V��s ��l����I��a�JPDh 8U/��	�CW]�5�,�S*5
�J�Od�TGu��/h*v��p��ѯ��ސ�p�7Q�� X�@���Ġ摳M{��/�ew��PZj��-�F�p\i�0��\&S#GC�s��|0�QDn�XI��J5�2��J��ޔO ����w�lα�t��M+c��-zK�%�N�p@d��o��tD-�`ǎ3̂[��T��h�n� (���7z���.[���A�
���;��_���-��6!���<1����m~��ERYk|<�pT>�3�<J�aÄ!_��a�en>��˺4/�n_�
T�ꪬB,4m���ʮ/#����\n��o�TE)��ƛ*)`�a	�ybM�P� %��1�(Yf��=�������i�8�IZ�z_�xЏ��B����2މlT�m(��T��Nn��U�}�d�����2n��3�������J�:�;E-������x>�YO�V�9f����o߼�����9����QM�V�,Wf�����:WL��"���֐G�Q��E�� ��_�{��(���X��~)>_�}�.|�/�,o��	e������\C���u�ݰ&��xfeЬ�Y��ƴ
u��D�N��mW#	�\isHE��|�$�>����2���\�V%�ful�"�%i�]yRz�>NQ�Ң:��5ן��7�ke�m�}�'���Q.����k��
� ���GIƿXի�����w������_U]č��[�"n�#9�	g����	�����e�����C��U�)�INoN�i��=No"�܀*}�aC=�x��������4�P�)������V9���hdY�G��P�-�I J�qKֻ<A̓�z2�$��؏УZ!$A�B��T�ۡP+g���نA6�=��E�@|�R%����u�q*�No��a6�U��V����H��Q~�ؕ�z�y�E�N���2��oѭ,����1/NڙP�yU	؉c--�����/3���2#�?1 Tž�ǚ�9 v�Ҁ|���·k���|�פ)�2�%�l��6I�ϸ�����PK
s:�"�y!W`	u���_S��v�щ�BÌ�l̶Ӧ�4,%
'.����s��A�T����Q��7����-���Vm�\�����۔%㴌o�C�N���wF�`a�̻E��ٝ"6�I�n�.�k�뵙��oG�����}�P]�\�}�{	�S����ӣ�|�QW��r.P»?Q���RRB�?5\v,��L�s����p��_�",�������J3�|�96����G�\��X7L�J���G�����!u�j35����̚|)��|�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO���{����<��_��Q���U�f4��]`��m
���ܢ&.�c�ڔgH��j�G˂'�4��:u��[p�~�k�	-'�,*ҡ9���ӽN�y�GS&�G�u�l�"���j��;��j��r13��E�V	���¼�1�	�����Y��P���Di-�d�:A�C1��/Í�Ɍ6��%W�%r;֥�����j�:k.x�~�K�ˏ��G|/�M���)�8�9��ȸ�+�2���gW�� ����3}.�uI=��օ]1I[=�gL�<H�D^�����֍w��!4�I`���ȗ�ww��@p'@����Wg�`�0N���YG�B>�]`��cI�t�?fb�|�Us�.�ۚ�q̡Z�-x��x��=)�+�
b�88�����#J�y'�(�U��g��:���q�������a�	�s,�p�K�?w)��b�\�Ts�倇�[{=���ebU0`��%IJe>�����EΧ�9�^��}��)p�A�1��@�����D퇺���( ��N��t�;������K� }]�N^���)f����O�� ~GA�9�6�a�_1
���FFP(�)�Fq]��ژL��c��X��.P�0���d��F�A��ǅJ�����p��#6��Cӝf�(�g��'�``��w���e[�$8Hmg|��٭�T �}'>����:�co�~6�:�x�bP3��i*Xӵx���z�t��z�s}�L��{�z]X��I$`�Fۚ�q�l�nL��Y<��Q^�a�`V��[���o��WFV���@�\}ߏ_4JؙSn��zų� !|�g�V�~����+^��}q���bv~�Ğʯ��rTyY�F%V=?T�������; Q�@j:�{����R�P����{Gq�s7f��M�K�l$���|z�ϙG�J�:��{�����"_4�T<���*�Y֐��\I�|!bH�C؃g�!
�d�^�|�Ӏ�Gpb��N}��*��	���D�&@� 7�[}��6��{RG�-��ƿ����y���{����RR=��@I�;!p{Z��E�vPu���4�bUV�6�D+\��~p䐝t�m8��q����ߐi��NV��sW���g�t�(�C�1��ޘ�FF�{}-+
�ӒGG�(1�7�T���!��Я<ǺYj�X,��`]́d���ۻ�^�/�1��a�j���T�� F��X�%w���o�E�7���5�����xWH�+�I'ϒ�LJ�����b��S���E[Ҿ��)�����u����3�v������[�Qƺ�E�RM����j6�=fV��RP�>��I61��pc0�`Ԋ@���{����%zN!n-Byi)@?;��� Bq�K=avk���ن�E�
�+�S'4���¯;�d��`���D�~'�3��<#�ȿ*0]G�������L�g&S��q=9h�ɩ|�@d����>o "+Z�H�X!|&�����%�N�7��Z���p�#�O��H���|�v�pe#�(ge_��
ބ�V옃�|Ū�庴+(� K�B(f�a��N9����J['��c���ν9VK���%��Z�tW�̇�fǹ���m���i���j�H�}��¨���g��(�G|��iF�	� �0������F�3q�&Ql#��!��J��!é'�,�qRt=�]ЍGZ�+�c���@��G�b�aU/� �^p��Ԫ�Ū���(�x@=
�zj$�h?:�c���������Q��|q��t<T�;<�������l�zMF��'�f{!�(�?�
��p����.-u�j�q��R�E��|���V���<M�x*L��̨�4|M��;��~-��C�f]5�y���b��9~��c{N,G���LmCV!�OУ��ݷ�Y�b]����U������pU��&�:3ufR�Ʉd�x����-���R���\�q@sRS�{�?����ʡ�Z|�����|�M���:����OH�T*oQǿ����j�6n@�`#��S\]P�����A=�,��&8�t�*f� C�j-C��&,�-�ۀ�^�QgGP}l�~��ݔn}=i������Qs땏��,iS]�%��\�H�V��C�l�ܑ�P��q
5�w(��d���3
���<�*�@�)H?ʚ-T{׎8�Tf9��Z�)���\�� �iZ��o�M�c�$5&�����a	C�Y� ���d��W��20�ʝ=T����T<��
���$���X��21�h��W�%Z������l�c`�g˂�:�]�d��^�UQ�t�_{�Ő��&�	v]�7���cE"�&�%�O��gH���_Iʹ+��8�)�7_}�$�14A��Q���Yv�^�k��Q)������� \�I��*�WN<d��Jk`�7Z�IڿͱR���LZ���Y#yOET ��Gt7h�C2�?=A��;Y)����M9f��G��<��>+A�xc��L3'�I���!aV���^��
V�s�+�T��k1c�[�j#�a^/��e��Y��"�G5A��?�sٷ��H�9۰obP���u�����@�{���b'w���'�t���qV8��"�3�]����䴸^�t�g�@�����b���-�9B�C@�T���G�uuCE����G�	��}�9'w�#���pr��i=��J����/��s���;�����<?��5�k������TY�\��I������ ?-����޸ziG�H	G]�S֧�S��Q|v(�qei��rh����o�.�)��W�C^�U KKvx���+}`��s�C�������l	_�b��[�Wdb:���mTߨ�L)7��lL�=$Q�r��y/�`ꥭxc)�~"Vy�E|�4�)��8oyR���c��C޴(n�:,�=����;ɽ��͹7/|D���B�;&��@�1�u}���§l�0������}�,u&�{�[_����.l��!�x[�
�6�0gPA,I��kMv^�փ�7T�$:E��N���jm`	��ySkq[��5�nEp[��G�E��-vON���U��	�C��@�3@C�V���������gN].�m�0�-�E���,z�������:j��\�o��3b8ot�h�)��G��s4��`	o����S�[˩��>VS�R2 h�V�`�oSk4n�M'N�aP�W(�|יn�|�9����J��V���������Ed�:��tR�G(�ff���.��� ��,m��Ȧ����w�UmX�$s8�.�sr����3��+d3_��4�R�y�)��6�O�Rh`�[Q��ֽ��s�|'_HW�w~��|�O/*��#<E�[�pP[�	�����M�Œ,~-���k���䒧����/����*N���O�}rH�@,,��}�����_B,�6_��3-�p;Eח��%l�����Uل�^����W�! �Wr>�'/�:�0h��N}ڲ��T��*���X\x#���iC���V�{��^5�3<���l��7[�ճ��x���vOf�Ep�/����*���j�g{\���:�M��;�ŃZ�'���f}`�\P�9V�?ܴ��i����E�J�b �`fwĺ+,l]�7E*����O:�u�a�ߴ�~d���9p:�Jh]�E,ut<K�@���Sy�F�j!�=e���9��IE;\,�jnf]
�<�#�_܊�B|������
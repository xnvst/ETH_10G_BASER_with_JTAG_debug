// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:33 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VYvnR3Fvmz4mNIURrNeBzvIsQRVehDRtJ+89KSEWDqHwion4B5ki0UFp55ffa3y/
TkOlGt7XXWeAlJojeVzDhG5XJrd21ek+FcCMcaGehK/rA2rWsYbSFBn9L+j17TWG
vlPtf3MbcA6DL4Jmg78KlYdkNUP8jMKcptnfSFSPsXY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7888)
/mFpIQnTDlP6NLSpzkrksuF58Mqw/Tty7kkC7dS+e9VfI/PDT2Crcjx+u+T4osyD
uv+xBIhwsZ3PsHVJsaOZtnVWnHk3cwVP7XfB+KpPpO8uQP+Dx1fCTBhu44Y8Vt5z
RN1Jbko4xBqGOIq6Kb1hP9AL8uOF5uXnkMgOcOwAj58LVyapmTT6VU61Nao3Q8s2
rVFoV+qJz4VvhIRuw+0Gswld8UyguwVhDAMpWngHUTZDg9rAZLB/p2bto8HVAm8t
HZ8V7j5c6wrlcE/F1bslZtrPSDkznrVRoos5VWDffTyBNiELr8/r4VavUcB4yDDQ
2Cqqtvp5fSLsA6inEEkyFLvT9m8ihVLY1g/k6i6pQZDPGf8iJD4KQeUD/wUQ/sCc
zuLLN6ddTZSrl3aA7ZT1QJAtt6u1qykFASx+ylwi98m1p1UB0Ms3o8boUG+wzhwe
0pFGVoRQjxu2b1NkPCpodSCn/KsQWZBmpuiYFto5ro87PZUFyuBG5xaBF0tbARo1
UpcUyjEpEIEuY4/otc3D3teXO8OvcS9nzMnMCdcZHuUDzdJ6t/T1etAqVW8FfWfG
oKeVktdCRYr4hGRyjUoAT/HdBJ0SMupGLJu2VSoPMRW9PFuOlEyIWpNCIVyywRJT
fXg2em3cCywJzNvmtR5tWp4Ue2LBSi+VjxVjKSWHTshFm9GViQxLIAylsb3kPqlK
uxuhlof9i6yB6KvGkwWor9u4PMrfA2YiNIykrJBTw04FHBhVwUEVsyp0c0VIdP3u
czReJsWVP/D95EuLmcNld4LNV2VrhzmZrFFeYO4Wq8IC3147I5u/Gh81gGTyK2Xp
Wp/1pUbHRfBhrWUuOXFw26pgc0LD3AilnfIyYUATlkKkLOMtPIOq8Oc+dHnDJFD/
vzFbrjTlmK0nurJ1IYwVmOMmheuXxe07CrH7uZhRa8tVYTGWQD2j28mNMdWqW1zr
i2QVc8gRwMPiMVKsDtlpnsglAiymVQT5VGzBrvhmyQ+Bsa8ZxJbVnkBeQIT8K763
//iboEatW7oCJutpRKuij3smu8ynpt34MRamPcls4LCHWmDwjHWkfpzLH2ypNJYl
nn40ksFObVtLI6UkNM4Y6NZyhJVIZcLswcXdMhxcmHNUv78gVS6+9ot1EI/gnxJH
j1oW0K4HPA26xX9jMFHeT5Us+hrUMc8FOdp7KPacD4PemGMn39f2mYNZsiO3VmkA
E1aS5Dogiwj0a20STTmSzwkN6YpmulMKVcVLQN7oo18/DK4d96E1f2vajdM2Th5m
SelMT1Af7g9eJ6IAXW+7ntKWzy871eVEG5lz8Ys86OVfHMH7RU5v0qopfpY6kHxJ
BQrl4CPsDwCvfB6YupBEVMCnFgap3raslQ0Tx7SjUE8ofBk36p295Kl6Xp2r7bdz
z+5WQGVZiDwdt9P03LwkkE+VK655VHKIDrywhMAKKV70fZOXgg2vRM9VItOqBIsF
+/k6PP4xwJHkO0RXwVnR++ajpO5FboudEIy7ZdT/pTtsFQG0hSmAA+SAF/k01vxO
tf4w3OmWlZU24euVnwNl2Tq1QX4X5Khj2K2SMrf8bZi3GBlnl3dbfIaabDvFo77W
VUx4fnFaKiX1RJi6c9L+obmsshgw43cJs4SGzka8jETZXRuFi83roKgya+CvBq8z
mKyc5li2ZuddeXNdXktLAUCN8I3r5I2DYiFR2EKPyK4c9Rb2R03iUDTxn957Dzpe
ftfEHwkFL09ss3xEOaTK9SZlRhsCxvEmzsyShEA9QKbQf32paR52Mj3PiQNQz+eq
gFv/wJzieQEBBFw526VG1YgFogsNbOIt5c3tTSZJumzvaqaZE6mkGLVkNWvArhNu
bWpL8ewIBP7mxiNr70OCuJ7kIkZcummDNLyXeSibwibOQkYvtA5LYT7FYz80ytgi
bjque2/VaGdBSj/+wdcMyf8H2uQk4nNyggSJJvYA/vwnb5OMyIalNewq09bndua5
pYkrTgXthD8taM635ISAnghkCOn7qC3k8ChhfpFKyLOg/ib0tO6Pf90OQP0cg8cy
d1ML2jmDKi6xtBSF8gNxbYuMT37aR2JJAVWO+0/qibvbPzqOSwCzN+Axp7n81LtS
ptadRW9GBcjy7BbteynIeLRQnCKpGE0q/PMdId9m3yHufJhHYOMOgwDBACdkOMnU
9M6m3tVtGt1b1y8oBLzezSQ6o5TZ2tSqurAmM097x88RniS89pgkvJpV8QuC4iYY
BsxCJ115fNMgwFrBGwfJ68xul6LhAFQzwjF/ghc9NGIxkSBh0hWvqm76sbsLalzT
jHI2f4jeuFD7NcSTII+U5C1B5VWcJRGTYYXZfm1vGy4u4IiLIIIo0DG+o41f0kNQ
Zu+clE+O6Wx/2uDpFFuIoBRxy2xDI2Z79MU08yY1htxwdxEGPQFDbFKrIfs9/AnL
m8aQ73Qu4HeAqzKgG6c9wY2h4L6oE6rlkloRdelVlqFxqn+zMG/Ee7npoKgnzQQI
PyP5Iz7HuaEQMfgeZPJTUNE93UmeiGe0lmiiyuiEFOZ58+PZhGE0ZGZNEPlYc83m
HJr1vaFItCA7YVYaMJhB7IZbh/ztWgWb2SyggxepJlsVF60d63+Oq82sLEg+rzRW
oLA/yBMC3g7c/WQqw5/tVV46hewiZZ0AkFNXw0QYYmF/r8H0KkWdBL2+4qlqE+bn
bN4JFPMF/fT3pl7MCv5vdsuE7pNPCHBa/FwqyP8L5ktmV/X9pTaDemzNN3Zy+pdK
xC+5MQPnyi2c0rvROx9/6WUTs/pSQM3hEhBGids5iH42sjMLCOaW7l7YC50YTy5f
4NoDQpmyyD4XghOae/5k7CZrDtEg6nW6EkpcmaaUamb1ugVPOB7ZW+ycJqrBwpxL
IOvpdRktzAchGBi3XqwogEXnEEmNk6kIUn80mwZ00Ccnto8ouXEGWb5aCYuaKx5g
Z/t4id2sFWorzinBF2bbUxk1bQ3XU0IhcU1nYM0P3yd/7v3rtWgdphPugRoIxDRf
bIUL4I+FAIWkWk6i3JmEJSLJ7KU3kmbMFPgCSOZm57uxl88R9JxAzegYUJtW4Qan
36PnXjtwO3SqtTSl+GZ/bmpAeh22lbQOuTJIAXCTa277+sHh/Ipct5OE9rpkf66b
MWfBa8yd91+bvDuiWCp63a2jj+URsAdpaX6WxEimWXlRX4ku2X3SANvLbH86ROBs
E/2y06kY3sDR7b5vq9lGw2qlX4i5sm172iR/Wp6csrOJysl8CDg8S0lC564wQ7NW
mHxbdhv0vsG0DAeJnBH/6gaiPWihZNqWcGtpWR7Yd5GoTSTATrg41u+XzPJ0ZPQo
ZujImOK06fJlSGQ/RemmI5BzUd6iPp48l7oBDl5prI7+e1jNg5qwOiJacVW/6XLV
usmLEAlkZtOwjQmqntC/VoeJi+lr5NqMMYPTWdsUs3hrqXh+ysX3arpW9XD2/nvt
B41wZsqCJCKVzJdQIazd4MvFXb5jlklQiTLToPSxwdQT7i30P+18WSuXTiw1wmE9
kPhlbkBe4ONOQ0HnMNtDAZgKGUTEawQpDlHLXVMNjdDRQFqYHPZvokHTcW4VbG+l
Po9MuFBiMzoKy28kia8K6MemT/lEqCKMm0HZO8jHxz3RjrtCL530BZlyr/57WtH+
XeqkKT5dugn75/RWyCu8ggjCAcF/ss8gggTrweqRhC2Eh+GM1Rl/tpqPkZopf7vG
cW1P3GAzy1pAH3dx2n8zMpyUjE4FA1dWeFvEXrSwUuuWeOlGNC2bWunpdMZWvWw2
qWDguG40qPYAB93I9wFVtAv0fUDx9bqc7ZXLbfTONnSUAvBu3Pyu1kIrmB7JunKq
BYlwX1oK+7L2cJB8xtuJ9KBiL8kPDGEiyymPlwDVhDd32C7sNHpwFdKKdL8XY3KZ
eIc9cwdWjbtihx0HQBgV4YKbVERRQQJ/iOBAOafe0iDvOxLxLp6f9mWyb9I0rIVL
wD7+3vhYJnyZak2qOpJZmdrvQzDdyi1c9PFXnesCTr8jZWHQ9i1SV9jokh16n5v7
mQKyFiWfLTL5kbkJYzru3nYJ7xyQdobbGX0ixemJZ8CuWJOQbL79u6rS7ofqmXVE
+jl9W4THg9eOagCV9rugwML16MR21WBLSKg1n8bccVPermStt0ERQmCmty4WkmLH
/JsK6NKKZTuYbWQmIdvZVfPII5WJfO8s3qdaL9tSJr26UgvOUd2jYdMzg8SYhGvE
Wwzz4cBAor5PtCTZgXg7IB1AOmvyERgxSwsYNl+ICaHbNO+Q+1qmZfy0dDWMviPi
zT8SyqP0iWNtgKmVie0D+HZCxsxwe7Y0NBJZD+L2bBDbmlOPGbWbBchRXv8oa8hD
N4JHygouwRtYnUA1dPSgEW1AW9OWM1QR0JLUUlO/USbbDfhrdrdk2X3ycfGZlQOd
ExGrNcECG9bzZclK51VVNOTBPtvBIhRrhQctkGs6zYIxtXDq9LP/PafGTDtdgej0
24WGVwsEW/xKCA8xPlIP2jO/35TGlIF9uyymTLUWP8VE/N9SHSNdpVvvkZBjYQ9Q
9pxei7yN14iTjhk2Gd/G9UfNhhcUlpB8jTKGvftOAC52Rt5YOekvfl0D8kn9Gzn9
SAcDZ6fgQb4PNDyn3d1cbc4ZJI9VVRkIbfeCNKbKaTEkjmE5AwQ6euFsuGU0Tep3
TUeaTLN9WN9xiVQpxt9SjgxOE67hR9ui5hj4UGCRgT78derpouejjgNQxqEz9+GI
npEi/zYGaRC8572t0eZb+Sl484N9dEvtoHXP1oXXOBnMEdeC9aaL+YTMwwSFaqnj
fTsWJH2IkibIDXvmrtGyEAdNdRpPDd/teEg6oG4taX0XAXkH8V9ua6/wfVcBssVL
4SiLfOnpUV8Xwg2fiHBC73kmhHDVp4AT0sdsu+nZRpxAlU13FCE0/2p5GwI1GH4j
zO6oR6Gl7w0W7V5w2IVjuegNWeB9MoPevoPJDK7hJOHWG3Yw8Bpe5gOsVXjJRO2G
ATiooiisY90t9YOWpkNEFuMCQX7PbdgnEkID6fqe1ndv53P5XHQ7OVLWUZGrBpiO
TpIITyMdBMnoS9G7CHXNUQK55RaMhw3LdDmE2aGSRGbohg6JmvldsTBnaBkIaM9f
53JpsB6qRavoKf2Emv7IGVTPm9G6d+9TpEeS8K5l4BV5R9rk0xzpoIMP7a584u8m
WdP70+XA5FMm4kKrdOJSRJmyeU6ss/D2CVBuFYJ+cjRAz15lwWajsjaAAPcGETM0
9qBgkqQ4Tm/LL0DIRGmDhVTTb2eWtpHEgGVWI6rYvWbkRVVjW8uVcpUXUHt2Kfqm
Kwr+uSeYNVCQwo8Y9vcCJLNK/CH9Y8oIYv57jhrbOfGsD3RBn7Ebdv+L5xPq1yxD
uJsytgrfocpsqVlp9RbbG1L7jkKE0/LgI4y27urUQ2PQ+O56z92+eAdH+XECnF2D
FXZvlV8L6OCFKWe19yp18XzWZYOIEMMcTlPWqrlvvnTcj5pgwiXJJegZ4gIkGibJ
HjQ15ZnZ8AUt+e1kMGQva0SrSsdy2bgMm+O9lHHQvP/ZikYh4E38sug5gJa2tdq6
B9xP//0i81UzCbRKvJGDzDUwxrlmTPy8CgywG1elw6ce/x+vIz4GrAORw6Refx5w
GAQSPnqxQbWDhMgAVLscb8cnplD5rk/V53jOR74s4pfuMwLh4I/UxyjRp4riwaOT
JJXuj0my6DlSzdc38GZmVDoEMiF0WSE0Fffz9Zx8LTziF0ecW4Jj1e3K6c60rJrT
fAM/je2fJuyXatZ0qMkqn3ylaiApl5VujD4dZ8OeGEjnOpgf0C2k9NhudXkW9j1H
pUWadlczGCucGpKhICF78BH+H05oINvz7cyNIiSfBd+QQcHyCLYZ75oVweOPTcvF
4It/bnFxbTEnnVDJ/8FmKfMrDHexdlLO++yDwreAQgzTweC5R+kUVsn629tQvKlU
ufivb+am/YoijbyctJwgO6+lp9CWNflwIYTcP6zU5fEo2ta9SjI+vNRtVEhOCD+I
vfvC9oqeatV03VPuU9cgSM1VDBgyQHBkK6UP8GDcKhdHCs2QuDHL5YWpT1cygVm+
/xeED2QPucWsi05NkDEN8QYL5aEyHOUTaa6zicxlgTRGJAgdgzUPLY+/AVama2EM
OiRzg841UwSVp9Z6L8YUUd8dp0ztxM3oVvtRYz7YMRoWXsP703VDYn8stp5o66SY
3ggEiNcVlYCoYp17/wCma0GiKZ4EPtGXQWm7VHqKlNqiZqzALfToJ0eN+h7KOPkj
2dq6htweQG/yfUYxXnsNE8rN1hDEvhqsQN49iq6bYhblBi+vqtShd6WnhFtkh7un
7XnzmcOX3wftf8x7X95y2diCXxebpGLicVsG8rcLbVeYoPis0nUZsQQqX8FahI6N
M7UOS0UvZA1jcRlFefZueWHl1HQTbqYSOcot1WQ5+wjLgJdAsIcPmg/c/g5TuSvP
s7mI/zD73dTHC4SYj4uSJijswyq1nSa6RtTtQwY5AsEq7Y5u4DYHSKAKY5638Le0
PfH1SIeBcfS+qQCBW0YrTIw2s/pjObp2bA4M8wXVZiZvxXh4hk/+3Gz5Kdn0zMD2
2B9CYnmnqHjq1wwrepip0JlFkc2+bBjvRXpihXzqH3TWzFFErI4yjnxTDK3DnsbO
akq05R2QlrWw3sBwgO+Jyi4NI3O+zg/0ljcLxPzNFTM+p6urYKxg/RKT9hSKaeXH
qEZdAhHry58d/hteavgFBpe3mEEbWab4m/zLmSlZKyAOVbZhn7SBqUyN6jJ4au8Z
WO/I7xcKQrfkwRNZLUAkJzzfLvYDUtCM3B5d/tF6W9uIec95KrwMHEp7GyGnxCcq
SS2ru3LXBlbNsNGdfP3eq5sbeykJh1Lr55+P4NdOfYk6rkYD1Ix+6i9nciK3MtWF
LycG5MbutPgKt7vKp/t3+OHQlg5axSc9qzsmmvDF0WZsYAh45ror4YAczaei3hf8
Njx6Qh8/61KBVhuqE9qRC5sEt3qiCnl/qeaP/1wbq8wl0D/RTr6POHMITeeb+u/0
dKvnKXhD3mFi9xsxHTLkiLk7nxJMe+u4frDOZYXWqIV3Hn0Yy3tVI0j1/FdAK2aW
hgp7jyFPd9lgvVWccD4zcGUXsyj/d5wtVxXwgS43QGWjytc84EBUYg6XVhyULsVC
0AjXY8JzeYW5T0pG9hZ7wJ6vjYMsOR94qvdmN6DPUPf8DnNCaIZrHyNOdKUiDTjZ
N7zxdeSG9F/sD/WZX43IAXOLYsFXmjEfNmko/fmWZpUfPbLJ1C8kCnoXpm1xd8jR
E1XwlWdKHD4jt6hj92lTKAkIrFCQulw16Vq7a6M7l2cYO6aM89mESvA5ViLNhP/p
pYat8ZY6oqF3W59hYx+wEVOMA/1Xfp+lWA7vXwJOfcOWisUDjgAcE/6YOc35OC/g
/kCeiI5hiAy+LwNClFJXfMI8UHvTtkSTRa+f+Tihj/tahe6dqtANAMn+r8WDD80d
Lu0aBjpNd6xFBsyjiKPiPWbsxkrG2+yi1kTABamR8cjkqwPnkweUoEFjbDIVvsoY
r3ZZauKg3Veo5OGvizQtMDcuYRWYoW6M6ADekBOQGSDj7c8/0KbrlGebmFiNuM/A
jTIMsrtZw8hOSW/M56gze+q60jtO4aTLf+436LuBtJXb5forZyp4WcZORHT2K4HH
W0ZhJuHmcBaEsQKOwcoLv/uxbZAGVTLBGNeZPeHr6r7V3IE2H9G/gTiZpCrUeVQu
ODmVMh1NBAU5maL9pL82cSgb7OKyI1By1pHMxUMqDVaa8iwQ+32EUvHdzxlg22mq
6WgZmHd0JHhR07YyIC+NAgc2yU8tFBHT+yYfVMOrJ9jyqlfCeXACWzVphRGGpshp
bKF56L+INaygqGiNHuofTQgTGU+La9jRHZfNFCLjvosgidBKbCDAove81GLZVpYm
aF4oRJdhux5Y+s+5rWJcKvrk23mvrGH/lgMKjDBB+4Ht05IsOFad/2K88FZhJlI3
i6FDijWeecv0f5La1VxYPcQ/Z1Bl030kewlKvkYj9RZIKrgvpO64cQdjsKQAqjGU
VPZDSaT8EZN4h4XJYacaHMogn2VvZdIvwvgYnrroTAH0Du4IHm2r/SQYHOIUcx51
Ax89TUWYRg/DBNS1rkL94byhvc/IP345s1QcuzPBrhIXDuVnIJ/n0mTnNuCEEkLu
y073pr0I9iPoYD+hRF43StefbBqAewUJxYHFZMKIB3jaEfOA9OXdUSQYAxxB7pv6
7tlHzZx/IzX5tdWzVFbOLoTbQO3ICYxs3RyZfqlsmuXoVcxSl7bF3gDrQY9byDX1
d+mJrbiRXEUFYj+SyP53968IAqRdzaJYsbftyQUpGS8akZFKu06tTLkKYtz8uriV
6ZHQ19MXp2t2/smiOxxmPrJWeC7HquIHwFHHrVIWu+68lk1Dr5jrXsb3+IFudNV8
yaXQePBm6bBUr82tOBrfNeCMstFU2SVR5oLF9kqQZQMBb80fA58Q0bw0okj2R+t0
P3c0xIVFAZzaap2YVUHDBvigcZ/iCxLHgM8+9iFCTcou3XPwdoQsLf3BldPg16Ho
Q7rHvGpzC590Knd+qcBn9t5FDEDmuVUq0yiYDjc7p/3eVtTgvLtf7emQi4KQQQGn
Xa/G1c1FthjFs4OFHPYgvoS1glM2hskQWaCUJqw9czgYalUOVMfft6YvXWQ0bQnf
57TWuaNUmf8lcQUZVqizDry9d8JN7DKu6WtvYCBRQudf2rZpfcq/9dUaRTI4bMDO
vWhzTmcfSOqQK2pXr0IDCSEJGr0AkoyCrX5hqRcwOznGyvs+BWOZ3+d474bxHFR5
4y/hOalADuA//N++hUHz89KGtcgPUfjW0c/YOw55LuMl+0/vg56VgDtIk5TDUUDe
K1VKoYaRDMeVTWZ+enmwugodOkYFSZIHO1LAuZjdEcS4vM4wBHsCwS2vK0NvZrx2
j9EpRxWQZYamtnexGnZI5SrMLxmPDI9qpiG3POnyHCqRFV4uXfAUf7MtQUNugCcr
uWxoova3uPDwezSHAheFcFZ91N/X1A4hvnZcPU13JUN1QHtXeOvKhL2FBLJB42aY
zoKjaaUM/0D4wqsI/1oIZ61dd/aiXoF+7ttojrMc6b+4GSlzUFszggRHqiHWzBjM
ossgUxKf2uHqJbO9RvOTdMuVOLSPLY9tQ0XNhFvHFzaWLo2arfhW35m+jvIRGB6M
yulycmRVpiEgAblqB7qkfnKZ5PO5UoJ8hEJSlBhH6F8dr8ZT8BKXx3R8fUjgpXCE
Dt70mmc3OGQPbISvKCHsKApxiw0UdIrb8aL0pxaOVI+0m6tUJ8z9VH5Pp73a6fU+
u8bUb4y1akgEKkQLnnNjmmq12iYlFBOLYgTKTWNEK7wG5av4tj1tdYBMqqeEqxFg
I/drv6GtH8DKh+w3hcVZRL3EDeB7cB14f78e7WBODHv/le8mWj5Y2NTmZ1mnEIgh
0lokK6/D6C28f+DC+tMXgkr7jIVsSDyB5nQOwGVN5sKyClswPPZJXxjm1LFRAyB+
XrIFQRglebLi5bOTSbuUF8AC+bDKrumudi/i844Qb3piPEMmspHhv4gBnF1SXmW4
iGGNjbeZrEl5eZ57Z9ab4vAt5UnTdvm8iS6fJI8+4JPbl8Yy+dYL9wUjG0v8Gz9y
boxuPrfpcObyBfeb+tn1v5YQ1swYJovrX5E+BM/wX7PB4VNHcNvtHZ6qmAyXA9A7
EYUrKUxbloJM2STB5Pk1cU9FNZydxM6yotvNgn2EJHxFU2tg25FRF+uIdXOnJJXf
qcc5v08U7XIfDcfgbQqh4G8WZ+r9lBTska10xy8UXLLWvs30a2bCohkbadI24iL0
JXddQBr7JhBbq0BLYATodouvjaJVrNh0Fq3mhdp7u+eVuUz3l0bWZ5IN+28p4Gg5
Rjp/f6iDzEOxDzUg0vQDOWe0mfBMtpx2roxscaJ8mKbCl3QjxOEc3tnpVjeoVUJZ
KaaSrznxEGrwk7sgPoXQTRp4nCEoMnzS6+HQBTCy1kGmC3n3l3GLp4r7NtkH6fYA
L63hmnKLNFDomIv7YqZ9lXIDsTmHqtmjuH5spaydIfSk5iuo1mKgBNwhD5B4VDDv
aqWJyoOk+vNa+wpPlM/CXO3ldqNbdIUwAC8QTpDeyM9qOwm9DK5uiPvCpjOcSCjW
aF+LppcwC3yH/CQNMLR3Pebz1wIcl4KTjcMXjcxWz/1Qt2S1z0eok8dv0zhZvWJI
kc38ee/Zzhyw/aHad1UZktivvOy1vZcCez/Jx4rvUHGS6c+i3z6UpwzjOYj8Cp/J
YjjZkxhsIV7Z4XaHtDrTZPwPlavXol/FJNWrT6sCh6ioNZETLURL8zHS/lpAFjJx
tI1gkLKHQiT6XG2KYwEtCKSLAKH2TTzyKdBIMVC57DSeb14JiuFlbEgjr0I0TYsy
rxkgt2aM1gFFy43qB11sLQb6Us80sy8oZvAJuFim/UhdXMMSw+1FKlOPgh1lQ8N7
l0z4czfIq9PMpZx3/kDysA==
`pragma protect end_protected

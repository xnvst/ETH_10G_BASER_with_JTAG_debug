// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:33 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oWvug4W5+T79PslhMjrCaXNvFRJLcMo5Hy7vDqa3nYgM5wNEfqcKhpzQzGAZLplC
hqAKUjwsF5dLpukihYK4Xm1Og5BrQxDDg+vHj9fXfXOBGPnb/SBZjscIb147sPWY
kz2ZSuytlQDdOk/ymTHnq5ig1m4c1OrCgY5iNSHskCU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9968)
ffX07Abf07eReNJSh9j7dNb2Kpv8uWyhdoc7eIQO4c9f+RUq7f6slxQrRnhg1C55
UB6vlrTiJucfARinVeAM3pZnzR4DXGLN4j48XAwb62RLt3JJvOWszA44/F2vYRfs
LopXgWM1RRaFSedKJLC9WM3fXP5VTYKo8gWaNIHGn6LbCjOhq8LWrBzOryXhrLzA
D1Ni2mJS84CcnLdggcptXiCwlDvnYa9etPv6D/Rc+ig8T+dY7tGGpXaCyIVaYzIv
9Bnx7B0+4PaVJ7N7AZsJONPBa0o5EZ/EtOwInp9zn/O5xseLLDToQ97qPZpPVtBt
0rwNLSwzIpnD/Vvwxm7ta3evrGehCObMziWbNAOyE50j3T87pKkVdNY50XSzVY/L
/aiGtmjoVR6BkLcvLInNJ40ZOtYBlyp5SQFlvQ8cSJ5TT3/sWWOgE4ZCRbrMsss0
Y7ir+lv8sA18uTmT1npW/K/SehvGDQ48KoMsHILZmuH/1m6hp8RWtW1ld9/TqUNC
gNNFGupnKztKtfDdwplC7ccDMG1P6j6uOvVKYOMmKuf1vHFZ5wSl0D6GrueenBUR
BvvftsVzgBJ8hE+ChquuhHArHYYXkZtrjW1Utjw+74OBGFuVoO2wFL4Flja1s0yj
cuiAR2p67F1Xhf/qP48Y50OelOvs8W1CIW+eVwi/+R0f28BMbKyK4qbStNprVGyq
ExBskDYXPMuyX6JAve921m6Rtz73e7lReZiK2tmQpVfOcpN53eNbPJXwu+2IbNfc
447fMsMyowZSEZcYSB6a3068/l9qgD4WbaLqhRKdRiejz9bRXfiqIGuWry40NgoB
+Gl0RF/yvs8llGc1qIc5fJhV7UPXcT6fq543SqH7g01vMcJYoKXwQuLJ7GXCXT1H
B2DAE1QUJWd+1ntliHXpZumG2CUrgzF8iU/dET0cDygGoTrT8ZCOob29BkZGVNpk
imx/i/p+JjVxWSgqYMs67+pnN1yCmTEKzyZKYgx/DBM5/RoH6ze8fCVY2difW9IZ
CfdiNS2CLg4cNY0NgC+tdOPYlao4QpYtIaqCjqrecWOmpDAZ7SE7E06IRsRidAgE
9c8CL8SSiXlrUKeaDk+Pv9LeIOSQlqaqImaOQO/DIK+QabISMMlFQ6N8/5PxyQbY
M8rXXgE0GZgX3fvYdA93z88yj6eR7dN7UT33fgULNwHp4NaWZBLAUHQ1dwPu0jst
UvbtKbpOz0GoTuy23VrsnHVOE95zm9V2qdMxpix3haiZ8AgUl34V/KhLRtQVjpPU
5NKoztne+FFgmIsKVm7vXLQKc3SHB1yCg5geaLfsIBUVDeQiaL0lVdso7KDRQ5kf
cNJYhev2AVlg6qawxMPu7mq94OQWFAUNGb48xJ00pZ4U5Zbhsp7LRgcZODimVtt0
YJLU/5EPUtWorgbV9ypmmAHGhibcxCzy1OXFSm2PvpRNpBihAk3qSe/QVVIfcjDC
chLPXDsOla33Zft/ROIwn0GJx35aDomKuH3c5RZPx1ZcBF10VySRIqsGfPRZdqKB
35IXCTMeWQ1kp6sJE6qv6GEjcPPqpUJ6yXjB/zOtgFwMvjUjk7xxBVQ7oiLb4rGO
614SawZdSmQ8HDOjPCeDDOzUH3DQ0FBu46LvqJL9RF3hv1lFHgtuDd0PmukkOpa5
6c6XxQpd5RVmH/VTSG0/46nWJQY+OAzkm00hgTfLzcW49Xods0z7iydDX2WT31t5
W3LyrdAY2H0dIHIKjkqa3VZTbvSswaAgpxsz9vcbE8DgPVoZbwEmofjd4Ra5ilFK
x+Cu3zquBVa+L5JQVAC10jHcbaho4n1b54WDde/3ut/nU7liounG9paUO5yL2oVw
FiJ7T3EPVtWd/Zi36REbZOSL3rOlEd4fnGoMYZUlKUQjNGbEkbzOUR0PQmInBpzJ
l4gYPdzs7SPhIGNxPQoAUzZ7qoFj+tHyj7S+rjIBdptudjFB/sKX4HQUGAW4oadH
pKD+Zkd9kLq8kSii6cNqcxaiCFEdTvrNfDDNYC0zn4mPS8V6y1ODXa9PY/18uS0K
rnPTrs4FbdVlCFvGfMMtZE83xVthn839QIJez/bW8x30ym/UVdtTCdCYeNsPo3el
5/y5p4v0JeYqDzcqaJaVBgM4PFg7LnC+Ot24J9FxfJh4R9HxW/nNJAomX+UZqbDJ
PsD9cobNVwBpT9rbZJyam1p6C1SCv7G7xjmBklnEtzJGrwzYZJ2E9YI297TzKwm3
wn9HmpN8P+yXPMs8dhgvkUCLHOAsgF+gX79YFICYZCOiED1vCKqNnNGHvzgbYF80
34e2NHwf6TNx0HNU47de//VoEY108d1BcHY0+o3JYq/87OmgSbw1PFdI3YQU3gPf
7mwBHFuto7LkbXpJXGrlVveDxGH+vP8om8fscy6RaLXcKj7ml4jj/gA32UEbFTqt
ObFvcZ8muYFuC9mmlxdK9sKZOr3e+cEp5amGNbYgLh6odlzoNBIsZ1iwiy1nALN+
vqqcg3e9iJdVNa4dvdPf5LVgOv7fWcmAbmHOj4YLAIahJDKIV/wc+GCpUPXdGTjU
rzze4WHrN3YppfIipsyHXXrK1krcuVxXLHDscG3Uq1cUFMCM5pD8ziFE8AUDiIIj
x3ussvRs1CWamAamat852Mc7UcJU9NejNXZFNLsRh1lS5RbzQx+mf0o6wp7fjBC6
PqVQQSMGGuPNcIH/xSj08/ku6oFsTcOPBXkDTRBBoMNJRMA/HZW75hUBtrU8ra7M
nwf8T4tn+gacHzizHF3YWM9lnNjJncDzPpF9K+hpgwbUuFcsCF2E8uB1iIy67kkR
oy0w8LUscnGvHUW5l1jctf3aM1FpEGhMfFnWh0MpxAUTlYCdjKGlhEJYQHUboi7g
czCyEXUceQBHgY0UD8l0OhpmYLR2uHL9i/5n1iyaAJGgRJm8D94znjTRxoNbxd+G
fl+YF1FoMZe1uoXJJiiR8SeGLEUWKtlez2otQfXLnNyUkU/v5W5da3jwe4d5wZRQ
+SBbPYf14TaLXoMkWTc3z58eTFVd5DpK4nunnixx7j0XqOxlB7RbGlrGfz4S1LBF
3Zt/tyiOf0qhO9RrUK7pDy3nLF6m00aI6KgwuI1Dh2fieFrmORaQ5bAqcmdD4sTS
GtVdDNGYXrtXBCznYxooonNeyituJGAeBbiirnOYB8b76xN1pgYXYQVfBIAMCWE7
ykulUbuCioUKZt++zdWf/XVq5t0uLvQHeHGUufXO2hKJSEJJV5IpTimGCcAGkdCc
UbFCthwKsJsLDnXmBYFae3CvMPKiUojGAHijXavuulUiOi/6FnKIisPTDRr35sVL
aWHeWNBIWJueCgVFdMF4iTAPO9gINzOq1HvUlxi+W2qcEj2AechUDDU/WEmzAaxy
e9A+3jRz4t6NJoWw/9CqwlNH9hsNhL9yMgiyrmWnZtqJB3ogN363PUR4HhROdjKN
Zhb2Q/it8yRF3a3bGIoVk+ZjRj87uHaDSbGI1RDoFgCod8QPpt8kKTY0ooW8bm/i
86xCgr8aNszUPZGUDE/3WxHmZAgdTl0gWhvyAYIlid+m1j7nI+Jo10YRb9+oPPKZ
XpVBAFsC1eZF0+b5oFuohYJF6Enmaz/J/Im2uxcjGa4Eiy2cT62aISPxivhVbY/Q
37QbKUDv8kM9qSS+6LwVg2iaV2T3tFbpVoHpCsfHZZ7Yca1pG9N+SdYuewis93Tf
46NVLsVg79hpZHBEyJiwjxdcAARQOKgImdbaiL8NVNJGIpAsjn7GGG6aL5BK7UT+
HLFKGvfkvtajOjCST7ahZwXWpFOG+ERO36RgN+7BkNJYaVPkL5L13lnvFg8aoGIs
68YhAod3HJSi3j4qXJ5W+lMvnti5rYfnU+BF2CDIeJvY0zzJ8aSpV2F5wIey4uWW
BcCG3JEcSbxomy77X4ch1TuR5K9G7ozo2hHPxO6+1b44m3zSInIdyJn8rlJsxxuR
x3LMBJHGru/CwEslhKOqg71Pi8ErEVzG0/31vYswjZgFeVXDkAa9slEGSByR6D6L
NljacPkM1ZQxvEl1qbwp2h//oeo+8/VMQtK/tW9DgGooH/DTM/RElpDyXsrtWjBD
NnXRJrefRZQp8nFZs9gcPoBzkO/n/YaTutDDWb3lepf9qcdu/SmPcD10UyTwDjnU
48D/gEQ1z1gXRQqdCh6BUwPoOriIwkWt0MlesY7XcD8M7Tb4UGYJsZCjpEd/9dpQ
K0lM03SlS8DrKyJ1wC7pA1gAKxsedIUqiPw0ce8+ayLwiGfSxQmBTyTZac2OOXD4
6vdeG76wutXIym9TslYpmtMvvd9gzsU2ZwbxyhFaLua+bZLCu1afVwAhad2X0yEr
sud9mDNZ2iWpgdDhbAxrhtwd2FrUCt5kLEeb4FgEzQ6TXquGbzxuq3IONK2rnpJR
t27NEHoZc8D/gXIEZpnWiWaOhSWOOP5Vf6Jyq2mr1g28JmQp5xzYc+vw/VrW2KwZ
8ZQV2SqgEKqnfoFWTSGTDYd2CnDGkVygRke8r12Z69uDUQggocomw8wDjyPanJRn
ETibe6BN2HxHWJpG+WrDDKO1VC0Mh9gLVnOQkiYPmmJzwToAxqYe/SAnKAlDFI5s
8L4tkaIT0WK7m31QeZNNHHIOVdF6Wj9solqLTITrh+sw8qF2ogaKAyZMXZQO2zdA
XPWgcrtCOyWAmAL3qW5NSf2k0ExlbdNFyyecFJCcfLFGBzGzoqiL5fJI1i42qj19
hEAL22PfMakWFpTdqOeCqMgsqf0Y3iZmzdo7CajhTPpzfbDU3FfNWOqlJUO5z5uq
Kx5ZhHdVNUKKyPMaIFGrCx6KanzCh2IL+MyBq0wNlb/wiahQxvttxEkcQkEvOvnD
6BpMVnecAiLJNLCSTiy3mirj9M6Z4ixjhPBImUH0/vTgPi2SDo+ZrfdMif8YYaQP
c20HusNwnaYpY6C8P/RM/jeAtkdlCNyatW/uVJFbeLXLruy8B+F/KAxnmfAvnkCf
BxshCdolp44uzDYngDi2ysCJHg2NmxqdnlRKLEKkwUpoM0GRlZNe0VyAa1NansMT
lXjEbAIk8KN1H4P3CIQoPrr/4Gm11NdT4pTgxhWR1nPoVE8CJWKXT7kMfUskUPFd
I0oWQUw1ygCFlUWdtUrMKtfq5W53wtFiA3XELC+50US1V8Zg1TzFbXe6Ng0Cukul
wFGWZj94jCpGJFv+I2shJN+hC8VV+aE7bSl8TA7FOW/lfka8XpzeeLx+r6C6RjzD
6Os5rzJ1WWQDHq4Az9UuWkNKWKUAgidK8dfsQForEQ6d3w4d9pJNkbw1Lbgfr/+Z
My0bc7HFLD9Oh+mR3evGJG4JBMloNkFYA+a5O5nIW5lC/DAPxDWMcrRV1Li88CPu
/MAMVGzlB2iqNa0S/5RfRHrP/uCRWRwKYrBufEoMDTQ3hGP/JZuRQDUr3SkqyV7U
Flx/M8Wq/yzb1l+HFthOswW2FiIfUwckSDSbikZKATnZg9X3/Si+bXKOpF70Zw/H
qlzG4MTtvVyyRXvBka02oBzCwxeoBk3UJ4RmU39dhW7OgiDTxHhRReJKqs/V6ro4
DAGF+858wd3VAFpJ0f2SNDbsaQlHiKgXn6kqzUpf5wRK4+soEri0UPD//EW7skNP
fr2zgNjhjXD/wXURdlMCxQmu9GykxYx4cMEMtbNiCvp7pz8QXcKy2Y2sUBOB+r1Y
mTh80vG78riNYAKuQ4XXJRYc5yPJ2zuwYiXlm/3O4aVjEP3gCQgsrihp8a9TDspe
BrwepBqCLCybmAPVdBCM8gfZaqr/8sUxcuIBRWJP+hsCggwbslAyiDLJprg8I2Fe
fvD+0iYDSyhZukkx6ukWby003mztJ/y4l1cyc+TgERLqToyXxJtei0qH1T0mqP0P
GVKeL0pa9gH4vIkJ4gtaJXq/VEqA+DJ34eT42olF7tLA1pnGsGYdmc/QzpFYxAiw
F3EMfZ4DTmZUjZsahHWrHrW7IXuFfE01oOgpMyH8XrpiL+W1v7xvozXRdHutAGsX
ZOFzEPsOYaxkcaul5b7Vg5EoScXaTdzPdpPfQ2fJGac6Cc6PXC/5mYKtCw8D/6xW
ljguEGytO5DcJNHvCQMmblyQYeBu/6zhA8meswqPPd3GOfA2fb8ybWhPlAHNlzYY
cLxUtOGoQSU7D/5FECXME0nGqiAnpZA44fUkmIEu/peZnLCT6UC4s2DIDGtbqcQY
XjogGpONXf3gPghVVBhYS5h1WZ+hiUDupGbrmxmolE5gXMIshax9AophIH08r4qp
Of2oClAig+LvWpBsShQfediErmq6qKLF7fii1WyUai34DEeIDsoy63LaALCmYg85
s2KWEi7/IKc49PvUAW3XK5n1QXukCh+UhFV4UJpw7acIpesGaMH5uF3NvWENFcVz
f/4VE6hkj+el6TjYq3/DhsSI4GZWPzjpay5kHpDq0fIBYdKdmOcu+CXMc/h5OLjJ
b6kyJBZGUdIR1fgsTuDKRRl3xgkt1Tq1WZ/IybW7uPBenmo2juBQCj2SW7OBjFe8
TW/TcqUF4g8EoDXAJ4fJ298OaOQSV8TnLViv+69DLjVg/ERHJYj5PXSZpY80It0m
pumOdlXu64Fwm1CiyXt8OdyXBV7zkilnf7eqs2mR/JM9HPeRNNhtD2CXfiKD3wC9
2V489kH6bO1ztjNdwBKytfn2XDIqbPamVioBIVU+mK2QQKTnEb8UxJpdB1IB9zxg
vJl637wijNZx2Scqx8+UEqQJYBqNFuP47HTJPc+RfKsXDtTCpFuBsleykwzSIXDC
MYOJ/0anSSs9Ot12uyoyzefG3bBlHl1bfydbaPMicgMmxN+WqwJ5amFZRuZPUmGe
CN0KwRT5j75cA9x8s6fsxQAEfEg1F65D2lujzPn9aOwYPgDeRb0XDHvgut3pIAQZ
mkpA9SJ8XSerwWawSH4j3Y/nf43yi5cU2OdxopkPmucWYMjOofrfchg8vYgpPgSY
TeUkstF4FkKHQLI5CmZ21zKsTRqpx1rUB4cqjfa0iCghvOUwBLz8mqRe9qbXBHmh
JTiitNFbb/MNFa5ea0elQRxbqBscgnTEDC5ChsZz4CdjXxtWB8hV3wh5PsfdhJC5
0sEV0p6qAKw3yz1p+nXyqclb6r9+fLOUzuxOfBWDprtyJ47EEJRKC7VNtBIxkJaC
kP6qCbn8tRT5xcJFxQidCuKrhzEJI78vJ3k1oJ+7ZX2Jd7V/A/Yd78GQUv/GogVo
zXdFdmD8ucZfZeXDmgPRg1cw6H+P/XVJ5YOOQ/q8C99yJom8SjlsRUzP0WTZGxlY
H29rA520rCVbp2K+MXQxzUIut2hApMyNFQoJJ0RAwoutcbrYTF3C3qUK6/w9OAGF
UASC3UiTQCtXXWHglhF2YDOgMwVuFtSwdIPvHg+JVNi6NxEY+n6CBszsB6YtFq1p
IAzOvwI9H0Ex1YzXcVlNA2UmwUa44IVMZQvGbSy2YLUWc9lFEd7qUtKrJ8XyME3n
XtrTnE4nEvqLiDKhCPIKIeAdI1ewZe/aJR7net1D45iLBmmUqX1P1C6zhmov/3sj
IdEwDiy7wGNSYciShy2NaVZb7Pq1lVhDq9cy06uzQhwD1wvCywpduikyclx9lFxK
tKla9FlBZm2729CEXXvX88T7AhIE+7aot1EgKXsAPbshGjaPuBjwgp09NxmnugBP
vBLBdRyyKlpNr6hEljZVFVHUU7+wY6jkZHLD2ODO6h0E8QIBLvqwD7lJWLomnGHh
VpfyJQQcKzKgm9TXtJAOFA7GzAjtaUYKFLZGqmyACbkcOpmK1M2WOM85NATWkXbj
E7CfS0B5NrI1+Ozctaek3VkEAZ/hCxxiI5uRU+AqPtNk5a9DqPHPG1jsHdOiBDNd
2IZ4aS+VPsjzQcSlTvl43czs5PturnJfrzA8HAIKNRk9MuCa5nYYudVCZqNABBk9
sYm+h/sbWAJNhaVGpeMLHF65HMbxpTMJ1fSpvoYpj/NIJx32j+5+ySiV82ATQnAN
uQvxuMe0tiyD6A6sm4JjwVdJu31Dfckoj/OdqN7Rv9O+pUcFd67CSfxX3ZQJ5GpZ
Qro+T7HfIQz0vjoG+vLOGf8j+UKPCA6GGQxVscaMWx85Gjyt9rg0MM7R2/XCTRTe
7dHIn3GYw8S12yBvHuMsQ/DC0AHsMkuzuYgkuj7P7pyRLk0hN6DKoagIxAdMR9QE
yJulAyw/9mlZPnZmDEDpgX2R6HE6MSkiKrsNR+yE4NZTOlkRNSemfoliK6thk856
bH3CmQreX0ub+O5oO74bGhP2E6d/OnR8BQlyofGvbpGQSG4arHJaeDdK6I4M1TKs
Hob36EoZ1BUmOJtxgZAjGrUq8Lthab+2I4eAP/FqMpnKF0gDHRtl+mZJDDplKJiX
KzgmdGVZ9kTAwyJQz/GCOP/RTuf5PfiV9Uf5VDQ/tZo0HRJGfrMhLsk6e0lp0Zdd
oQ3819sxAY2sFGtWSnzEMFW1GrkKBZ7MeunMCqXADk/ZE7NcFAvuQ8IaUUvx88Cp
6rVC707865HEdmTYCj5gH5CnAyy8OfrLHEiNGQYTvxcnZVD18qsyNw5xMAjZcqLy
LX0Kx5yxeoGQhb+LXpG81m4zAzVV7L2OvY23FjG8wxcb+xOwJQdxPwIfNXNLcCWD
xCDUNp84h0pSR7QV8uAPRI/yigCTCnXd/Fi1xBzQ82cUZM7L8sOJ+FasWW7c4+JY
CxIGj8D2zdvirqofZoYfVmQm85SxilXqCizeVRZ/XhVb/c6kRb+ZhY9zvMwnX/QY
r7vnRKomvRLRshL7Q1F3MH9ssT0vIGTwkjXrvFSNW5rZ3UicInTViU9N1yTAV77P
7hmJtjbWLeNk2zPESHWJk55hR1FM4Y172yg/LzPh7PGeY6Gxw9cyeKdzq2KNevRf
tPEIlJJ/0SOUI0JGkU63lXT06jNZQT60vYNRED3jhU2tf8E3T55HqEsFuf+ZomrL
1r6vuhGKW4nBlEu0KvOr+pAlxIj2uFIwjzwCWTOboFfDfuR5GNVGka41cqWJUkfd
O9Q3SNvajkuM4uGk8CM6sgWc6MRrQgIqtjWg/urNX+UFBSjpAXTJx8AAvuB9QZdM
YslGO8/o1zHI47CSI4CrzriWNy2psaAIRKlFsaIciPBPGaN/JkYDI3GUlaHzjCY/
HKbB3fR+g1YoImjxbIaOB+I4OwJpMgOUgpAmGo2xHO128EdKwlhmmfCLpzdh8mut
+TGzJsM1GL6q8cr7LSTJgl0gFtQCistdHQMoDhAGI+P8ovdZEqmP3xevmJGXk67S
PvbWZUQLO9m/bauJEP0d/6QDCpKu876EgK8C63EDAoRD25fmd7N3Wz42tg7jbqao
Ez+WL0y8WxImLepw77YoJ63I6nqY/jBzMCcwXSl+6+ipJcoV3afQZWMirjc+mgdW
/qvrA4Vue3ATg6/5VuumQZm+VzlaFXTkPITnvyDEKkKKiNUVNOTuMJdqVNNVG8SZ
lFemtlrOE8JcMWKVUphvXtaNyiqFA+hXgC0l3MX+4iyLHD6mVC1G+umdgmqW4zOg
qPj7Hi5GAezZ/PeA7FPe+L61xsu+iT5dSg2wz3FL6suWFxRpo0KpA+z8JCH1PMOZ
RqMtj3ric1d6MnPH0hlTYq/TUDoIO1rfxjXSRB6rCfPEUShh1iInz440N8y1HqOk
+PylGPCwMwS7hjPQzU3iCiwYbKBqSNfSv8Zf+W26fvZJ/FnrHJwe5o7TTr/ZAwTG
7gEuaH6Py2RDfOXgPWQdLbj/IoNXvF4y5SGWhmBkGCW2AupE7Bu1wpMyTa+M5PRq
9d03nUxCnRR9EIIXP4VclWie6lwHsN5Gj0k04aNph40Pw5EPyvJ1kvVN3pdKUrNR
JLLm+RdNEV9UKEhXircGLq59JtG+MZ30bfNa73sREo01ldSwzKNr2LRm03sGayZH
Qt0aIeCa3Uk/gqUGNcCrzhU6aEybAoRgO6KTkTbchp7vpDLB6Fq1Y/hbg75oFRF5
gth4XRBb2IHoDbuk1WGeF0+egCXBe/SXwzS8Uej8agh2jmcQnL0FcOuz4k+WLVd4
MxisKzhr65lOKir372xdjzxZ+aOGmocC6v6BPPGiqC3Zb417RiLy1Fsdu74NJ1Ol
iaPNjV5V7E8TTWLqet/QXPWrPB4eXOB7W12h3gI00SfqyrAVSxKAy8k1TCy+kgi2
VlUwg2kB5/aMASPNV86TbpB/IprmzWu+HiQtDB+7o/cJdHxj5ji6+lPwY23p8/x7
LTYpCP/8j3jVpRLBD5z78qWrIKIceA6Tq+/8TIiE3tTdeM6ZzUI93FE33ZI4oetI
1rvN+mdPE60CAwanGDYVzpXbItCqi42NthTovXfWgve7+n77Ew+JK6MYACXGo4oi
n3D66/qck+jmmbbi7zni0oCYE0vYJKxf7fSLTe8togVElQkAAO0PDeMygPQla/rs
LWVdEmCWbxt72t8yj0JKTe1NGBpY+URX9Pi7qZAeGYRaOh7GnMK1ayrSnitYsI5V
CLbrFbwgUoW6VUbUJ4YxS0n/pvY7CyacspWJfzCxPCi+otpdvzd8bkOTsr0nQR3J
8OdfTaYZisjp+hsBUJEdZn/l/qQ6xFUMtXIJ2NoTGBNEJngxec8qn49n8xVc1D/N
uY6B8epejsAAuHekDMhjRfoj6d3wH6G1Je6iQiz/jw78nhM1SZ7OQiIT1fSIOnsW
KQbSmcTm1CLjvd1vUkicBSVAnehSg5D9BogIa6aEz3FBVIyGt6tx+D6RbkBL8UrR
ck6mwPix6x0d+ifqlSf9GdZF6rCgNIwXG/q/ja/PcLE+JlVd1u20c3E+JpKDTTsM
DMhjexoX+QZCEJkN5bMFYHY55b5qsZWaTwhcNNK0BmPr+XnMkrhmmWb1lWnJYRHt
Ezyub+yDB9nYD/h0/NGKdidcTCLBPf1JwUZ0wpWMjrS6yR/IfiDCbJP0EbGjHi+j
fLxsNVBjdxX4rWg+hDYwgiowiKUXDFLb2itcZr4miG+gY+BylL43g+wtxsa0ijhs
PlnsLDGFx5ppjGcVoHtgDm8U9M1MSP30AF86JEDRQ42nh76Wx72Hl0yf/WMlvT9C
AFINATmK/7bHTqIXwNMn5c8SLLYMoQAEChOwrIILfFENK51tlELGxSQOWg8k6mXF
5XoOaaIlSE6WyROLqVvpeH32nRqz21UB7yAYjYclBKjrp7Iz2h5vzsrSLldOG2gg
5HlFauwOxhANcrOcsuO6fCw6vduditSpRpEU4peFdlWR0hNoWhLFFkrWJMGUOVAQ
UGXoJ9U+t76INwLQy124+b1fKnSX/lprocyxGRzl2lnEsN2K3ePYh57vg7BbiKmU
CuUJ/jlKiSqUL3klYuMlsDjJ7FsNqL/MuMsR4oDhEqxR8HjBf7z8GtcIKxZuCSJW
iSIbdHFuKAUaIVOftEKrmpaAKFf2QzZPw/H13H/rfPrWz5Dblqv2Zs0lTMF7SCE6
j3v55ZJKDQlOoAiI2lhdpABsYSpifEbthvnvL2Zx4qwAMulDdoDHHZ5AmxJGFXbS
Kmcip1HCcUIJtyU8SFZmC0/HQZnpFPUgryPl671q8HyaTgIqsZ7BAVnyg2WTdjcL
6BBgDdBVmBIFx8qY94DqXtXLaosrYCNi5owSozsqCJ3FI7kukfj68ij3JmquQ41l
yBnVY/VL9Va1jHOP1Ins5GDBX0hTm3gtAvHjdgaV1VrV/YSLbdVmxAyrHjVtakyX
gBXw5mV4C09UoyZ2Ctf2+uwS51Qben9DQLWcpCE/woRTxRQQqQyqR+u86ODUJdzI
tiTr5X10iTiVM9CGIkly/EfavLiBTq7zTFjlC5zrXJuzSLl27FedNimgxNH2IE2q
RACuCcYlnBH72rUQ1D3ldz1rlzNnNb3zjcY9KKPV+Ls4NEQCSKy8KMkWkiDDM7v/
JpUuwCMLDb1dLHkYtyx1HRkFd4YvTRkFxoygVBXv/HJT7VimIq1aXv57LBn5WD7t
wo5cTlOEUwdjn2Nt2pJPO2eag796rrp0K5eVt4Ovf13Fhs4Ly9lV8WMnUC2v/x1Z
t4kqnbCt10wsbjOZQTrHXlalxu01W4BRrFFx+g4OCzKMOKMufWswzZTv3mvTGL3Z
79ov7pSiaxoDvztgYB2BCn/TEfumAyvWCx+5eHSon9WG2rYfgjezn7B0bkhnoJh4
VaTYiCAmnD2RMD/R5ZMq+Dtu/ndIvtdrps35D0mjwJXFVI6ZNrZMt5SKMl+uL7JC
L8ISjfs3PGgrUaJ0syFzfPmihpg99eMdz+TMJ31Dh/vJSY1Pjkb/nMCqoc9xrjQl
q8tTxCLNxFVz8B0c1k/bnJMSG/Id3eeDOxlh5aKOg5/YPO/r+EIz/gTpbtU7DC5Q
wuH7TSiH2yEmdGXqJsy6RkEpWCHEH5xMR1iTvhe/9K2tct3/JPkaiYjpFuFnapnq
ECetIkZnq5SndQgqm4I6vVTWdUG8IkLDKdlKGanyFDnx8o0Cxi0K66sGh709jWRS
5XnLJWrfMbRk8NsOx9HH79uRDKZoz6MPfmF7ngB7QPFBP55bPi+59aJqiwrrfVJ2
8fZ9ktuvYAFeVEPJjzoeT2NM0zLLzBnEl59nH5yN5ZqIctEH4lK6bq1EppHP89rp
Ppr0v9/jkUr77ZYo8uP8KN8Tl71o5tGFe8zTRNbUa8nM1cczEXfq5bERAI0OxgOl
XbW9UgT1NqbhCVpEh9xaVFQXImQsn1VCWlkl1jnHMurOEZDJjShIZSyGpQprtVgj
TsPvPz0CtDaT1/JJ8U8RHDRPFeADVZLopjVyDOsrn27uCHbcEVji+vKGpjTlohS5
JktYLOstMWHDmue8kE12CZ3SH19KML62t26e/u9aG2v20Eo6bWHwRhc1nm4Ddp1R
tJis8/hySN11JtnhGa1Xz3zyhM6tgRE5EfWdDZKtQpnDCskzo4V53kbpjVR6oH/H
obVx7rijeOGb7UBFWmpkKCg5Cdeb9SvSIOGRJENNy14qm+WWa2LYyDKrikHJVU24
SKpC73xc9MZRiKb0TUufs6zCGRY1x0kgy1d+apu4S3mn0Ep+mlHa6d8HmaOOr8nP
jw+evf2IVhDRwKC9hU8yhQNSBTxbDE5CiAOkHW5/iPGmfDC1rtbd5vSD6RoN97xQ
XrJI96dAtLR1XcaCp8FVk9B7x1/T1GaSNIjp2xqFnJpyqDAUoqr50kMaPbIgZ9HO
fToM4libREXFRMCR65tWvW2rDxMjVQnaHcceOLBjZBbJ9tHPjG1wS9eFZQyTfSaU
wMEvmS/c3Dm043RnEmMiov0xOdCOD7Z87YlzHB/9XYs=
`pragma protect end_protected

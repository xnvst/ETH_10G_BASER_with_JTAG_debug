��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO��smϪ�Ŕ[��;m��Rk_�6�T�[�:&W�O���Uu��A���`I�H�xݳ����I�^�lQ�������G|n̘��p7�d�>�V?�P��-��ӗ��1S�3�9m��#5	���1�]��G9k1�'�.���,����0�Q	�.��b-q�-���{�j�g�9@���L�k)Lr��O�f v��7���
5:�" x��>�!�� xt�m��V˨bK?s�J^&EUw��ҥ?���"!%}蔭T�]��z�r Ͷ!��ӕSԢ`���ϰG�^���]̟��:�~�U�d�/Ϭ�����F�l ߵ�=�M�P��S��i�����m}#|+�pX���!R(��z���R�?_�2lg��&�I��!4���t�ƞ`k�[�?���`��4fۍ~^ȑ8dH�h놬���W*���)�B�C<��ӏ�و�F� 3gН#�������#�@!��@�=pP����7#�l�*֮,���0-�al�0�.K�t9�j��J�aGZH����r<>�x�=����_�;VR �+���tS��1$p���qp�"¥�f���j�����´�BX���y�;�]	M�/�]��'�uU|�ʓUu=��O?^�:�e���մ0�
�ϡ�\��u��2� �Q����<$}��m�6��X�'ل���Al�@��~J��&��X��X���
\��5�ZB@0�O�fca(�X*�/G������4&./6�itPx��*��0s��W/�s��~E#�pa��5a"J��U�2.��V�Q&h�4m}����+Պ���#nn�B���*�[w�k!����j�lq����w�2 Ö
"
��©��]�'��7墭��j�vߠD��hDYA��+j�t�XR�7P�;������g>78�G��@��2�V/�J̞��.)WZ�U�='O6�~/wmd����6�]<p	4�� ZUs�Ng|�ΝD���+�ș�,mp�������>�,t�a�#��Xjr_�'��($&`�L�8�Jk��x�Ή_�@�)��z@L�@�� ˟��t�����`���TX���Ч�7Lx]z=��uD��\����o4u>�"�y�1��Ej�$��ǎ w>�<;���wL����Y;(�"\ɦ!�ȓt6�ܣ�]��^zC��ܧ�Hpj�*j�,j�aV�5)�������u� 궄�)+�G9���<},��;����Є�۶�̓�A:��}q�������ߐ�:k��?W����"��~'��z�S�j[%�p�+M�7�֘8�$�R$tՒ���Ѐ+qS�,5�/|Y��YM���؎)D�P�E	l�Qľ,��ڬJ�NRT�������G J����u��	i��x���}�vO1'686���!����,4�.��{�:�PTv�w��)��������ɻjt�ʹp,�F<:~�B����-l gO��^�u�|���S+�4|XjP�s������'i?��l�+Kb��]��<vij�B�ѯ^M��#���H Q��ۅ�ja f�d��K�UiO��@0x����ܟ���-�΂h��U'q[<��w)��D�3���m`� ~o*�Iw��Hr��R�h2�԰{���}\�4���'�E�6����lt2�=)5=;V1��i>�a�� �۷��}�t��?�(Dc�G}�/�h����H՟�F6��G6����~E�5��Lo]�S҃=_ݬס+y�.�G����klV���o� ��1��ɗ�l�	�L�����Y��b�g��K���\T/}�Y�̧[���t�\�<���
�@b���H��'m�Hq�֑H�6��V���l��4�*�8����[܉,}�1?�l�)8$
vc����SX�N�cl�����c���W40�����|q�K��Wɓf�]�����J���ŢV�>���_9��T;���B��¥$f�v��	�Gt�~��M`����=����a�M���nK�\G�V&�e4�P��뮕:�(��2��A����1��κl��E�5 u��������4�e�H^���tդݱ��/�' ���Hl�=��W��<�NO��ڎ����͞�<�4r�����$ۙ Y*L�
� 6�ׁ� L�C��q�X��'���L��L��O��	:h�2��A}��'�LV�iW�H�������hT��R�F�d% �iJ}k�Ĥ��+���3��e!��7U8L&���O�@4������t����s�KN�������#�,��̧l9��rȐ�%�!T᩠gwl����'On�+T�V���Z���EdU�$և?����к
��Y�����K���݈7��(W�z� ��X-�������ҙ�<=y���x@�<��C�{�����D�]�2ʏ�@��vM�lpz��LI]�e�m�é	-�<�x6ߖ:��is"('�K�Q�E�����4��D�>h��܉��e;ˌ�+͠�oK�4KU}��$g�.&N	�V���s0
�v�w���0�I��?Ƌ[�$8~��%?l;��6:߮'�������_�S�=J  ș�G�+�m�5T�	�	��b�H�C��R~���U[�a��//����cX���OD�S�'Y4����f{��~�`�%p�<��*/[��3;|�#�BO[�&�]-�5_�a.����8� �N;�%�ϒ7)y���ڪTH��f��IU隣����zwı�rQWvB��C�;({����.K|������'�_�����[��R���zB������[^��5ЎK��2����WV��j
���g�he�'cs�p��WDX�����P�y��[1H��%���`���o@M\"�X?,æ6���%P�@����������K��Y��	�Ғّ�o.��lS M*�/䎻鿾�Kz�l��RI�s�)�6Wn04�h �euy-.���h�ވn��Fl���Z|��,k3���Z�3mm�?��'�޴I�%�zEIW~�	�d�L����N�  ��d���]�| �*�q!��(8|r켂�����g)����,��?:Ut< �@5s�6��'/��zhg/2߫&��ƍW�����N����[4�����#�Q@a�RM-�A=3�4���rò�P�½�Kq'j��_[>F
u�n��n�`2%���5\;�ZXGq�RK���C��2
<��ٮޢ�C����{��o�@�"M�rf��b��P .����	�C>ѷR���l�4�C�	�%b[$�̧R'�~A�)l�z�I�V*�6�D��Eh�m��[ʹ+�mt���ȶ�q�ʯ2�Ϝ�7��Z5�T��%��eA
G�C���#�vV��vK�r�7Ҿ����Ec
v���*�yn�û�"7+�]����D��`/����Q�l������9� w�F<(U�ǭy�V	E�2�Z�%zc'���Ú#��E:�����V��
�XY�x���,�Px��(�b�۠�/:�!���7b]	t.��D�{YtҊ��Q@�p�I�	SA%�>�Y7D���V�}3�ܓ����>��*�c³�Jg�v[nU�|��/�p�W�36��XsI��o5��.u:DkA�nr^�PthٕRqv�ϐ�r���Xi)ֲ=�����bc��C�	 ��j�K&2�4�lʝ�Q��}lp;@�948�Uj���,x��jx���� ^p΅'���i=1��þ��n!�<R��vw6�"�{|���h�ӏFnl(:~���3��=��?�1��T���{K�:?���G±�k�Xh�"��r���`�vlay�NP�P�@����a�5`�Ԥ� �)�0X �&�C�F3I�~E+���X��N4o� P��O�7���	����(��dt
,�N}=�U&��m�ʸ�������e����*H�ik��3�']d��@��4����J���:k	+��?-�yLz���L�V"K����_�u�<C�ߺA�.u���'��4\�v��Z�jb�5uH�v�(��q��T�u?�ԓ:�h�4^��G�TՏX�PN_Ϯ��S�S=��OLgXב�<qu��k&鿛+�B�����S�<��G�>��'��%�,�� �h󏺃u|��{=-݁���D��]V�������X}�qLM�2���a ��Ӽ�)w�$n;4�wj5�q�Ú|�,m�H��R9���j
 pe���s�ce��B�Ǻ�h>>&�MBb];ո�E�Cgd�;r�ʾC37�� u��i��1P��_F����@��*\i �*��),9��`1�����v�qP��{��\�߇5�T�C0e��j�^��km7�Α���4���2z�=�9%C�k&/�o��{�	��E�1e��F5P��T�6�%����R�tW��$�>�f�Џ�^$�S96X�t)�q���&/QPm&��n���h��	��2׾(����^��Jp���)��A��5�I���Q�Ԕ�p�V����Á��3�CFl�m�yG�8�������Ti��B4|s/`0I,�R��<�Ӹk)9qE��w� �7�Q��@�lT�&��F`A㦙�����t���>A����)CQ��ytM"���VT��@��<�~O �ԶTp�9�2l���˸���aC�gAG���w�H�z(�ÆM���'�<�fxe��u�h3����t;㩘�r�Ɠ<>�v<b�Gc����}�M��QG`35��H�u�A͒��B�˺��2�{�݇�Iu!�G�I�Y ����t���^�c����[;��7����s.x�����蚫t�2E�x���6;b�ւe΄�V6֤�f�j1�I�����D֪A���Mz��9� �袸���N�[���� .����������ܨx��<܎Tޮ�M ��&�y�vm���14�����b/�8��[��z��j�U�z��a���@��&N��@��Ot�w�LD�!nГx�l�����E'\V(:���Q�`!S�8z�
���RY�Ĺ����������7�)���lŮfd�}Qڬ��q/z�(գ�*��5��ǩan��ay1J(fSJ>J��Z��}PE����i�Y"ޚ��+�%�L[�ܡ��6
�P���m���Y<],Q��x�>�������j�WL��uHUa�nA{�g$�!Ea�)��L Hh�kB�f�O`j-��{(��<��`Q�\q��C�.��VCa ��P��L�=7��[>k�0�ģf��ܠ!E��F�BwA���?o�#�aGx����t]�n��q)���J�Y������~V��a��Q$��2���47bE,6�R"�6����
�6�!M���z,	^��{��7���m�{�w�3���e�1��!3b�缻}��<~(�T�P�U�F��<�k�k��ҋ�'�7�vs�[�fc��Ey1z�N�Vܸ�}�8��ST>>���4��­-|�����~o,�5m>O
�`	�YH���r�����C�ځ�7�B ;3�q��<XQ�d�K��p�'A#h��#�/�C�?�G�%��v5}6O�m;�;���i0��XyI��a��[���b���XK薝g�Q���#�"�9I"��t-�B*skV�/qA��6��������#C��(����J(�4�d v>e��t�M�*��
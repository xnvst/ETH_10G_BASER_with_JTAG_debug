// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
TkhuxDIjEc/RvpRo4U+hglEOTf12VaZihl6ijkmyE1hza6RRMcCNMjuKefZxXMRA6WyHc4WDkXTG
Eri/c+lKqQjohPHne/MroE+m76na93r2dia45WgNwCAN9RX4MjQLmAs3yK9uuin+XFtt+e6xXde0
vxfIThIk+PhfXYGsWPAnE0oI7zRLAohvoq8MDmgvI4nJoVbag8OVVh3l8mC/q2TL+rZH5vm0CX9k
9CmUqjVXi/ZaugbE3gP3jPyzlHi+kg+O+LKPaBO5cf4rwF6LDq/d/ngBmekwLV5VVpf3eFlXjydZ
GZesPTN8DxkRL5tRc6DSOOOlLBfN/d/7MPXwdQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
nThRAjmZ2vWRMOZaWZvR96Kq+PlrJBFGIvivfZNg5aMIgBF2yxPlBsklxJ7CoAx9CU4tfTM2KVQK
n+Ot7L8XJ5QPdxXqWCjQVQKK5oKkYz++A0b4WLeiAXmHvOK/Lx76wmQtRn7ynJWfE9/JnXHOccbM
mVbvuivCYDPt+QNsCvDWKBtMrzbyB0vAoykhiglTUrwnUH3PHY6Pa9tZ43yCU5MKLvcTs0rDYqca
pYM2wm2P7QDv+klqKVHLN22zMgVQ/hLffDzgwe8bQ99y7Ow4PTYQs+m7BHpoWvCtXUrpTyI3EvGX
4xc3X501AkNyesJtdRF0Tq9UX6L6RWxit7BvoHNWRU5gUyiYHT1r8T+Is2/fxj3lLyNNzWlbbf4Q
ah7S6vmA1fOaiWcuBeqJ+lbnmAAlfIdCfdl+a4i8S+NSx3IeGHSDwoSu8gQ4sIch3h6K4Dhp9j96
7C3jzn5y/UDyVat17UjuUtdqFW+k4gDRsVv4GnkjjPtjksjGn93DOniiiUqd7xSQm0MU3wa1VMCR
H8k1r5WTYpSFMtYn37Hig8xUQvly71PTAlclzSjKnJqSYj6iZytogP91beFaG5mHqwJjnKZ4rSfg
S73aEKFVZ1uX2IQieMm2vDXLY/kO0RQ7pJ91eIBCmtohZ74gvnbJj0rrvSoaljT/jYRsMa9tb2eC
hDJlY0SAp3Xx1zpIiCz+/u2xA51jE0rp57x0Xx6ym9DMNJQXBKdslgmgcjdJ68cIk2Mf5zRepiLs
/StCmdGsEjNBEeds6VMvFv7vCRln6E9mHvwa+u/BBWrDuQ+/gL9hXmU8PWWWQkYOiklWYDTqL/Sg
yPC6t6VPzm7TSmsLzznvFiDl7eUipOASAPEy611MGJfjtLRZJ2pWUFgKhl7fHOeTZrnBwjLBEm5y
pKDyKVZr0umDui9TeL3GX/3ww8pj6enijk8cu0gy1KoWFllC7U8O5tciEAcPqcYBpN3Sn2hNbbeU
y3ZRq5aIXH9zW4lBFr2qQ+UpPojuzOqY25gkv7VTkTuIx9Xbcv2UkcN84VR9wycTqbYBuOC4pCoz
VbVUoy+Ub506+l3kZxdJGrHvWqxi5pkuFhZ6q50zlxGMLN5GW2u5UfQquSvl83xXi5M6yo6oSsDK
QtPdkJ1OkZXxDX6KR/zRtdDm2ycMCICvSfJWZKobJSw2FEDW+haHmnZw27ralhH/vskyOBn+EdsP
jKRbbUu8Kq3owaTccAKbao/jwPxlXF4Wbtu7MvWly4rHIP31Dm5WrGeBxtXeEVbvuDVfHYxDdJWE
e5xxwHNxBu6Ljvz+6KUvvQ3Qse/x1amufhpht4fhGCeI8CIlgiNljqvf2tQV8R4qV6/b4uO9XAwA
7P3ijsVCZxGm5uX48Z8dhjMITVoJpmx2pumf8Kmggzyqwv2lub+7nSZOJXL3jwvr+HN7VVvF2ol2
25ZgfshicIrZFNdybhrfx2mzEqUIOJOaQsHGpTkD+kOLsv1LpkkFpr5W+jlJ3NAljHNVmow+93yU
gFJjkr22lgsdliu5v75sFxtOgdSRiwVTSV/EpwAGTSAcoWuHq8dFDdgbWD68oEzFHSFU5XOTTRty
VTFNNGCcUt65AIEfWIorHR8nVtaZhGQv5TpUgEuroZbloFUB5XNHdtQMo+Ti8hdP3N9Gi6vK+gkR
Qb48g2IL2PstjpYLnW0pT8sguJYoxV7bNxo/L2zfNUkVTgQzSA4rn/ZXzKrQeONAAEdm4j5E7NdD
EwkhCuYkYZiagYAvxwhJsN/iTzYa38q6qY77X1tnTLl6v7YlguwBXJ/98IWis99XaNzfX8MJXdEM
O3Yln9XHI+LYIYo30YUIhT5BhVnCtbHw1ZrMF98f6kOQeZy3mbij7mXsQhfOmGGDx8ON8KXPWBUU
BsHPvuVnrVNDrWTZ7Z71K3pTAntxe6PtCk5FA/zV9+HkVBuvGiQu5wgu64fu+hzYpeS4QzTXXK4q
vGFfnoycgeb0EaFLGo89SnVqP5KqLQW6g2nyRZyO+TzB4vfZ+XTOqVu8UsDTGuDxv+UJozORb/X2
mmqmftZHg3znWTd08VQAhLJ5It0KIwSxI0/COWq6d/87kbSd4lB9Pz+2Tef2cn3+gj84mLnBhihq
Qb65VhGCDbl9SeE3evJV9lngHruxbwKsI8ZMQNfEk7dQCsTs+xUWRe1qpAeYv37th+ufk5vDYZkM
tPLz45aCDE2J7NL5zajxLzzA0cQhC+Bar7wi9MjOpFueFvOgs+RHfNM72Ug22bh6QUxHbgnmcwC/
Mt6irxBBdvnyCQKHSIgL9cYYIprtLTAy4be7uAVPrrvsOOoxevX4w/aKgESNDOqSepgrZUxq8MgM
WvXBWaImL5qz+bgYCTlauWFqh3y2DlcFhJlXF/FTHFL1GdYjP1RjFz815xmVCgAf1jeVm7YG2vHK
bypL1nAk3nll1tgJgggyI8M6CIlR+bCSPJT5YSL4sS+EbjIVVhLO8FuGT/jmcBgSy+Ajy+4pJ14J
4X/zOwTGK6eBLLNLcFRw/GS3/5kWZiBxhGYESwKUaeioTP3gmR7X4flj27QfE11BFqmuZRT5AsGU
5FaLO7pZGyVOj6lw0U/5enVGGwaclN4bEChHk2xAG0AujXcYG1bNUQvKF6JqxrqEpuKxOLxHZDDl
DdtSOEWlvEIESEBBo1ZXFK7s27pU5xxrKxJFfQsjR4NpMu7JMMd7ym/3GW5UuPQ+fiLQyIg5eW+B
981wSWV6RZfl7VzcyU/ES2mBZMkCAZKmH8GG0rn2ieDmzV3eRtW0lqjeiWi+RqgUbMmolZYKJwoj
bIVh58z3ns8n7VhQx6lrICvxivuXYjLMeYe2H38SEktdYWF1H2GZHRmXONUg5rS0UKLHwzJbNLGj
waW0LSwXEpbQra8t5vV/K5pyJtU54K/bE430GZAckZaq5LvJfVzJRcM130NO+zQm/epdcrJYEanF
X/idQ35rUnhOPgmx/0sKDviZGNbbBJ5BUxn/y/NTkg3IavCWIO8RoeMtcT0zLGBiy2gMNDn8L4cD
0beAZpMRDND/F9xMXmeo2nhaYQ4J5s1ZM8CQBHmTYRhvyishb8+b52S8/q2Z9+vVjSgVzQx5mbpT
jzFMKwOJRQFSlc6SoocA5l103Sb3b2v4y0we+GVhS4FXJdWzXhtpaFP2Ph02s/+eRtYgcFwr3gun
iS06db1YMj6461OudZ9f6Z+/YbMpOJPJFekluR1NdMXnj6VZYZS/F1f4HbdmQ1xlGdEesOoZISTK
fOqOtTBZ5kC8foJZUJFDVGQalSF4C6UCykr8JJTZTyKKUgM/MateIuq8yVidMsUOKchHceQ8/gmY
+fbembyAX9wk3WN3/Z7lS1qFjdJTyeM6OLTdp1guD3CJ2/onrhDL2rWQypP9P1W2/iSDKlgS+9Np
JPTOmFDx4AIdefU3IKmugZTJQM9KLCOPOwT8tsebeBUbvRPgyPvK7L/lnartxnBNYCjxPAjdo2YF
x9DueToJvnj29gzdv5Znk68vumD/09PZ9acCgSKJsXXugUxmpVwMhdsGGsLU+8tr3yyFT4w9YOZf
gScFeTiuIORo0cskOSgd1Pm+SgGaYr9bhEddrJjdYU2ppfImqbSU64bpITA+NbstGnB3YkoU84mX
Uf/hqMLdSDnIg2hJm/uKqM/tMhZjRK/qoyQCH7WwnmiYeptckDb1GU4kPuEpPPMHAjthKAMj+MIR
nZeQndvJAnVcduJCQZDISoSLSeE09RU+yDLgDSQ+0T5TRm++qiPtJyb9uWdMXzS6ivS7GVkJMb8C
PvXfnDUkOcl7vFPXgF6FkjZKfoRckwAWzi/8ZFrCERnna+qxV3D5Y1SQtX9K7qnDIPtvzkukudfv
XdtAUJFDuN+jPKvuIbpcsj0CmW0uuxHW+v07Gg9HRRjldnO5kl8cGyTCkptLzFiaUjpFuFCmkX7Y
HKncMAyZlM0pkEHwyiwIbcvMhL7ZrTCTPHqCKfOuVC+wHu1YYbHLxQspVqBN+T3xkvV2yDgOn45b
VR7V4grNJ9weVa5UcIwzjN973oUnPP3rpHtfLvIyoHhy2IZdowjePX+WaY46Zwl6huX4tMtC4lLR
xMk9LBS4uO3DrqznjxHUA1gsY0y6KtBM+9m8TXXJY8oWgg4Sy97fcRDaMG/pPc5jYZJNgG32OWRX
Lw0BnJ0XKJ5GTdwoXG8Ydm6MBAzXUBsqw8Tkq1GCV9nJ3P8RLvTrev0yUEJEO4nd3rhSnqr+Fj6K
gHVSPZzw0hd0RvtSK/cibKgtjm0K+ycJFzC/FazwTLZDs0yJhcrm8/sVL0V8i3T6I2lmAJfFUpqx
yJT2+L6FvbDsUy/4yDPBeQsCc+PhP6Z4sBSeFa1JCfgVrIggUkHmRa+3Z/7eGaCeh7r13M3OyoSe
6H0IKtSTwdc4tLJNHf3bnX/S9dfAqaiLWK+5/M/AyaJqsDN6g/Aa0JULsjKNTBTBU14LeDVik4gj
mWYSYvJDFm9zFG5EtZkFV69AE65jE2bZuQVmd7jCTVgOqETNssHpmhGPWjafsUcQr5DFwdojmg2j
5ApyUeoVQIN+5O98sQ9zpcMzdMIgz2kiJCdNqcRyZBS/WD9bd7qspBoDhnBF9AC9Bh9tDEmz0QXH
pYeYh64QCqra+eCoduqMuH0hKmXHSo3LO86GOhpBRP6LnR92RFoqUIkVaDxUwWEcTXO7xEdE0bHY
irQH+B2nc4LHm0egyBuAGEWYERrFLuvaeUM5tFDThWbixx0SAqLdsDCrF6Pv0wpaegHxq8ko/JmT
Q3OFY5oNcaqQbsJdBh8b0b3m0i9G6zTrmsX25+NBh3hA3t6D+IrGw6hv5Vobe1D8CXVEcCEuhARX
ySZm5dVExznIzmObTw9DxZcT1Qhc7H46xpc51YVhYiIo7vLv/vYJAox2XkQH4Pij+XiSWGcp4NDA
IxZTM9piulgyde02CePZJaHZkmlklmjzjhESPFXuhj65BMMALKsjiagXmHRTb7CBkN0e03ACa3py
3svjik0EudAUqso5M0vGEN9BhUXA+p1SlslHxB0eOm5Bsl1ehAiyYRPQykGA1N2fGPzgyq/tNVDc
V5rqI+E5RFpIaHSm/2sDbwsqeQgKLi6vCOmaE77CXhwlQRW6BTHbwGu37JfZl+Zr0OW1FiROG+AS
NjttzHXURvpgVL1dymyDWnoBWRaMmeO4vp5LXLu9NwYzVeU/vB5uR6lbUsUdzuDto4Dkc1nsFQu/
xX8foiYij1XdJlZPWLlqrhEi6eJhKl28oyuW5BjpPYDEoJGokZxCLlO8zPvy+eAbKdBgUtl0jfgV
wMMovoMDfmnzibaXEGesshjMs3SGhjY0APtiyMDrvm+AU5QGZKyVJ5XhUQERBr1CBSHVDWLY/MdI
oBQxIkbrnKspDmUmuAg+SpG2F0ahZTkx8oZSFVR5QPHWi2qmG2Bwhl/Fqp2hY6e2iKDSh25Y9FM1
ZDpn4DKcHYyMRPERHfX+nxhyLNADdVSHeMaN0Vwhnnrijwv7vm+0bKPUVj468lgR+7gFfWJ1ekUg
atVBtIi7vHK5bSOeUCdhZb4xCP8rwf3AWj47KfXIQh+P8N7uvPMSNvmAkWHHUXD1/ubBuHr25Uqz
iCY1Kwd7BjQuubP+Fi/dKSgV+NYTVC7Jq8CIDtihBHrROEdJKZdS/beIlLDAmUVfzhvHHB66eBT2
5i6Dy4SKFJjfKte/Abk8iyjnvD9Gp6brDVCtiYRzh8EuKhRsPWzKyy5G07AGsZuIRYvqeWy/XluB
CulTLA==
`pragma protect end_protected

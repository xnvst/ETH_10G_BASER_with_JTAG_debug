// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NNcisgXuP8zftM47s1evZUB1XAnYZqW/hwKTLvd6hZoWH5y//Rmon4/qLTeCrnjMTTbE24npcSPJ
BmkEG4Lcjm8evOU8+GhsQ5J3GJJrvnFgcZzU0Wcc+o6hKB3KpPGqwvaNvgLVL48X1E4pnVEIyl7y
vPpzqWDwrgyAuM++CCC68UVLOz1/GU80mFBWAFLxxy8svLFHz4IR1Oas1sNJh3V5R5jwZDDE8F7/
/UjuwVgQl4ezTu0TujLTj2iqPpo/+xsiyRVfIq5Xq8ybSmE4Vc3Ow0Xd+aOU4+Ui9/ITa3uJuCnz
TtT0Y7LQCiCUqBdKF/NQs4K1g+kpURYwLbqr8g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
7ppauMWAs0H0mC3PdADOr4xqEozN8M6uCn2NEZ3E5qeIqwLBuXzMH7TAFfKxML9ftFukTv7sbebn
MSFgRTzcd0hwuGzNEOIqsJkQogKkAkL1khSDqm5CPKqkSkussX7xblqv7LK1eQmtmPbfKbe1z42O
l1VloClKRQS2HCbwn9lLOse7uzil6nyl8o/v36kSC2HrTyQUd3liylv6cUl7XWjDSaSB8zQHFsw4
2QvGjQI30FjPFIMNRumEmEgfVmbALR+u7wEQkvz1CmrfOeF4I1zwY2OQy/wedf63UASEbyP9hRvR
6ULgGPsUo2VkZdJjGu4LhFFUPkxyiv8Hs3DXkBbqPE5dnk5oef1CSpWmS6wUoNTF61xNYDwYXOWT
RRf0p85voenaahs3OEIMwae2rf9a+uOxLIKL1keM0Wh5f0s4L8xLSMEtdO6ennM1OIPOp+fEcnm2
mLKZdeVMTj4heMMdUx7hAg4b0jfcGG8pp9CPLUxjajlC4sA8eMRPBY1KbsdjlC/GkC81Uy8toV0Q
EXlrLfuYcX9hIIw4fxY04f9mY39XTPmuhHaJAMQG5v5e1yXxSpEOmqRtDjVhtMcHC/G78n4oH14s
fu11pVfvZaUQrN3kV3STuvZPmZhTj6sYc0NK+XGhnVtLUXHoIa/hUcnWoFDXoQvoR1d1RPzRZAxQ
iACtvCc0eCEUIn1aZt5labDzOgqQDPYpQVpVRi84drecObv3eUA7mVE+QzF3u5Szj3Cw99hidqUe
6lNldSMYAP4q57R3XEzs1NtscbOXg2OUR+Vw6o+V6mIUNRCTno3SK+T0v0oTLrgyATwCmYDO8lQA
0bkICIQ/iKtLaHlziEHMWEiSgqxQNLPs3Lx9kiG+4HMuzeUubUH0yOgs8AkFNyZ8c7Lyqy9goyD9
dCcj5QYg53sgK24dGbkHkP2ZC4/kbY4PuopTkAa0VPUj304di53ptkPDsSlXDLngTfc57PAXd7B/
YeP1yfRuubwCq0KYM/COidahiGfulDcy3oObIftNEB14bUjm+vaNIK+2r52IyKdVQLi3xaeauIUG
25vzGp0TC0wYnUVAQxkNFQbUMCkuUBsC/r906Sryc/e/T+wgSR3i46iPWQzuiEqz3+La/7XMTLgN
O5mCt++3pbEzdadiJc7Z7bwRAV1n1TjA2KxD1wkM7cnfkYSAtGs1TwQ4dkGjTAZ4PGwx9Yt8vI+U
zd8XpY426JaHLqrjYPuCt7jjLq32Hf744bBojwXniAe3CbhbU9xwoLJ24DZnEMSg1Ok0T6ikuO9N
C6Tj9RpfDWtr2rjZD7q4x5KuXqWx2J/wmwwNlYtM1H+nsXUY5TJIQKadn4vvxt1Z52ZrMIt0i4YO
yeH5FPg+lxtYFdFV2/NE43ufxOlSK5tcI6U2dTsYGKu0CGYCvopPoM9ieIPaSQ4wuMnDf/bg0oOu
BGZ44g3ctFGnwOb644il2zAq6bq7c+UaSD+SZ2QJTPhBSEFJMPZ7U5GnFPFOUU/BvvAWTv2YnPs1
cXBJdvxr0v/PDHD1YwBtX5GyD8xjj9FhXBSw5YiNkkQJnif12V+XD8Hczkx4qs8k/hYg2AJQ5Ne4
98fVhUTLSXoL2u3yFltXGYpzOFc888n8EvefU7inVq8x1BqN4FdAPbkyAGvzFHOOA3+lz0qQ7Lw2
030xmIEoAKUBKxFlUzRnFoc5ZopYXwFOpWYYL25rHaVaCU0FoCIMQs/DUXuEGIeKZU2EshrJ4nX4
R2VTqxcI5k3/LJE/1h18I7rU+pbf75rcO4q1G5OsM4JIGtpgCU4c0Pw4TX1Nfa75R9nYVKIjjd2n
qQjKjaYatMRwjrWMNhuhj8zl6/IE8/jV3wb0wsPYpZC9EBvDnn2lv2LzvUyWSZ/+b4eln6+RMQbj
r5raNMcHvgAMLUNN4Do1vN6o/yNiN4JZzknBpXx0cYURBdqwSo8ZqL/2Q+8msE/xP4RYo84n15UO
6u+boutk2uPkp1aDLoVUnPphXBbSkacHsuQgs/Dba50ThkfuP92jqCUq7CGP/xPMmb2OJvizOCGc
tCMFFicWRPdnexMJZ+wKo5VRwkqqpX06AuqUJthTTi7sEDLfnO+UbjsDkkdIcj9ANG/nfn1Kz5bR
o3RmGVgtNS8mOlW0+7MI/ipo3G7U4+i+sRzSESGSEod+caSkmJ/xaqvqyTQ0dDZj2CGG2nMd79ns
8A08P1vDxTOAepnJzM6QEdvBxdrq2MMUaMrELM4I82U9iTzPbVfVZ3OhOqFSoFLX16rBxEJQzljT
fxIz4Wu/e3Y5CM3Ig6JztHbxlrlWtEpd/RCWZm3SkFEInl3vZq2uGQAIMsQD1FkT8ej9hHA14gk3
iUAz28e3cQFpSoOJsfetYkpES+JUPq3T5YoQAajO5Pa+c5lxwg0vJozOFFpvh+IJrGH3OaMG2KGf
u2Gqz6PS9DgUZJo8IDgXshhziL9q+UASplV0+PPD/draj2/UdBXkL7LA46iNF//L8/T8/U+8RzF8
4qjh75auqvs64eEQXGdx1Tve1oek/9qmIFT0BfOyCwJMfezRy9l4EM+arvxuCbwruFkzEznbs8QL
gkaQQ0MrShsUJmNBT6x5H7i6fECnqhrb3muGsdKjpAlJfBP8qhrJ9t9UF/+CDHwUNeo3xtPgWShH
usRMjB9HbkSAZTjflM/7Sl8sckYs6Y2MuMkhiQCwafK9Q7YgU+Z/he892RwqZvpGAykQK7ElbSxM
MCxhm7m8Bp7THfgUsrOYg/DeACkrz12FuVMHE1w9+RLieTvVdMKkTJa6/eWJtxG5l0vl8N7/V8Cr
NbWrJTXV40PooPpeXDK+VaXGEtrqMbYpZ2+eRwojdT6EtZGxizEAF5vtGg4OUcG2VKlCOjPucYWE
lIItOEb7vhW5rcaD5vg5maX+0SjKfizjJSc1swvUnsw2PPiyErfZhF3ioOPqcVnkM75imH1DwiZC
NX2sL7HOccbhHL769QKPjd3dR6GZeMsz5zGpFM9xxNOlqw6s09oDEX11uAwh8X21ykP0w1Fpv1CX
w01zr8ksKOHylhAQnI0QUDC+2y7PQFH4TE2W9BCDfMfjRIuzt9Suz7WlAnex88l2wRiLZsHpvOgG
sK3Kxggb9EKl/GANv2EPOt7OK8HousmA/NCSGtVBT9em8OnymZJlLMISwu5sNrl7R1ULdHpXIrUt
yqU2HYguQ10jyO0O+ZpjHT/KkIb6dC0WwiUe035VO4LknByUPGFcHY/19g4iw6O/g0s3o7wSsjnE
ErBHumRMda2CYTRdLl6Vl9feTwjrqXimdjdke0PzhgCbEjSscwaQsncpE+DRoVvgtJoxutBzpPnr
PEY7x3H+MI4jhkc3BoUvxzZ0hXDgwCNsVIDewSkm3A2etYRQkOJUVi6V1ogXng3Tp+DYB85pwZh9
nSz9RbovB6X7S/Zh0NY6ccWSqixMWOnXKiGg4bl0Rz3T4dHBfzgmgaRMVIw8w05XEhrMOTHsnKSM
dNnXgw6yisaoaKk9/ZhDKVs+wMwUu0CZduUTgntPqzvvzeDuNL9kLlp/XrDTWBifNY4ziR9hnyTN
setMtUmacqxwmi35eaoz3x1k74xax0+3/etqbXnMXAD1eB7j1xnjiuRMjWVS+O35wOCep1GhAlNK
9QSq8KLojBILmkJkrrBtBlBH3M3rB8kh+mmVYhGhYDiI9rqlNyvV6B9LokVfd2F0/ej60wWSP2mY
WrVysh6aiQP3OBHJllcvOh2xkjjU+aofCRzxhS9P3BtVji49N7JXtvvf5Td2cZBvSA9Wltx6cT3x
yYQBGthVuB4GMUoiV6k3drRqFNNdmbkn7uS0MNt00MlxMHIleERJ9gj5dw+9VASmaccc1khpCxje
z1LRVuIfoG8DcYBG5LgJnpZim/dZvlIPLUfYegf94Q9n/WsuWFQ2o0mL9VYO1C6mxplyFL1pW7h1
OHmm7mS+TMu0oeb9wofv5jijNLcPhC6dU2TmLOriDbyXkx4tNomvhYnNC05QW1Af3ZsFB0/PZTma
YkcuSFj952BU5t8Fum3W4IKUgnakNXMqH9SPNP3ZzaC4h0jmY+6/HCVDFvG1rSd5czXDtvjgWZhF
oGyvYl+rv0rgW+m62VLWAJu8JTv0P1lwqoLxYndkEQqT1gECl/MxrdM9/Y0jfUebYcutSCONKTm4
RWEJAJGVybT9Q5qXOCJCtewEh38OLCyP7TXgldNKXeKuvgS3O/DL1oKFD0hJSrzUbg4kM4I4LR5N
wrIDY2/LCWzk0WtSLFYkZmTZaOWWRt9r4zk81H7TxlogIz2gNVnb8a4spdP6qw6D6sM+pg6AwqFD
uBzdE+0h66ldxney5EwUlSKBaKbympMJ+4HCW6Eh4RgNQj0C+bHvgePDgPkTEsswQex+9xlklbZC
0LTsnmw7hApGvqJKnHXUasjrusCMHk1f+LWacHD2FFGsAPRxZea/cXIfujB/mAGArczAyyyleXTb
P5EDsZ4OoPfr7uxx9q/pWynLaYd/Nm7mthDIgEN8kgTfwapWVAvHDDzl/rsGhMf/WdxX0n0SQAxa
N7P1X9kf68Aj96luS63Dbo0CksFa7TKyRANr67SwBTSvakMLF6PtCFlzeQ4X8bgx87gKgnNjSXOd
aKbuTXNSABPcIR80ZhMrtkttYz674rJxYXT+XGGfROpHAuVXDhM2/PgKp1lmNN7SGmYj/pEXPmz3
OTKH+j+TkEI6OSF7yavBqU6nrOWMJTWru+tT5UliMAU65uEj7k7DSgjTvzbhmPTYv3EDrBgENloz
Yjz5HKVhA7haJzX6n1SoMdLj/Y1Cw/V2FhYn13fzdz+qDKxL3QuzWKs2mH2jALKerl2KA2knlRJz
A6ib5IoORx1Bd2sEttngIm+Txel7iomBQMdFWA8lqcat9lpOVtTn2a15fAGNJUPmneLKDKgMdqWu
3v+0GDznbBMUnx81G+3w35qcdirPB5m2AdtnjfmrLFDr4bG9lPNK45xY2gZGbR92KjCFJtpWpOjS
FkUb6p89x7jaJhYqjy/ybL4shSN/6+pTGhluYDxffkgyqwH18TbrQWV8VQetLJ/nNkNRgT/XF7po
eZmuAjJOBKKpbEcBp3hm/Wtj9s8+FBlOfnIU8u0lUz8rHV/5mGnuNPIIU7UcFbHveF8N3A+2UqfH
RTbAes6cj5AkDuMuwoUuUqYJDAnZetTYTAPBFL3cAN/Z+flMU1eiUjJYmo9rVzKvSfru4MmgP9hJ
NgMUJZSMntu28WmPrx7LewMevAqFlmoKYocwWm6JODO0hr30EpJVMQ6wwtPw3mOwThc/Z5sWLXF7
hYskwPBIR1BcNNR6gUieVej2cH898c+EjTiK76xD576R8l14NQ8wJGkpj/SzIfbJnH4BRnW/ITdN
rV0gHjIbbN+CxKkowRIRQnpX92SOduEYOK7+1SljSW0TSXICRrX+BV1UkDlsH6hgXd8+/UGtZKsu
ctzilOou/1IOb8AeU4pk6BT+MePMmN1keHl0A2Lu8zhtVx/iFlwDGPGFtENbUQhPkWnQBotA/9Kt
dlXIByHRRlMvVBszBPXYua35iQkbYiTHe0S5hX9q/vXSQcW63kXjPLrhW3XjcHJ0Zctu7p//gzSz
r3arwlUWMe8qFQMm7iWT2tk2CBQ8da1+f2ow7livY2O1U4UQRSRnkLaG7kX0MVyFexrebHZ+uRi2
hTJVmMC7K20GzUHMtcm0dm77qKT+LRhcz5jzwSPmCyTyoLspi36U2gw18zjGfZ8qvSlzH5hCsJ3F
+qY+napvbZXduWgzosm3Dr8yxq8kxeaQRu8WKD3IRca0oduiDri4fBBXa/XIofKW7ybZAy+8aYXt
jNiiLwvKd7fOOslCwvu08rKGNit2pNHi5tOI1ojVl10HUYUJsLE/4kc1cO3bxV/t45nNT2ewwsjO
3U5DjE0BhxsHLfu58n+d3aB6spy7+VkckLGBwlTpsboYoEs83vrhVi0Uy2i5BrSG7Rg8mxqMLh3F
DMHeAykHSBBIqWC2gKXnVl/FNWt4jhKNAj6t2PrwfXEMzkYUL7rQg83fSoZtnoo1Jtbb6lX6LLnG
UNL5Gco823EX2s9MVc6s+3FC2doheTWC+y/CawwaG0eW9ISp5rQyuv94DCn9whY4cwuf/VTX8Ien
6GMoGGYW87nyk+2kZIKPLJgMjyIOOWJ50f8ororR6adDDeZy9KfsvDp0OPV8bQumFJA+tY/l971u
EwVlk48XocWeYLd2rSOyeOFlEQfQpO+KgcHyMPfRoQ+N80CBLSdL1zH+tZRhY0MZz4m9ivTaFNmV
ABbu9776KEP5/MD/C46Fqfgy4gawlrWydDK5D3qmzk3xy1t/hGiNETNrRs5r20GBsS+eBPGP4jFQ
CHXW65wv7vFXmVFHALaRa//j2t4OOcZ2b3oFBQIy4VFxP1IYAhqZcbhqaj7UtcccoMwJyA0VLRco
mFPmbvFh9zxG3m66p1JJYVDZ1WAPcXMCNOW+XZKmLwGfy5J4Dv2uC06RtWvDxhXDa5pIgL8yU33v
2Zkq8VpL4wZX7axG2wOkcPiuDcX7Yby5cm4tv4hs3d7K9jL+95FKr2GUssdXnvnoxovemvmpnonY
T7SbIHIUTvgcGnnIvBPokikIgdF/NFsmKxPgDGBbI3Hsows6YRFSkNvLaS9aDuHPzZeCZGp1rRt9
9Pb+qK+GDDjKxG7R4XQsVA2wdJKNn6TvSGS0mRL7TYy26aKdoNMVDj2YIr0+cM81FpXzMM+UZnB4
4q0npmTGOq8gaOVkixEbK6WvZ0RnrcuyZNux43IdQuSMq9Ok4qaM5jgQ0oX5yPKTIM76gLGMyYwZ
Gd/gdoXnwbzDcCpGdr10UpNvHGYtIcD4VJDXVEw/nW3J2nMx0rSHvtXN9tHcOLsC+XRs1eP7CMJz
HhvgZmRecIq451sKMMttzPF8elU47T5+ZeL5yuI0zFrxRDK5YQvaz2oMc6zBTHOMyRit18y9LQQh
8+Fu5L8lV/6k6V7x4LMu1xG5n5OFMpaAO5SZc6AK/dHyBLQ1MtLoFklUZH97oX7doZNlPKC6gs0c
N3xG/4wh9ZYB/pgS00QlgdWmvnVqP6YeHj11uAyfbDwyOxCiUCFlcR8LQ9ohwdMabdSwr40IjIkU
Yf9Lzt9XBWWwr9x0/SzwlVlD04o/nNLL8JOZk13nm3MnOzXMoeO17GPJQHjWQtgOv2h7scHPNC+A
xyqDvnSgIf4smPUgcd/aNPuXxi3UZ/XWUw==
`pragma protect end_protected

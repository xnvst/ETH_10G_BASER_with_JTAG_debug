// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:22:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
q7cSL2cLz7vCjlL0vZ/1Cwv421+FL7R178o5wi+wsTo84cTMP3lI/KgM2bFflA7Y
DmpUd2vwJMI1lJJLVEM+FavWilK4j1KAKm0o6BPmWQQRkHnSjj4Q1RfSE7PzzkJA
RsazCf2gS+YJu/6JfK59KI/XfOFt9ZAFBpNkf3aD+Kw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16096)
MvtvaEnQMiKD97N5lc6oNd/xasWcUiy/IR9M5u4DoSe+UYr/jZws0CZaK6DRsjPz
vU6f591yGj2YXJdArl4iHMpEfZ0fvspBC2OwH489ZOizKPHNGdKyz/phgIapyHhB
mzaT8nNTgeUFQbHJbL7GLEohZoBSmrf4L9sF4UZ3kNRav668envEcE8HO1Ky4NdZ
QUkf6D4lqPK9rwcTk5BY8AghsslAd8euqlkkHyJxhUsZmQAiPKcp3AUDckBhIy9Z
duyICJiIXo3UyMeLtLQVFvgxy/iB5H2Qrd7m3UHQmFihrVgYKacrZUsxt9aXrGZj
bIxtUH2YWtayyjk15tAPcdtjm7LSLS/EPah7yJb+RhVIvEbWEOnqO4JXfjhV91jB
zyG9ogYYop+vq79t21y1IJQXbsQXszGQLj8ikz2PEnI0wq1wZdfwbd+F8JvxhT7a
d2UKnL3ZfRq9TJs4wUm7DhMf14g5t9TyoDKb8bm8gVmR3+KHZPnZe2eoz2/e/3zl
nxGRRw8OU/zUgtsxZTbzfSYnf+faABwYLv8OfdT7Uyu9GgT29jDsbtj/3Gv+olV3
fYPSbr/QByLFzq82FVmhZ7SvGjTSm49gtPYTQ/or+A4kJvysFvObNpfOEbeCKZdb
M16evWUMQhNeQzpcofJiqqKAzztZPuQPkrDmEQeUehAprlaWktfI2oxz4s8NypME
Optkl8hagexZBi/g/4sdacgZq0g1xy1VdcZ/5S/oU3slWg3lbbS2gehdhOX3cqCu
PeAhAPbIAHmKQAY/yYQ1YxZ8rLsVsLTlBNwG0+stn5OTlyWr4sGX9vjb/LEDjh6g
WDdQ4EcNL/YxoY7pZGdZWJ61XZrwgoTqAO3IE+LQfoHVmD8WoQdDVaiaOCuN6RVH
PLrGEQMx+R3h17IQrEs+npDGhDY9exNTP0tqIUPLu21Ix/hIl5Iqaiiz5jXP0YdV
H4yAEfRrWAlxdlvDLDDNsgmi5IZjR2yYis1ClSvvIcOyTCTvkrcXXMXajsP/Y41+
AMpFYixNR5+qng/fvbrLmm+KBXBqKT8bzPy1Y93NfPYbul/bWdGYBGBKTLxqC9rz
uUptojZlo/9chNLQ1AC0vo/R4oT3cVoe4YHTS3yHeZ1za/PUIOapi3Dlgf/F3SpT
bBeFG21e+5wM0dsbPQiFnGgXJDUGS4ZHMV9CotrxYZgg269bkbY1m9wpJqouPnpu
+pNfOeHTyiphNkdecLmgcFc8SCkTdVcbDtcGEiJLN3Ls4unxNIh1PivwyQABO7uw
wFkDsFo+ngXSs25QxG9pFBxweWc0BkTKS4tBTX9lFTKWdbKcm16LY+KKIphlfnGJ
Ejf8V9lie1ssIvFFhaOcIz9Mce0B7rkGmwjSkHLfyNd1OjXiCpvhUb4jKIY/3TTW
1VcP+qMUmdbkQ6Wa7SSzR2O1kbMpxB5qw9vbO+yop/razmYVY/8iK7IO1sEaJZLv
U1elJKds2F1fP7zrvH8h1GmmDop8nJpaRkx5c2LWDnI1X0NfllX9yNuNltmn1c+C
3/7mkt3nfTYrDAzfGs5KZE0nPv6xLGnUe6D1Pt63LTZ/IE36D0bMEMC42o3baxvp
rIVE9tcoB3Wi+jsFOZaN8S4D5gOZvKkvDmMZV3/OvKUqvhloBnCEsd6Dilyj9mtG
fJpMiP4cvrYvTuivdqZq9KF/JGj/DSN6c2kS+mgheNp5rHthLwxwt7bWsvU6HoBL
lkTjY0aZ9zQ9IuxnZ3TXneycsOnvLYbZKIYF82MhGv6+XjXNz0bP4MB/EUF0Y4uJ
2x9Kcz0cm7D7MCqhq91eOzDztiX42GlUhoAP2rA7VDcJ9Hcm3Z/ozk6qCJqKrNyx
tyhOAYd7Jnz0ZUMQbdeXwbfKaVc/T+y16x5TvLdA7O9QUvArZ2H1ICAd+Z+q5IUc
Nm724VpNshvq1RnijlA3lmmG4YgBk3nYYeaR5cIawFcoyKnGe1dySY3tzLQFwUZL
Lk6qlp/J4VuBHnfk0X3feDJsCGod4eo3MuchixckONAcx6ebn46O4bxDO0Or6Ak/
gnaYJzD81vwpNwGwNRdjzw75wRUguF4uQnytav8p6PCE1nWyb032NMGHoCJ/7Y0E
18LvQqsY9ZIKn7duFLR/rbDnoUUt5TDWFo4h7bNBKdmjBEuCvLVdSLyN/fUTjXv5
dL4S8MBocOyeYBR6fUrkp10IQXitHhxyakizPsEJnjqdqSQwzAA2/ER8+yqZ6kyo
kR+rwTjHh3WSiAdX6924v+02X/GvMVnpRQODdcZ23ed4czqhdgtJWOYC4kpTOltl
LdLOujeprj9yD19XXLvcC0ufxlmR8ilUYaGaxZbD51/q0pGcV8iodX71Y+IXAgMr
+Cn/Pq4lhe9aLr1kNgjUrhGnI8wL2IlTH0LLNYIxwGnZeRplY3HdsVReK+CTM+7b
LVbNHT+QsoMmRkd1WeW0iMQyO1AHp5hluPTNL552GYIQuPIReGVbNVt8s+MLT/cs
9FFG+3GFrnHbe4G+j43p4L9EPwrLjJP62mAR8ALIIQ3cL0LyUka46ZOFhrzeD4/u
I/Xq8LhlT+gOMrPu3vZcMZviQD0iJ03f5EkIMYXZ/y9wmgNc5rHDHEIktT1szRFJ
UeRmBJbaZUNy6rNnGtHckZ8qB8X1WTVrNRr3ObRvgKmX19NAciaUYn4vje7clUff
X8IoJNFfzhKqh6MjeRIfm3RKpuC3Jm8RvYtgb31h2qY9+/pwqA3ouB+O43wHcU7J
kSCwuqxbQM3mTyyeXwaj8ZWJd7y0F3gI9hRJ4qON22vtXf/8K3Zt6gsYSr8Dq1tp
UdYZpXU9wlj5GLACzz322BR3hKoipa+XOKyOQJdK5VObpDZLo7mLK/1KcI4B8W3g
qUqxJmFdwffY5RAWW6Z7b06uB6a+8oYEQxwKhD70ws9Z0AeGpqwdnrv06hrVzixS
QTmx6mDsaIkv8y5/P8vGR62fBJjxpKaOOXWlZvlAx/+oAu3YBAVLMXpUKz/7lNBZ
6zOiPzYlAqjqrGsQe1J3QKK03b+TIS8Z0tcaqG0Ey87Mgcg4neXFGYFWyy1qCpQE
5Rlu+l7CMD8oJN3AWEb203L3oiuMZgxHuEyleK81YKflyl193koIYXyUjDegUO5z
KvhrW/oD3CDkkMZNzEeabsZ3quZ3q4B6NcSLm0A/krui2uetkpPVi2QJs6JPY++Z
+RCS53IjU6cGNklvM/7ruN3ZYpMLTNDhZV0lD2dvQRzCsqS+TD0DpMlgPc5pbQRo
odJLvBDqDGNYQ2NQkV0xGb/KlD7tG+TlV20yE2n0InXpnicLp5/ghKJjWgnHXFaX
R4+BCDDxZ1ccT54RzP2tI7F+3CNBomxtAmoMzqV2vaX1isF7T8c1nyhQuzxmb9RM
+e+xrtaP6XZsFrxXamkb5TeMVU2Vcc44O0+L2O15PU026NRQGIsl8fbkFknQZYUx
CFsO5sMatRHNC9gJwBMTjIL128WljH4FaMIgB/BxFvkVrlUK8cAx77j4yHecrUxF
BTjR5eYp3y+dKqdGCkWpzmgqWERf3sgFeENH80Tdtccb2aYd2pGY+Up5PsOfPvtK
W1W0MrT0m2VdG6JC3SkxIhM1T8uZJY2jUPub4dui2NLOn7CJjxbJlf8cKiBZndvF
RmPuPJYGq+XqOt/ipenStO6s6OCyCZtcrHUfv3C7sD3ZZDFEATyxFXoHPY3B4wH9
1tOmyDklzQWxcDYThhC12zTO8A0vsk3mJZBHumwAp9jmUc8EnZ4XG5bPy7NIIa/y
XMu/F3H/+nD+PyZgJc7il4CpxmmizWA+txzPR3kTIWMOwmMVov1v3GakGHLKpHNW
NVuykMbRdQerFu0eAMrBKm75RXOZ1pWuO4UG03iGEvSUZZP8GL96jtcz5tRbHeOI
JHdRSjGDGCM8AyuEnrHnjFdqvSpbwuHOEt1j2IIJWBGiGSWoEiwCBkpT7yx9BVFw
g99zuKogoqPjwPeichPVhWifWwuxYwhx2l++m1q+NPCBLrxjKeBGXuWye7Y9pacm
B1rRG7sW+u+I7LOQYwj0vaLu7mOe3bgG7787Fl27Wz5Ype/s8Lu+w4IcXfsYKjix
Idgh1CrGkWP2+5fHf6/hoWMH0QK6GEcR7RZA2YiKT+U9i1twkTCPxBCkqMD3Xbge
j+4S5RiXMLf5YefsYsyRk8IuyB8+mxQx75N7W+7ZwaiN7ZtferiM8orLFnn7Qjig
Tb5cHNXaZ83SwtFoWtknJhqcwkBjweFkODK3hhVZU3yfBjVxsbGOJR4MKy2WP7Bt
D9321zhQOt5sVgqXSNJxJmZZXwIduJZLzND6pOU/GHvg8vMsGn3fCN7keHO5k6l6
2C8hSWh0b6ldMl6mEoCd4e/92mCjfi+UELssogyrIQ9/hvhl0ZhW69sQBUG+wT6Y
/PU2nz9oiAbe0ltElQ+EBOuUUXc1ozOrpLEhnC6ZfJNqV0iKkypiMGDQ+m0d+n8g
SiApF5JiNCy8IB/7y0GAMH0ONYLA2BVBynEePfQnoPlrONNchB6hOyRRwa9WR+Vx
0Mnu13LtkL9qsgQ1NX1OSTf/sB+JKujqCrxhE+OjHogd8O8SFl6CE3X5UgbhoKdi
qoVja5AV9j1UqbIgVATGJtKPJ6V7Q/9irp3XqXG4fr8RzXUMTdK7OuBEKMlPP43T
Gs8aWKVDcjbcSc/lanXBT0WzOnd9Tmu/Q0G0acaC0bCB7K/BYK3AoQ5dPAZpI5hu
tiRjMagAAxJB+3bFExbI8y3QjAEtHq492Vhe9NlxqUZhInOG+blX4gU4kHJKmPmQ
YXE1d71569N5ug9kYEf0qj0CDJtk21glQ/WaaGM2GVN8sGw6BbnPdPJQ3wwlJG0n
FIqXH7ce/8sZ7UOxjpKGDHsnrY4pDDtv6YWKnD8BauIUFjf2swy2rSIkwixTrW8h
t7lZG4MijTHMz60COhPp8LACc3OukFfjEYlnvw9jcXfT4B7TYPNtwHN0bS7yVX4L
M/lfBuj8jeV+ZqMrBOJl/p+WkVQbTVipuRqc+tcY0F9mm1buI0CMSe4u86CjWjro
tUi0/GI+GY0RBz6Djj/psWBVhg1HVuczSCD/TBGyZ079rBHBqnvY8T39i558V2y7
aq91wgQ/87bZymLsxxrtV2kqXxa/qNmX7f31Ci21O90sQYOlaUKDyaGiIe3i6Xcr
TRsu09AYwOJgmgS18JWZxJBaqLkgFK6NsY4DFAnySr4m6t3IUqAX4FBMOUEzdoU3
U2T3ud2os9A/EL0YlizhSjgY9mXb9ha4xJs5p7bcT7vmw/Sf5AZes6ZeDixxIUPx
xeqlqAkWhfHoNuoek47HLU2s5xzOKr1aiOfDXlqDQ1YxFXm1QXLlCpZmdjbz+lH6
FhQ9OXUgh9vJ/Lj1oBdM/qjnWVq8IQQnsX0CAWlTnOxUF32/oAQYWveZvq87SkBN
wQaCbn0uwlxJ5ZVj+d0gx/CRSwvwjKDh6405ctR6Y0Nig7W9LF4gzqEvUS8vLiXD
QSQZPDpbdjUVGEsQSpsAD5qELig1YYq03D78mGL1WjWgQ4fn+qhpLio6x6nyHC/g
dk/woLdO9W52ovYp5vRIELqWWbhFnZxmczxNRNfzV4+Hl+YLUjK7jwJ2wIbBUxno
/7ndXGwU2jb/2JI6vI/ETTxwJ7cUCGERriEltsdAZGR0/rwf9jzUuoRLqffyhsab
euGrx2UPZBIyNbPKGolweYCsPKjUQzdKpkr3FA7wkNvCxYgNLmbha3e5381+6VyN
Np0Bj/F8mW6vEOyLuUjmlihvZwCAXtaLMAmdeOPZR7AwqfQaIx7NOZp3BTZAUWTf
iaax6zvKs4voA+ooh9vCyNiuIb+hKadqy9kOrlQQFc1Ut3i+s1qjMVJXzi4hwt+u
WisNzk0m/JbvpC2npTwDHwXyIiLcHIzjp+KnpkcRgZSvmA7XFeECn6vOOtwx3ftt
SUuLZLiaGfY2Nz+sLkYn1TRfUywpO1d/aqJ9zz8tjw6T3DUSbVhH/6Xh+EWwTjMk
26xJorZJTtPBg/odCxxgNt4LIsfYhVVkgcMMh3TCaIAfu5Cn3pOxpGJqz9JwpJST
P5S+K3q7qBfS1mMczx9/0/8pzr0g7jBkuopz9O3Q2gEwMURcstGBZcaz/7eWHoss
SVCjbf+Ps42HptXYiO04yteSXwo0EI2LAbHbnf8R6AbES5kGE+TPW09870iBVI30
rdo6zAZIfh87zR60gf6mtBvHa9Fmnn9strSs4sNbPXzzfmnjTJN2D66MKcNMhXeU
hR/NCkBcOQVQcDCL4YCt72iKTskqUSAN/MpJdSa0C1si8Qrm5B0mJeTnKoEzq9ne
HG2i/NAmm1pGq24jb5sFWwneuisCyBLiChM8TvQE11AU22h7ow1sATeSUALByNrn
6GXtgQw8bLM0Ckbb975L+L2B8Y274Bobs2aLrJ9xOp6CYq3j7v4KsMKVi7oULCFd
5uwJDYV0+HZoVVuAL/x4cqEkYr05P0yXqWZrJyJ8YRPXbkACH7318/niX0cqc54p
c56DsvAQuwr3TKM4sWJBJ4VH/XXMHnpvTLVrM5brmyG7DekSSDxIPnbETfgbfx02
kxI2K31wZ9DN1o7SdwcSBrAkMpZJBEh6MKont1sfITuW1RrDPG7mzRJwFr+tmPYC
USCXwVuCe6ZzVhT4RleSbW+RaApGHt+MYpmhmaDWDv0fMKPDopaMM5IJfvux6WfY
liiVgr7XleWkp78gZKlncH6xuA0WjfQIq6FAHeW7riixRahmUB1K5CBG5QPsq3x3
Psyz3LfS+ccaXhHG9vSeqYS+1CyR5RO8eNLdIWYQwqV8ICE9kI7S4iT2S1Ii0hQm
L+56oDTnQzvbtBgSk5cZ+xJGehzTrvpDkD2Lv8pCLZMRL6XBb42C+uXzRmRqNGRI
++pSYIs36LGW21z5ZBT+XXnG9Va0dAyoWxEXVDPDP0DdJhbjoFjVe5TtElqCFiFC
9ykhyaLN3XNUgVlrxdG0SV5+MPm7U5TXLNx0wHPiS34lC59ForKRmD3nKpc8K7DR
9RWeI1kSpOIfKfVnbd9tJFghyAJ6gZpd8iglaqxFo870n4wiTS88BRZ4FpPZyGJT
/7kyhieTFDr116P5v1xT4FG6cJKMWEcDvIRENG1DmVNgL8ugw5zr1q3QMNGvut8B
XAuNJblEiYPcrYBvr+g3dkiu/AhhxRlYqSJNDGrpLhWAdvbKZLrz+r2tj1JO1tPD
xPUbJSlNEG7JT66yxy0vCFWzPSDdQp2JGLM8bHJlxV8Ye+fI5BwHVjtGRM+iVyrN
GUF1Ef49t8t2atgbcDMOcsUaBHFBA8IFy23RIoCn9TK8Z+190jakVvDy1pNjTPla
fOgvvCSgYCSml+9/Wwni4k6AS/YaHALBh6gGGdc+D9Sf3RjAQYvzD7dqytr5wNmq
V24hkyxaJK5a5qailrITflQkIiBaiFn//yh8rNQsGJWBBNqv0x1fTyvMoLEb9Fjl
Te7wK6IgExemasZ8AxQZgICOQquSGmAwRvmE+RVj1F8WYjFKPZxu3/Gdggdbrbka
G7MGefNH+exfbibsTYgqvGSdpI4fLKlq3b8B+OvTHRh+JnKd7Y7r59vTVr4BUlbQ
wHn9Oyco8u7EjSBdfaFdZSDvRoPg9Qw8S25V22FewaNuZo/kCPWrMdQmiLpZBJC0
HJIU3K7xUeofcV023MECAHrm48STcqmLuUB95OO15u+RPBvCILhQv7+QFFevQPU3
OiY/COMBnZY5jFrHQhLzEhTjBonlF8IXYr6CsDVW4kYOQAapyH93BIkKQdTIr3Mr
tPq/xL6J9p/i3sxojdfcaD/AM1XLhV+1sV+ZbPYhfPeub1ZM37GSkXcft3uRQaLq
oLXcGrt6RKDD54OTvSbYWF+b/K2SGNwpdCqfBheZd9fvhjXas7INLaCKNlbg5l3G
xxgd8xfFxaB98bVaYRvguv+E0M1K99eisgaOswNkXzfS8BlxpxPr4Rplut60mUOh
FTOz19cZnfmlQT8ZUqrZe6PVL7AQZAOb+8k/1ojSCHLxbHL/aFDtf8YL1d8R6QwM
koXFX8OeJjXeO1c6pLemkk4H+1ni30hvWHCoRrjDIMuaHUoNNDxMIFS7yeCKrOUN
HMbuXqm4BHdKzSH9bCecMX76D4ooXINVfQj+Z105Ujoy21mvJtyutjVlDjq1BDXD
yUGPHShh1qc0EsPpffQ4ojylc1gCWLdAsV+EjQoRU2rQuCUh52hSvL61avfXyLnV
IOF1nyOH8zFtPLjs7siwb6Vk8q9AjNXLqY0lK7shANicWjQaHmdJKc35SEtIzPSG
9fy+FjnjyYfrn5RysH7JrRJnbecz6vX5sxklaEOKvd/rs0IAA2rGjP4DKypzJVTg
QXREGnrh86UuxO68L+tHd9Z6vvA/1QctdY/kTVyiKxWa688Gt5P7wgmoqF1uKEsZ
Bi4IJ+GYn8gsWIJ1wZxbs9i4Y/UMOeoK/v5N1Wg9NByijzznsZ6v6XdcJgWR/hz9
psYWE74UOxkaZGdoVe0gWwv9x3oUi5hoXh8WlklBKjH7gK4VfqGnJgwROHj4hq4C
aZwwGmhZulxHr19fBSHgKsM6WRcfgvL2IabM8uZ+BCNhrkfQEf2YzyjzXXdQOf/u
88yhZjIdoTQkQhPB8hb+cqNK5GDo021oby5fbDfb1CCWhq4dwsOE9TL+WQ6zTEcS
RaU1tYcvEQHX3UODphLwZsBQdSjqmWXfHUB4TWZa9HFeiX1DWWqA5iJyLCYOzbA+
vmxShqkDjf5pvi183VBNg4NH5WAO+nELXgRhxToUWHvf/L8cn6SqI5CGfxb2i7Wy
Pfni9jyivqOe4HzV/Gb0mNrgycWdogN+No7QC8DNtrb37sp0ie2p4mtU+guvoMnJ
JyJ8iJUyOAOM8YbTzwTu5PYWqpiZya07pDB4pP9b24VZTBKcmrKBndDFXva6cgrZ
mz4CpYSncBH7yEjRAsjwDwXjrY9XTX3WHwJTTdWrBH2BGTedEF5s7JfRbWcQGzUs
kAyGsoaat9ZyRjEv+kzF9pRJUv4xCgdxdjeObBemO+jKl1J/2CGorP0eSENerApG
LKBtgmTjVaVUa0MAQKiYejYusXe1/8ICqwSGBVbAvTUr5gdiIOO82bQYs99BmANv
YjMqXZXix9yaojtyj1IV/lIJ4/yAFwDUkr68/0CEdrQBdTGuDkxuzBcn5O+AhnVC
C+qlE5joNsa5ZXKWjWA1aS1esURIm4Di8hcTuV2/TGnjbqgvRKLoPW/Ubyvnja0V
DdTnICsmaM+/bWmWtwrjDBVoICxvu6djVqNE2wnTnENU3gxbmPeKRuR7ZbkNjjie
Xj0af6lO8D4zaftYPHnwVrk/A0IvJ6Mcvi6paPABhXgR2OG9X7fxYQ+gjpJ5HAtL
i2fpjIvHh9E0I+Uu42h+xD4cVogduzPjHcJdHLgxcepI1TETC0NndBHDWegbJ0QZ
YtWNxeHgM50q4HlHo3M96o7NI+afWDv8baqCz82OuJ3ppDn5GnyEn8Knj84ngoVL
1uIVh2P8Dnh9MSfoFDZQoHSjqLMXfoaw4Q+7fyvL/9T03HXdKNj9UeP5yA8clV5N
XqwRU1C1x15CtS4gcSiB5jG30uExU5L7vqB79F6yVrBt5o/Tf5y9USdDqKMpbMwu
I/mIw4WhyNVR2hDLKBF5bETybmmfn/mzD0FnWFT0+FfRoopRw00hFyVFa7TCuM5D
KMTUPoytFFjgIjWLO2atVY+e/hicwfxJpljQda9sUjOWMAMm/SnLdwqwuPpPTi66
xWjrje3vGlY8AGHqg96ElIkf/i1HUUUAtOF9yTBKlIQX7W67ZHCc6dxYlpVbrS6u
zG2GCdvRK4coJ1j0T2tW47lcDHpzxFCmM2vGshzpqk0RXIV+oz/kvVJzL4EOAZUD
5WHw0lHLYT/zurRdnj7MeGVvv7Hf2apMoFHh7yrUlObaxhnrO9x4QGtdpHn/w6IK
qg3kOPhR7GZlYX6zcA7Fg/YrgUeFJm51/beNeNXwL+iUXnNVbqiDC2xuCp0FbyQ1
/B+WPMtFMP3qDT6a87ORXEWsmcaLu/2MFL590DWviEYgG8nSZVlBhQfCkcAiuBMZ
AeTTKe4VM1GE5pepmZkN8juM0cOjxvOusxs1LWZavsxldAZG1j6fHElnrfcCA4Ze
fz6lkE6S/12wftf5rWcDJwR4FMSFYaJ0jx3EqiRnG3snR4rxMeLJslFhfKXr0DpP
jy3PbzroAcpLGVijD1ccMBFSqHRE4nh/P9xgE7gvK11mOh8dQ9RMfsmyXUdqwibk
ffOwgDqG17scXxD2gQ1MPQ2AlDN37M+oT9v+RuOQWhcnzgbrfKfI5p9HfWkcRFiI
+JRqbjdYn4N5XQnUPOAayBRfct1EYqbpyJwaGnr+Xg/nI8AgWfW4UaKA+b/052Qb
UDZFRDFNf38hqt1BLwWCeCfOCeG2Q7ajzA1o0dPwS1dRqTT71ljPGaF8bST49wrK
O748SmowWw06VCuMCf+yQQpr0ckqlIcJmWuJL5LNa2a6lNJeusHhLBnaYVVy/qK/
k+YD0TBXHk5/V+vNlZrxxpg3SMLjEE//gjDdUwmdU08SlQC5h+KCr09QKkfPy+AY
ieANnJsWVULTja5HjHu/ycmy452iXwhdCknTY78SV+bIE64futL5rtGRn0FkjUz7
EUVCuVJn3xDZ7N7vmDd5lPnl3/+Go3L60l3FsLTrFRAhTzOOeYzAfQjC58Gub6us
BCqg1ZoNnpJdQPXrkGJVN2y3M2MaM4Bc7JJj7lCrVlLPqi6jDDAvf1VSPh5LFG64
OhLHzDUyxhH6w28rVYww/P22iOMjo5uNA734ZaE1XAtBwGTox/yqbUYQD4uP2Tpm
e/SuQ4POKwUip7eXPQW7th/Q+Mmg5cmKHoyfiFz0EQi6RJGaCMCLGppe6W+7aPqy
/QRBoQjz6pUQLdGjXgW4jOTqVKJUhz6OG5kFA9y2grbSw+zLaYXEamRtPpNml4Jb
rHoQA9cd0uCcF0a6N7W9Xh9eUfi7A90EyhtIqiriMrNf88GmEwpE13br0TJdFQ7j
if+/ofMPcft7kVG95d+rhngR64coZ7djT/k2HvuBBfJ0Yj3imoUxFuhQx2kuCRrc
Au/BM0QbOTvV/KtYU51UJVfKf//T3DAXGr4QINOkmyJOf995OMRjKIe1AclmNtuD
bNKUYU/w1gd4DTOQNnpHS2FKg0TVtAme4h9cHnnPah/rKVIQuBenlg0fd7L88VkS
wRsYhjomvIGcLhe8Is9BZu7T+f66YwBDR1501R3McNPrZYdpRaRUBYPoU5M4xfTo
bTNijZokJEspKT1TK+Rs1g4v1TeGW+/0vzwZfpg6dTBIFj+q7vPOvZ3zJ4QbvdkO
KQ/N3I/fjvOuwhzcwBqDx16vVbLpnsovtEn7x82tBK1Fjxgvzc9kMvKB543f1JtG
DSVkq5VMbWc+TEpvxnUt3veNUaEsKCd9wm1sVscdeqedF3nhV77nnOIWvY8TZocu
twQrm/IN89Pe/sFlHMqEDZlb5Mtlf/jCBCE7RegxeyPdGIRO3MIV2i7pxChruEh2
o4LrYtBWV67fzA0bcHlbqpb3qofihYAgIKJo4wKdPppThK8Jy46ANxB2SKvPkjS0
RjTsJyGrBFxDNuNjg+uaiXwQPKe1/YAmFUmjX776ujIZgPJkLzZ+iCac1bRt9bLp
I4/mxPaU/8/T90m412Wt/F6dI55NS9hTU1C5fIMV7QTtzJIHwmrPI9heiiZZm14E
W46c/+QDkyg0NcFVi1mK6eA0Jba47LUGkXpVM1BAgC8uG4VjU2//GODmGQvzOcLT
xYCQFiViwJSaITGHBIEVTIZctL2A0wl7bFmdo4x17GMd0X5aLoSEIFLtrYZfQzpg
um52dNrBGLhc64zjBb3X24PJsMeFjTmkM8OPV1N4kvbtF7nUMnABahkHi0OWfppk
piRgRylFM5emlVeLUQ9wWkUXH6euyTU7ZfEY9J6pEocSk6BBGzg2QakDqvC5Q21b
RWgQgdO9qniOWthqQB+aqPEb2u9PNfBkVcnwVWjQi+TMtc+JK0jjHqitcIlO2KPR
iNsfm3ekFLWDaLujfNhDHed4hfDmteRIS4LQchADrx7h1UUQvbmA8EASS/E1uW0A
IW5sqjL1Dtn2G4WPEbOOOBmoIsn44DzgY2RaGSvXk17dAW6qVpr5QoclRga276Ey
gM1wDdkYCnqKVY9PbmLIba5uYlAVJOtf4qrHNHXLxxZ5EGoy6YxNPczsyi/uDxs4
pRYq0+l2Y2oUdLiB8dEzEdm9uVKnNvGgy16Vxna+F8qeoZbpoPK8Zy3L4B4LjFeg
rZdGkR1BvXzLQ8hbPx/YMcEJ38CEYzbVKSlQJkuiGSyszwYZWKK/A8jhK+sc8+HC
iUD3Pkfi94U+xCDtx20BywnZDn8umcK8wXmZy+PTSXjWubhiHxrR+FN3UYtO5+yp
KQ08d2VNVnNRnKp6wDBpJinwAD/yD62aVb8NGI+dH4wsByACZEjyLPZp0sCuZbIf
nXrd1D7PyYeO6WItIWxV1rVKicNG3xTP9WAw2HvHprw3EY6Q+Kjq5vt4ztJhF5Fd
8IDAII5AmadKwxFP6kzJqfHzj2mKnLfMsTC6glbR237DHGzu23dgomeY4uskclGL
VU+Oz+n5RGmefOpte788Bg3uYiUcSP6yeb+LFZUN4CzaXbdrtqlIj7fOO7rSh7gX
KNRl0aMTOqVdCcirX7PuQnbmPxQ3XsfNMn1p/yRpT4kZfn8z1T6IqAVfEfIw5zJ6
TV7X1WNTs/mFaS2rmoKrozIVBM9CiW8sZ2NqMQc8gGBqdeUcA0U2G0tLRCazYK9u
hZXVN0as1KOWYd4scHV5CGLvTNBsZa1zMpGfsKbWGbucRFD/FQBmDC/OyXJR0N5W
ga1fIHWWRAAPcKXv4W2LUB2dRrgNgKsMnkP4z08gcmugx60zmfqEu9IvIlsBXb0g
JA5BXGbIZkdMmsxGosqTdJ9zxSTMrPGfRTlsET1O1w0oJYno03QBnPAJh4PMP7Tj
qS8o82lC3yAEjSdye76Svz9ppoW71lSfOQC+CyFprphTnX8XujM8AFseujxd7UuI
dOBZgg6xIIi5cXI7WhzkzzE65u4RrBxczIZe08mbRNDFYiTQpZyWrvID/0jhdrZ4
JHsQ3vjpsPzHkAURH5aUGNFZvACKe6znL3kjgJCDDXFtjjFNTnkV+WTMVtiqPuoo
NS1+/O/G1xYkVTaW5UdWiTRhX0FD0xnZ4JCeWfpZohbjLQ4Y8fHF5q6vmpbtbHNs
U+/1mWH6KBdhQwLj9ExGx56B+Y5IlypfBMyZv5CK0JpHQPIwQrk42AQJcmsoqe9P
vny4w1eAnsbkQlAkWvM5gvdfW7YiWM1sLVF2g0u4e8POfB+yOhn0vcLSxzISBNH+
Z6I6tAUO6fA9qNeQdiL4Y5batl+PEDFoGkd0/8pM6XWHjyhCLGTMPk2/DqTqIc7q
DdW5o9kJD8GNmHh3dzoWrZXuOcQKxltWkC5Jhf4E36FMtY8Y/BLFwGkliU3X8m5r
wP/l5zweThTLniOH8jchjp5bQZGEl4qnMA5ydlpLj8kYlNCFbKYk/zV/TQMeWw3v
izFONv0OXd18VGyv/G+gsqTmpBOi49O6IfNXyZydSE39wMzg/3+9xnY5QX4/bxWk
hBr9TLu/bH0GXx5u3w5DPNdtfiRphciHwUboAemBIvh26/jz70q6DBHEpg4h1pGW
nqB8FhGq6myYuE4WapFn846CaqwIW5VFaIprbl6lAzAA0Xw2lMKWGHKN9sBcZ8XW
DoYOoI7hL+7h26Ppf88HsEKp4YgWhyK5elFk+xh7k+31kShZRMU0vFk+g9jEo70M
VnT9hCACLqRUtmQB5XwptDrn2yqFFVwyK1JVO0il3IojHiNXb6jUa883sGaDy0nD
C/PAB86zTusxIPYcFsbKOj05+BtbetrdJRLIad7FWnq7GaJjMCopr9coV5qrHo00
Z7XZaQ9Fd7FOIOFZhJ0+NTuilPha5UKI6Klqb6gWmRcWZd2Fb3LANX93SJU+alSH
PK6LiSGq04xNXhgSkH/7akJDei2s7k0G+hYRCMim6vNSvF02vk5KxMDK5nH977J9
osAmFjxwnKloRbTC5ak0/m1RgL4NwWDaFP+8X5pjoL2nIGUIvlXGsd7BNQFUI0/9
Jew8Dxaz487+F0hlpilr3NS1oL4Bo0Q7SwbFGUpTEOweslKGary+63PNZSS6TRXa
GQhUMAhvVM698hBql/MgJUSLsStJIWSGq15I7F2hZlo4br/rNujlFKbS9EvIeQcV
lYil3URhjyrI4kS13IrXr7Ha6iAAWuAijNu+3VmDxvWW+yuKy0+RE5bgv7a7KSht
DGIToVvv8NnDsoy9TkF/0Z5CfWgYcN3lAtcMoPjtgDYDHZoaSsbyQAtBji4190z3
rQe9a3TE/rc20SeUgHkIoVGXfgNAjaS+1gfmLhHQr0E/36Xxv1ayKDGqxG8OYhy6
NAm8KRJVBuoSBedypenaX0qW/4KcADRnkJU9LdSAVB7ssrIBBhUG00sAxzbTLKZq
kk2dgOHoc+H0/JFY60+c9ZI7QHDsvFe4jovuyTvVOoYLP0q0kcxe2SlZrYCQtQJs
rXuPvsbEwTwxH+2oU1ZzRu9IxZ+5mowWZ+DELRYHNRs/xbY15dYW/aWZp21AepqN
c56JuM/lHbWvJtD4FtAuVxyQa9KQj0FkkyJU1XRjuqKhpldJ4GCsbMfGJTfRbBmL
G72Oukyj6ZiVCZzZ4ut5c7lEtV+0jKMZ+CwYpJj8Q6Pf/O3WLFpqviH+qkmUCvQV
8JuOffeAz3Pi4fq8wi9fKrcoY0uMGmAa/ylKOrVNKNo/lcZ4Y9SahcYO7wv6cf/b
plXKRI810n8AZlvBZf+r8TYnuDWno/fgrGueIBOYN1WWOEKk2lOlUnssRfQrpXMt
B3JeJhu9yAg/Vq8vOA2aNBi5lM4uruFP0joT3F2xgvKQGUcV7ZVLfZQcFmikfk1B
aCXnKv0rZMSgaTb3nd2S2H5Yyar7ALzdax5/mPEdy+Fpqp8fkjMbdC3SALEMnSYb
6ZyDEUV5to+vP0RrO2BBeBbXbiJ/PXmwZKCyn4d7NybDdChlHOexvctPIoWfOM5E
BQNw7rgvlM3dAYRMsjBWepWU+DLhn1YbJzuvPTudv6ecA7U7FujrXnbByIRpPUWL
vL8+rXN9uAGSR5rP4MrHEEZXe5PUrY3HaBmqCvUytzCgjhB/0fKKU9AZUCziqsZy
EugLnrpX0LdncKAp7NaOfQiiHBYIq4CRwbl7MOftUuEotS+IjmynrzKMjemsl3TI
nKTJ16OnPs0ivk51M5PgId8mpy2iI6YjSYe55YU3SxfU/9FEp/IHcFa4wsOtFK+N
EjcuH8sy0YTrl4psqcqbVphmjiSeemyS41CZydsXJ7I3Stc54JLpRF+EMnrT0iQ2
VNHKH8uXdllBu41fWzXaYiEc7Q/43HUSaHNEbpCT6s2TOlONT498HYvNhxVyd13R
czdaPJ3MBIGNEmfmSB7Zx6uXbuK9SpzOuClg1AZo48v8wTdB9dZstAIuRrFyPBgm
s7gFu8aVVQKFHP8BDktWmnzHBOtpF+RYuaJKyuQ9zVvzQY2Mm0BEAhzXTf+lruqf
+ZqBNdsDaeZLyOEwmn7buM6h9XjSEKsIP9sYHh8oX7jftU7yQ62UsKsIaPCIpZah
fv6O95d1k8gR/AhrGENqdt2K3CByt1K1nSWI2bjo5ibbYo/x7V52KasoPrb6gzjw
B/+SUHJScIzlfIOaq8TkB0QhVLk6gpbkOS0T6VzsYq7uUSoIV53G/GeBjzRweS5C
Gw8ezaUvhOryvSav2AAGSXUOGGH4lXkglIWkvZdl8khANc6kYqF+x3MlmhTT8ZtK
kOERPCpz9nQi9qu0cMNf7Vg/yLpt6JVHAn2a2ldoglkCFyo4Jyjeo6Pc+kI4Dtn9
Hm+uLFemKxL8yByrFsWtnhJKftmMD9wJT/ONiSYz+hL/PV6aLDGjJutZddUlIRhL
xjeuuwJAxEO4Lyj27ydtXx6GmhYRff3b0s2I6o/mnJxXv8b4H950keV7mpr8aoZT
SbHGMa2RJg8byIGQgOCWa8tl74mQ/FqUUIwZJ5f8HYdmjfTySKUcvFjiE8DptzMU
vqUY9MM4sl/IzlJzz41tKBLLZ10m/8tq4KDkvIOtZ9cwJWVaNCdiNCxy0pWwlSEu
JbgzBkiRPX4CJxb3Quv6g8MCekzpQQt8se8y0d5roEmTrjMdnr9lJrJp3PxTfZak
W33Jdm/m1Nyf61pER3WVp9XGnqdyzaekzjw7Cx0wyJo/rWF5cMYP/nFQGadSScMF
Svr6cjWyFf0jK5UrCArYqIdIMD8P+d09i0sjEQNYmHylYKas1cKCkkAJEywsIojB
3tP1rNhhCbRE2OKt9HAzTAqcunmJwgaj8XhT01DUHgh/YPmzsYoAC4lbZE5u7YmQ
GsyljK8okp87lqpxJeeuGc4jDd+RKfnjChRjt7mxhen1EfYl6oL5ZLSdM4q6MiZp
FYWTUQLkumSCk3mgQSb4DErLb1vTe92e7zKSJocRf3wUEscRVS9mas5mcqNd5PPb
O87pvKXNY8wxL6eCGEY6O18uijUmFbkFSSU6enpLR++Bgf1nqMekBLoaniuh78+S
ngczgRSY+Z8CxSUzadbVSpb/rSFmJHvi5M+O94maaz1FIlhDK0Jh4htrq8NoP/I7
iizKnKlS8EYVrPhv2tbrHMQ1dihemDtE+WqvaNu41zKGqIOYg5c3YBVoYB760Opo
KgUnxdJO84pc097U3tpdKb0KIVEvs4KgiDwBd/9JiR1v+wxHjAKtQMufz9rreCpk
MBysth5ZQqBkDuAY4Wq+g9wEaOFFAKC2mFKWvJymi1SN4zSGR7+l53UjCSl4PjYL
aQr3RF1uoesUfyMhjGImsdVeJJJJGCI9LgaYlQN1R+aAajr6NcH5wkI+bAt9131c
evNgFIPzec8dJUU9+aPckPB/NYcaONvyURDlGBP2SIWnV+C5zJDNo2Y1ARYHsGEn
zjWAwSA/AErKoxh+kCusAupxGYmruCFV2340Vn8+b+J+Vb6NUZz2At4u826rNxuU
/iRa8aMkkivotBAfophJuWfBHIYbhiLD00bC5WH+toQGDMbSdih8HkEGWxqDaCHS
lPZu96GouGNwUtpATplPm6AxY1k0WbJCqq4FQpBoZwEzfoNEaDoAhSTAPfaPO6Zv
H3VUd96KzXgBu9aO1prpDMRGh1fUm205AJZwVSu2UAqSSliX4qc7xfibw8oBGTbq
Hf+pGe7VE4ionZ/KCyHyvkfyZweLUYW9a4HPKxfRrwkCB1MNrtQ51jUYCiSaSpBc
sAcWdIucacJeWrvPC/bIp8UyQPixhAG6IJ81TBior1SOsRK/2BvwhvZuZjwJK8Nl
JazwLTS1hnPbejqQRME5UL4/np+BYAUal34IIhncY5IuY3fA49Yl/FzBI8wxoRpG
njZS2cdkKuVABegzAY4/x4ji2s50ectQzDGMmB9wgBIb0iLIL2lYfMbUjqEHUcnA
tcN5Sv/2T49K7jzzOkKzOth7ZkTB0cofMVjUXmR0UetxqF31gLe93asTFeVzFQPg
YqweG0PA5kllot94KCWpmVyOc6GNFlNd068pyGgNN/LxEb8yzc0x4Me3PSo4HbTO
0DglMoQnraPmfKhVEM9W+8lmYylC3/Jk9LQtheRFs0pv1+du2jVcoirWl0G8Xprb
0oA+lgjrY7QQFxSfUlxj9cbf8tUZcSYt84kJDI1LXn2e/STyTBT+hJIWkzi4jIXT
osGtYmhOwFXNXjboHFCmPwdTzwIZ5NE41kp1eF4W56FDzMC3Eb1yOrFUoD572v7J
odGIBCGrBd5pzAbWLTToWq/22OojSLLCu+5A/JmBBt+7ScuLz826oEeIBA88WXNH
9QnJ6hXPscgRWNsrLLmKlW105zmKuRjLAjETIswFSjuEkNsPIsQVI5pvF1UnzzPM
jvPUt4SWOQd5UAwdzRLJ5pYtMkuBZRfOJWZ+pC0bwj0RMt5n+FYrNS7+7mSFgsx3
4uREfdGsdk3/MUZkeLPIJpa/NLXPu9mq/KLQgf2WozpPHdWTk/gBstCviIu3oxS+
u4lf+J/NQqdhh16YsNnziDSTW0iQAyEwnjF9fBfT9G+EKwF3rVWm69iaTQU949+/
jVIiJvHsMbJiatI61Tn3n09q2nZMc92cGf8KQasT9rvzkyEKj1x0bbt5ERynKWUI
Iyd3/l+QR+cUflS6f1MDBcL9kwwojENr0PdlI7KLgAVJsX+PSKy1jCVu4s+EzVhj
KkmOEsd4AFdrmcNhSQ74KFggQ8q+VeZp0SnCg8CV+XjCWFYQ41BLLVJd0PY5+qL7
LdBzvv+xMwiS5PTDiELV41Cb8wXpfv1aqlAxHtv69G4BQLTaeCCsMW9Pbjxbzxse
xNJ2ENQ8+m6uo5XLOiLrjfM2QR14XmzKBHESKa5WqnNpPuJmNWLFDRw/XVO9Ya+L
iZdrKMIJol5QIwLAIC+/nGkS3d2FaAc/GLza7HIS4O+04NxsBpf4FzeB5DNhXG5n
8iyn6yvB+f82Z0v2+iOiaZRBHdWnQxFiYbWlDd4yZ+ZzzOz2orez3Rp4q79f6tZc
BbXluolkyt8sIK5tNPcfXkdQIMpi2YGnDhvVuyzL77gLEQNMaipoHRs3vTtSz5a3
KHeA3Hy0M+rybmpqDhJKskbC9HGRGVo0eQV1gG4p3b0vFd1h2KPd83DCqzLslwNU
uJT7QGx9pYHaPaSFiQMGkbFDXDrPOFJ1vzpFVzSCAaYrExuVux8ClmsPyhnV1ze4
u86ecIkT+FQn0qN3yZPAL5KC/Y16LFk9QnnVRmv8rcMMtJRMkXcQXl8A9dC3weMR
X4V8lIGTkuFvvY/0M2NLovumxcAAo9l2BbQzHKqfKXXLfeUsQmU5PcRbDxqksqxp
4xvv20ZKgK4VPbdd8RcJ6NaU6yNrkLYv4lrI+YO6Zb3m97AYqio32fZ4M7jj+QWn
GtjryC52JazAMFj0SnMLzjOKAFnYj4Ai29TiOwzLn964pOxNAWE+aEKmSZCjBCpY
rYZr0ba0K6MINeAIZKxeBEQ0d0Jcl9275rmBAglRKPdpzkWqBhCCLC/z1WTp51jJ
1mO20t2FaCaVg9xoaFMxL2Fc3ZpOTDx8/9fPYQpIL3bxQsis36jzUqT6pWjzfrky
IfPWTaQHfmc7MMuhXapl1k8oeFvJxZREZu+SxiG7R1T/oJE5RCeu8qghb1FPuy2r
p7/K4WMvxDCRsot+/aF+a3lDbNo419/TqYaR2iO+R/y+dKIFWylnFB+DfZMiZxDM
kyap+55MbXXwbN3frj7DFZhkyiJC16KdxlYRAUV7YEcqGzBXiv83sBUDCrRFfh4O
K+2wJs1Nx0vL9lpnMswQouSP1geDlNF+t9g54axMJXIrjkK5vaorT/cmbQ1pXRlK
qBUsWnOPVg+lGe05lAsoYVrGS74SPpkw4SHhtaDXYbjn7+Q78cOdsY132U7338xz
02Gr2gncMQ5DFe9jhKwVlGRteDuuC6zwfCByHSoOq79tCqMgOrKKFk1/6nPrLJSv
mFCxFW+TvAicenOtL+XkqR2EQgCY23wiiex4otI6R6g3l9Ql6b/WUsBbemdU5D1m
idZgdMpYnFBZUC4E7akqqkYvSIFZqyXHPa9NxgZW+65FQkoCUA6eyDlEMNkIlrzc
x9qImV7QULWAifCzoc2+tEmEu1ogdbwtLe4LAaYB4kHzyPlVFutmZVCL6AMJ3KOa
YzaA6q/qRLHDQWW038VWB7O08dfrihVXNz69509DBtX4Q5eBVlUBFu1APToHDBzJ
EQxeKiuhtvkLNE+Oi09/JRAZd9E7tKC9OoXCiMR7aW6ScMFxJ2dHYf9O+DYzQig8
gRyW4FHdPKhbR7xrTB+nafeF0Gm+xS7s4gNCr2GL6IxaNaEkysimto6KZ3d5CRrl
QJ6sUqapuAjordU7wW6qmefHfgFmG/9TkJ/1RDkG6hen/WaHDw0ET0T0GtshRfh/
gpHbHKYHSn0qMQwoo0fA5Zuy31nnlJDfBygb/eESpL6QfnBXgRvhJJ9r/Mqb7ClQ
3xp9L9hli5IrxrtO6kG0xed+miIKuTLYXAIEUPB+RWomcKfQk4N90DqbcuSBxY6r
YTlkFEFJPAlvkpurgTPeRA4oqhaT7K/jIVZznJxXmgsoA1o6WX6RkYDMT/W186he
vNt/ikX04GH7eQD6ogH3nYXH7IA4yK9snHdRmDd0rXf8XNthw4vLl27c3nhzZc/R
tPlEN7d+j/LoEw++i9yC005RVUZgZutj15a11DlPFiYOksqsxgVGJDQ5ugnybZ91
nw5yTk09V3P9Uhtxn8eqe4r+T8It04EH4HPz/KaIGoXNK3yZzYVqRZfFqGIxQAzc
nVkWwUVFVo3iVI1vbwbsrUVLTCYtBSfrO23q3o2tT/K4sreiZdNhr727AuwA/kQF
2zdAkjwnD8Rcu098lkPXwQeCYuramC3+y26rQcovxcQbCgQDgDE9GatY57xrtdwq
DLPEXQuwL2aIdRRhtmgcxjpGBW8RZs+8XsgaY39DLssO4VgJQxScEPbX9tUh3B36
mRp+liyNryVgOzvT7U7WW4Ab4ByvELXSZtxD+bDuCrbDMbofXNOIIl5dbAnaPgIQ
EgU4Bl7ZC5MHU7Iw2TfDzFCjsvt5K2tYzmW0XYvzeLCaXBJKDZbozBcWkM0KMD3k
TRvMsyelPdJtznL9ciJ9a5U9pqicqWLbYVw1xFpND5Ko1w+bne3FXnwAsPmQA+Xi
EO1H/QRdoCqxF2Awd9ZH7YVDGB8wJHITKJbU2T0xsQiWveMtRh4l60HcYCdbAJEk
IdP+sWnaeHJ2wGDAZxvl0AnaQdO7vy+W15LAdTEhQZbJiaZ4hwdplO5X+b+qi+cb
9gQBRUctprrE6PXLKG/VYO/a+vrKMcn3MhR8OPbJWkdKY0hcOtfgckN+Fub3SeYt
sqNPnpzRLVYwsAwCjdIC9CT4fWC2NCxQBroKLfCMUiHqj5rp3rXvxlovKfzuul5a
oMQLa6UXkbWF+EovjBA74d6veQW99/fOiYR7n0nMQSSbqNnoI3JPubGveM1PXvpU
/gK0jaYOoDyZT/H/EntbJ2O5cK1fIAeQT+QeDA8DyPEuRTIfqySleZHAmYOLfO2l
emZW6PEJxWiMs7U24av889ziRIZ/olf8xXCs6bEKkT+YacVJ5IRHsiFw1cIFEfc2
CNmxq9l98+xODyzrJbVDwX7q5U6dDrG04Xd7lN/6Thhfkav3xsmkKzP5Ov2ac8gG
VrPkb/L0kd0sQ78Ova77yiXOkCIX9nIC68Xa8XLlU/kVNKqlsVHxNh0g9RKF6v1h
xTU0OB4Q0bA+/DsekD/HwQ==
`pragma protect end_protected

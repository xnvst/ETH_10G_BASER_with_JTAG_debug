// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NZohjn7F2EKN1hlATkv1bMKWCkKVMfly/PM6bxbziTHHtpD2KTugmbkbSFNM1kUO
JdjEeFtcous94MT1foCwFcVV/PvnzSFZqyd150fm+Au5T/GtGw5TwZQ0I4+HVzmi
1clvbyYkpPqwIuRHvPsqr0+wbBWLyTvNWZpyB3k8fxY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8544)
4IpTRyWYphMOPQ6eTsvHpZNK/bcO9FOImNgR0IIlmHVShfF0+Ot9r4Ys7KD5rM7d
/CEtELjOxiiIFm/y1HEr8EOwf9P+uKrOxswBYuaU15UZqsDNyWAJNzkwH0yBDiq1
kJSZZ9LbO73CyYQ5Dkx+TvCBUb8N4XBr5HECxf0+AjCkCOVgeq0Y8wnQHbfXFFnr
nTd9qrgSVTchSBzzje0FdAnMIWvIdam1lMGBJylcGVjpxPaBA8rxzQ9E8T9uUGQM
lBqEYR/1woPK1lNUwOL47L0YEAfJAa6LFZneqiNmBLv14dqPXUrntuprTsX8lrMc
ket6EKVcnrD+aLJIdDQtmCM9jtCRP4x9xdtq+8UoD0qErzCSlgZJPqu2U0F1cTAM
yJF65TZ9ZTwzCS0e2Y5TYReZm2+nBG2/zgRnxxVMFPBHloe0wKO92btc5RZlxa2v
LH0wQaQ6vDVc3j+jMtZ6wQLhGi7tg1cZ9HVbjoBqpIePKgmfpEfs/eIfB/LbYkf+
w+DxNS2WTW0IncwifYQyHxYUcDlIHhOn0gv61SxNyHNVOFpfcsSNo04D2IU0u3Q0
91WH3EWWLV5V01fl6d12XlVOyy591yU9kVn6chI+WLvlN01q5gDWACiBemrQCZ7d
a46X5EpL+yS6dIS+/ZIjKJEGl+RW3ZtDvGomZ+kSVtfGqeJXRJZqC8hKO4MAtojF
iAfPl20jTYtfaJGzuagvgIM55kshUvmo+JgdfDf3zD9tFqwmvkPbpL7kmdP3kxWs
O6t+psOwfKNTJVNgze8v6Yyd5//MSkqQBXnwjOuWN4j8Sc3RjCrfuIT0AAPbsuAZ
yS6LaZtm8s0qvw9vMTlBmAVDQ1l5coFx3T7QKDrNljkSBPvftn+Byr67/+jyOKFd
B9SxbqEMqA7tEZ3/2oHb10YiTzGjq9M6iCjCUePUKEyFNJBPDefKRkyIjzf3tDBB
AHfaBKOeiyoIMr5K7r1+nJFBnKlPCWx+OxSTi2mCTwkd1sITRz7HqixBnwshgdu7
r4ss1OlCPE79UKicMfd/YCRVfA99yYtfMX0VHRkrIZ6ysdKo5/HGGUNkNWoF+nD+
2qvlxuZ9wHGbSnH+KygWQcMg5Cp/VIAzOeaS1YPw7JXSjS409OnkHfQF1pxU9vxL
2xOnFZDNFV7nV4MdfprONJnR82JqLA8R1flO+mvcNom/FSj0dGp0/Tv0qHf1uE7y
K/oiXqrkTwE0n13KP19UtW95N2x3S+HPFksxgnwSHKFw3yvuu6pmZeZRCPu1YILQ
7lk8EvmVRXc4GOXgCea43o0kY6lEY2OXkb0V8WcdtIlpSO6VTkk9Ljkgfvm+oS0+
WA9/OT9y+clAdvfqmA1a7WKKnSdMMcf4fonT0YBPPLz0BQOZ+Ci3z/LNxP4hraf5
WrqQD1SRd7p/ViDKu6WnP3YZ8A4o97bQHZfP9yAEiKXrKRq86uIBaEB9fVWqOc2K
HztttfDFsfhACBPwHLTmg/vskiJkvTihYJ9OKKTfUq1cIUSo0b3C+MQ3hglzvQ5M
HOZDJD2qk3aSLmcJfJrhwjWKMK4hA1cj75oT3UwxUHsoUCqqOHqhOVyNJprUzrDZ
+zxc8kc0q+oLDecFHINFdPw/toAAQUPVQWy6M6Or/DOHpfJiXIs/Ma0ItluC7lzz
qICOy0H9d6AdwyDfwHbKuh3Yd2Ie76gHUK7jV7x5HtiAiP0prBZ8yqi8uIDwASSF
rp0pVoZyaG0IDJGOH26ZJVDkUN7po6qLEVK8SeoQeXp5CYW09cJyL97BzQ/hnYUd
efYI/itA1VdMgXRL+a8oP/fQQF6EBGc39vU8W0dMgSr/+HbMaT0UEHWhYaiDZdmz
3nuERK4fG/unFUKSbuRtSjQg2GBvA2+KeSWLyWxL7ax2K4PZefE38PzIFWUsRGAt
Vufkjcbff7fQ312gyUvWStnkzg151aMIg/omc29Q41worcmUirLBWJ2CwarQSWxm
ZT4HMc2jlq1un6W5ZPTR9wuMJnIoEKDVt4WWuuWogEFHAAku1hbzlvseqA/x/vat
haaKskLcoUuDizaJcbfqlpSqmPIdPjo0vU9vaJAVl6XhkdtsOuhzR2eLrwYdmeif
9YvfqwCWqCkkVD0DpcyJ1jdQFtwNasVXJtFOlmkvlyBFBD2ZvsXNH+IJyVcSpwkT
unkVDu7bitTr/GE4zvZRDFrH/pURMZobFs4d6E3kzP6o5q2fj+KizLndBH7sQWOt
mQ6tN9hrgN9iAdl1pisTjw2MN1ksSYBKXwxhsH/YBb1XK4noJaW88gzxLbDDHKmP
/KUrAgoh3zL+ZbV6vRgGlvvFHj55HLt2nst0OmxGKb6xsQz8mwKtdYI6nFYZGDNp
AgLEvs5TrTJpXbz7pQBsk1Ngw8n/PZzsSjHH1jMrHdHxWPCn2OK77Dtm95pHcGx8
1NikM4mZ+n9g7F3QIIA2+on7o7FD1tpLEg5n21nAgLUUvtwza5RttQQyEVxPkOXx
ISejn+h16A3m4ypOnhrRFjPsCFc1x1YeoPMWHi5eqmROCvBbfEFL9W4kpu8x9spM
pTL7yDZ2vzce/U4bGAna0aWfKmDTiashYkiA+gAIKDZKG4CPDuD/lpd/QWT9Q+NT
IKGpsjhWZkivosEeM6v79gyDsuR0WqF/eWKEIWJLc0482ki52uv8oVTwooXoExWa
lykN1jzdhNx4lOzm7mzDz3wTIvJSC1Zt1gXvwpAQxTP/A5I6fbvyiRlb/WsiQtBV
AutON8Xo6e7Js58sBlPciDdmWz7JRJKx8QzeG5ySeCgb7rvTFwosr/GIJrzdhsCU
AsezvN7k98U/Rd+xWpvEr6oJsrfY3LIvwuAmpEhKlDbyoEVwR/+wvEzBsRouolwm
lagee//fVTUEGnAvuRQQ2P3NlbLuEDdJwjazQWKXTKxJgIyW1W0xJRdidv7H8dhE
Z5IkFcLYmI0BdxtswyICK+Xz5fcvROiAXTqT3EQn27S67cEAyFR7QArjKoAwhfGI
bx6CfbFvC0zqt1TsVQCqNj5UzaiTU1MRe4KTC0lpuX6o1HatR1eEJk/r6C3vVuEn
71v0mreTPLPJp8WbX0I1kFbiUMYPDyzBJUtsk69s5L5ul57k0l45l42NoDFoxDwy
fKBpwPHTFip8J4UVW/LU+chiZk+lqpU/m+frkiruh3vwZ2I/FCFRrzFzgvQWg6m5
2w5g6ryHzUjvwOelMALw8uY9H2X2OtG1sPceOFfDoYOLHxCYbgcsTVJJAVK9ieno
ndIfnp6brB5guR88Jas2JJOLszheFWEWamFmnlVI3wXWv0lR5HGPmeHgx+bMMluU
QKpCwGIZ0qaQ3JV6gNbage/ftq3YIEiYa3fKTd3x7s1yG9TMNAUmpToMLIeyESUO
U7Yrn0DBQkh5xFhdotnHrkYkJ+Ep1XVi0RFHtBfsGn4kmIzCyWC6pnLkrxVsn1wG
ndMm2PKrMfF55XrR1nm+YJVGnpA+J4/ZVy6EmKWBTBxIwWhM7EankM2+KB3Uwbzv
qagTbHX/RC9t1wFBUwChEvL4AsUz2QnJeIeGT3HwYpr5CJWPh81jFLGZEGDne+jF
NPiTBoNedidzFtLM1lqL1BCWZbTUMqdz96mkhluSVHOzxW6BNWLF2m5UrbWdHsUu
oaOIP2QMu38IKyhk7+qRhyiI1E8TjdLizE4BAe+KbNKOurc8tjZ0uDD2siioQHa4
hMSqN0A5ZAVPW5d/yTJ6UZfAcP2HUd2un3JPx0mS0HM6/+X8zdyLHYpWFSWdoYC3
Zqm+ojmIxe4RWO1b1sOUQunwC2iHwWMLNmig+THOsaS+fL+K7kQZM+45U4fp8JKy
BNdgJ3bLq6TqBIv1LMX8Dy7zzCuaiSp6GEawBIC5gVRTXhaPdEoumyrDSjkStqX3
DTuZiYILyuG/qeJJ8gs/s7HbEZTMjXP6vTgaJhRvEnDGfZU3bzQfLZ8mBfbCgA+A
MF2nfgXCNTwQbj/sSj+BbqEM5xneNmAt8HRwzdWKH0HlDxQavlwHHMRF1OZyoAbl
6NcQdHw4ljcJh2EP3T0ugpMt0l6CLSQaVJWQba5JUrWsnHhvetAWTd7ND2TcMXlE
OEKghk5dscGEkTAUCn8KguMHL+tD/RbgOWp13DZVHj4DHWpHGGDx2rg8DdMpIPb6
DJLPzvzjJ+2OrPJg6PfosBLhPBeZdVHa8M59OrbezXpZgeNRdE5ernDT0OV9Xv7Q
mWL/a3131sDn7hVyyKCBbEh3dS2epT44vWFd2x2XfWA3DwT7JS0UVZuWH2p5XHxT
bJijzRTzEiRwVGPEU8qmPDyqV7pbgcCn0EX3LNQyv9RSJXn54b4XaBDdK8J4Bpv4
bimPlvMsE37r2KQ+q//FHarWrRc055orThVPaKIZqW+5zKGW5YiFDOhy2xjq0Uk/
SYpTbRSPdApeSZrafoR8L7C+l8I5ojKOxryQP8643gfoJBmkphkKNuNqCS4+RuUO
obfBjqBFLZOHMOQAK1CthYO+kDFWPQSOQmU/blG5H1zmb2hZuB/jGiiCpwCXXn8u
3max6HY/PI6PTjfuRgi3LiMiFLHCNki+PzI4/NcfVoPvLik1reMwL4Mx44PUMGpn
gcv0TPtnt9OCx0bykAL9MplOL2xAQVXRnHph41dqvcNj5m7WpZv17hG+TrpbYaZb
10kqz1SF9omRkApcJq1THL9v9Bg90yXtQO0PWN9CvnN2WWpgBznKiTvZydz2SdVf
OPJYHAc3RCKu5VY/Y7S+D8EPiHGUs3S7LJpo6Fh6WAyVKzUM/VgSaIexSPG/UckR
jnoGWTFtTJUmSMdZdUkW81Ba//T6UfGTpeYfL7Lf+ygwoBr/4BeUq1Fr73s5X/FY
vpEvhVEEEwYY0U/nGJRlzWhQs88u/52sGWJcI8oKInfXTrI+cQQp70NlKQ534obV
D/28f+mNjmQ34uzchNLUjiJfJ7gvUl0M6gXpqV2bmBLZX7QvdNZJvyUbnW4jIihA
oHJz4ujUYHI/GUfNvlMKuGpWp82+0mlkgo7ljuCpLVt1EaOpfdHIVppjr+1OkdcE
ZuOFWomOmFHYLE2A2WQZDoF6TPy6ZhPfewd3BobDlmlIXQLfEMXzuk9UrlpLNgr0
3brCICyhhvQVcjijPvgRxP9weSILY5cqNtR/lXSFiVLNk/zoUV8NdLo9zXy+kBl/
GV+TsEygdJoh+DJaVCsCJ1nENIaM9dInoW3vuMQMN2lk9wQEa0xFNU8gIGNUPNji
BDbw7XkJcgG2k5EMClsU5JZrxDyKmr4R9naueTJXasD7AOfCe70GvBHKz7bkIw4A
DMYlOdpDzW7RZgkd8NoF8Xd1ImYy3hzn5fK/RnxmpiWrmOALL/BgY7Mp4MECxCQP
743kFokN+CB519LImVuUKhVLcEZ81buj1v1z0rh5vN9SNhCMof/+8glUVSqiVHCB
uEe4I9yklqp6ph8E4FsN9CofTdvpHb1eJafH1+4F7Qpb8tDdRFeYRzBWxnKoISlb
fRwnxo0WZOm6JRjX00GkA0FM+A3QlQUh2iHilv5KPAkuHp/UsCijUoruclLFSw0F
S2bgfhqa6s63/JXhB+3D+Ias/MqDcUmRV4ckIY/Dlwm9ncbVg+1BDfKF+DulnRqW
9REmc3hAajl+N3HwdZhze5KGDeVbeY1VDtSScDV4/4E2GUG95mIaBohEyJ87zFH1
WFftYsBSB/B3R6PpcagrzBNLK8tVcr4Rc3LTECflY5ooPe2bnH1w/F8i7Tfu+d1V
DSi0LEBdN72CsmR4uzI7szAmTxd9puGX3dOwESmID+BDatk4qKAWDW3Q7m0pQgkR
unGnxAPBcUGM3cd0MJXygeRHakMd9Thb84t/bu7AmGWjB5wA35mRItcCoGuMap5F
e4YvnNLCcI0JJYArAcShqmdZKRosma9lyHp9XwsGKBxwtwQEqpTD+54sGsnhueOX
gH2XbBFxAmx2E7PhqULfJiWitIjCYdbENHRSs1ar01jVaYUWrwjF6bSUXyE1rQi1
7QelGd+8AmSX8jLhxY0dPNLd7S08Yfx3V3KMYRcWuCHKOnSV0JSlF8Kt5aOfh/7u
rp0b8UatiIZcy9Pw77miY/9Rqgd8ikXY23aYLlO4822cNY7rzMT6NVnOzwLhapIP
KVtW6gWeTF8n1u8IWCJp2bfAj07WejXnGc+PHHgnpKQ0OrDOOXzgYsilbZsnvT6m
dt/+w/kIQ9CI6642mS0BnMH2UaPbbDWqkuw8RFHjBCAfcwxDkwFqlSy7MlCWRr8o
aWh36u7MnigP46nM1xoslXjCEODtYJIA6xlCCwUVPlLxMz9+5rynl4dVfkmXjkb7
Moxsy/Sjj23Jl6a/gUjaR8qbMvKt0XIh3COShAmCvC4xioPVzGCBlafe2o2pBXlH
d0edLfZvgzdGCl20HUMKMhX2Z8vWgM/wP55LQ1t9SqGPY3zyCdZ5+5YETF6XNKxk
mUAJmaBQiv0+7ypewtYgt561ph2oYrFlzC7WQrPLfLgkPrT9oa6cua9pCntZpx/o
s/AY7tKZvKf5TeOhEXabppJNfK0dCogQcpjKI5WWL5Uod46LXnD6/qIQ4KhjxxcI
Hpu4Uq6doFyYEQjCWE3g24Sqpr1x7buwRy4ntYjJj4YjFqk7OIbChzZ6Rsw/7iRC
MF3RDtEKdiNTBo24E+q8sNTw7OepYJ7j1LfA+63OQNPyNsAeyKX5QRZdjOlf2WHe
+3Xov8OZqMi3RzQKqAGKDZMJatrx6wbD+66Zj43CM8j+hf9zCQC0f/gaJ2HQwd3g
E92TA/xiXIC3PaPjam7OCm8Egk1ny6s0UHZXc1zk6l0Iu27bzKHbWNn9lGLnSMkg
8gl46uPz8tl6UsisW/XFF2oC3oVvgZ4mpWg92EWwrsiY90gCvVm4Aj6ihCOiT0Ms
jaS5QOjVsuXqm+9dMKZHvXfHWZFRscBAHFrftB9Xa8bUIesqmCOsk/+WcaqeZhLy
wVc6sjGsEa081RJ7XgzcBYC9MG8fwbOUi1WHPx2HksTjZ97QK+haS+iRg6lci8ti
RF0EH8m2Q/TyYlUSsCqLCqcsj/vYW1SWcBBzQVXUDl0wxCOKefaoprJp27e6B8WJ
Jrr5xQunPtP2cGhl0/zrE57NLkKgXHZ0ZJGHFyxlvn5gnPaSE0et4AJDkKP90pgT
d5Lpt/ux5eFG2ZcmouwwtY9RYCGiO7raZhg3Xjpk5g1Eid+C09tvO/nz9yAWn87I
vJgejwef2qNaqJPW8zlmHQ4ZZI95P5Q+SA+/AqmMPBa+PDvttRGc5O3XwXDauzQ9
M99Fa7c8xJVVzJtCTWMq+iOIuszafb4VXzb16AhK9AEP0MdCzNhJw9nElfXqG8hm
6Me1UFhxer2spVzKWYfumndUesHQlOI+uEd9Z5gqw4H232FJlPOehsU9rpG9Zj95
OQYs1C4gYdo16Q/MjJw+ACw5n/tFOFLbD5AyncNFFxuJ3vHxUefwA3+Z40IjxhW5
Otdb0H4Yr0yZ8P7z+V/bf+/HRpDQZMlWa9FyaaagSHF+uJTEw+2+YyS6BdhHxqnv
xgMVyr660Fe0WgVsczYTqowDNHKg1cH2jb9vUWv3kWP6plB5QQKTsTesVNxfanI2
yreFe36jD7J0dohbUg3zSrjztDA3ZEaIHivsQAJ2Pwx5gE0SazY4ZZyfzh99iRss
IFkS9vkEseWdH2fO8BSdPVDpN8+E/CymlclTMgjaRWURZ1ELppfJ9UgQn8+PPwtc
mS2OjY5WraBvmgZ3NDg1eYm79sOplkiWS72XUevQAEX8Tkydw6Q+n9/3b87GB2sP
L/Qqk8Nd5Ueggu2xc14LVG0EvwfGY7Vq1ZqW8F63A9y8oRy/zzqMLpjgA5RFel/s
UmN0AmFg3kdIq5WQ96jRjYY07PvAWFiPIBmgzBqAqjhx8ctt2yTC5P9cyKQa71uX
Mm6xuNpQOhHZHI47L13dtcQLyTQ+fp66z7r2ZgQfFadudswCHDb4wNH3iJxBIKMH
jlvOD7EZTVhLP36I51qbdW2PL3SUI0t6HJgVmqgswRuRxDwL/GTSDe/fqmu6El4M
J0f4GvChhPfoe9RMi3x/AYJW2DsmrtijOz/cyiFJdnLiNv4e5YrpIPqlB2dtcpVm
f+sNmJwcJagwYk84n0NujqhYQkt/3uReQQ4573gFAvrP2tSa4ivvZNta1iU3zv/c
jd0DusHp+Bp8Ju9X+z4JyAA70vdtNdgzXG+Ypv5xk2hwoACECoSoj2S4g96EzEyJ
IbFpCwnb1Y72zZ06e3geEnIuH/iHBXvw4hmbumDFsXuNRvrZVYqBQeaj6iGh50Lu
laPmDcHA7ix8ZwVGExgzh/In99+HfoSx6ytgHobfgT7a4ySu5xtPSSzRhvlHi+8h
M0n+E+szANADxdSLrS+DC1PQ7eQ5Fwn51zNgekDQclGJwhJmqnhcqFqAXW0Yx3h9
3qExSwuD+RjjjHt17vFY4U/zzCvDuoPYfnfY4aReN9Ld6o6R+tin0QMgYb3lpJbZ
XevKeAB5xGWBvV6z9swb6oU5O2+nqzgaU0NkvMsza5H5jpRjI8wSS0zjMSJ+6zZm
KMlWhzX2hLV30wl9sqka0szDFDzmTliNkG0WGwkTKo8Yihdn2F0VGrop91XiWGiY
bjfc9gECDE/yuZ0Mwk9uhIif25Z/BEC/rNGuFFMFPizMBc7qIGZ5JwR/pmnh8du/
Yh5mDBlxNJrzYvmo8OfvwkdY2UBBBWmko6dLN1UC2EqsXz8jQuuBAGiMIlX1EhVU
o2Oo0Czx9uaa8+1FDEuJT9NtXIr+im9pw5wGsy+5lACzE7gq11CIcaqgfBR2X1Ce
TdHoXpm6YKF16x4wLuKbS6MH2nBcPh3XBzc7sqGxn9PzglcCoY6PcT503fJsTUc9
SEv5xnG/hDWY/j8wVHJI6m551V0ZC4mxN8lEubS6s2LDmT7dC6OxTDGI2T5lHvlA
oSdQZLYv8v1SXVxJLgJu01aQAlFDTAC4CVrVAwufCO8LWmt/az2+cGr1TXXWMQIj
7VuzASUYElz1UeFQASJkUw4mRO39bS/LyuTdHwtTNOv85pGXeOjCyZJNWrZBD+ta
fwP5DD8KCy+C57FuajiRyafuwZrcad8BqJiGJaFVMgpjrrA0+aRtGNaSY5Sr3rf+
CAwmOxobatn+Haqk+eFGFMlzdpoQesCWraqHDdJuL/j6oMwrytXUG1nNgute5+h5
0rfyruQlNmHqZGdApZF5nk+6Pj1NaOov06c7reE3YB/SQKOXEe6D4AXZxzquq+wv
RWw4e7JF50LvaZb/3+M/Q6hIpHLeZlrXMiTSzY5ums4gFSa4KM4NmOW0GViyDSgp
CAsAjwqapw2SQ3QjEIzJ1cjPQ/VxykSgR072E40fP+t6b2PkVAp+MARdRXmwVAyN
5al7GE7KUBg8jrTKSiXHyI1nXxOjqI/F8NHA/4d/eCayUieeFfc59g1CRgkYCRlU
RHhifmiKIyPhKu+yMAa2b7hhqONxSialMNTZ/kX6gm1NmatwCymSBsp0eO+zJd5/
TbXFYdP5+MbhKs64vXFExKTrpaFSwdkCy6IWjP8vri6LOX9DmzmgdQWvZ+y0kI2a
TSHFI6e74ASpCwXRBvaPOwxm8SwQkLRSNFkVl+kVo508o23S4YYVBATVFSBOL0ai
UtAEO51J9v+du2LDbO0CG107OJDDFmFKL3KB9hy3cvWf3h2yX+/ximpFlvRPqTxJ
PwpEUvzSeJulzGR2hqx/On3Pl8GjLxlYvxdsGLkPshyZt0JGl4hkiXM+SfBM3GMa
7UrynPRGcEjV9fMEI1wy289YJKIP4jqTHvbHsfdDRYD3qxCNgvg7IcD3QCD1PSI/
yL/Uj4eNyX95ekeAUlE6KllPeNAOivMfrQkdwxMq60R8GFg3KMOEDNJ+RDF/K+sJ
XeC4f8qvPJet7olpKQXfMP1vzrNN22Ae0u3i6TD5LRjYTiIGqACv9DIyYOevzGWc
GeTorSvUN8mpjyw7uwJPi4fn2lwRgUtwEjPNzdTW9/Wv6H08317mj4M2TzHu997G
eyflE8Rud7MIU+89uZMfZfIZRu5ezOZb6iLmTV8dBVoj3tFxzIDshfmGbyTitUHD
h0TdbRu7eU6nL17FkCx8P5k5bTUs5rSxZlbYNs7sR9sRsu6/UBBMXrrS7MKCZdEQ
ClMHEAykyyNJzNHcSaO90jv8fvw0MZvsKX5JV4L1eXxU8YVVPCeK8rJmXrnWswkq
URWPBmlOQOLF/ysn/gNlZlKgHPIA5CjODwvgZs0YRqp3woF1cayDkiLpZ6sCyaEp
VrecXARbq1/NdVbQxegx1IdYsf10dywC39stFCHsfkeKYgHYvgTwa0ZjEVBJ0Zum
tRUgzniJzgG3YA+IZ2jMoCMYLosiAHceV+FcmGfCIUQMvi9sw57X+48hDKfnEV+I
Anlb3N8M4AXF1lfG2PYozqX+DQaWkG70fqmxjNGbhv3dImC+v3RD3e+vDLBN/eS4
7KX34dC2lIyY45fdv3I/jFA56D/peH4wbwxt+NxNTcF+Mxx2lOEzivz/AFblT0TD
MssQxwNw5RPlyHjAWBWe/Sj/OVa2MNdVmb9KqmDgJq3lI6le5I+s2c/4MrmN4074
wrIvE+QbagYH08k2iD5E3SY5qn2CuRaSoR487yxA+4npjOoZRxA9beC3zysdKmdc
maPjwj3680YhVtLVyxAMJtOIrktvFhvq+NDzpoCsdkfW7wkAFeQbrV94mPlAPJ7t
ylFW3/Ade25nLaMpUZISxPxfGroIOz6YgNCPs8sqn7G+V3MROaskz78IM5tZOX4E
yFR+X8505NvMY9nlXh9L1Yj3exi4m5qTbObtr9YYRja86+fdo1qRUywU0QeeJDnp
k/XsQctunhhMC8kIV54lklW1+VSAaXw6O6p+p85kB02g7eBqlCCN16qhStNprG9q
U+RroXYj0RKzIhFAaNLNS0kW5D8/wrw8ufXgLxetKCWbXvuP+T71bqXuJ6lsrrN1
H2LmVLUl0Je/Jt2CD9s2JWmVnIdn3O1ay3BkCRehRkm34pbDst4F9ytNUFSFnfAW
QNX9o67pL27GFupoy+FqCdjlU1AgYNJ1n5/Oo4oIDjpI/ejcpCbWBERLhEHBvNo8
At6ATtDAsNLWBu0iJ00XhXftzSaI2+XxlMwihhqLHwDZWv56w1/6H6b5IR0NgH73
Sz83n9bEeXaBJLorRF0G+97kEvHDVIilmMd83H5n1Kbwg2RljeZzm84up/h7Gsqi
UZKt2nVOHHNMvgkywTyXUz9Bcdon1lVT+Ea1abSV2o6RF5G7oxQ/Zdipp5YF0k//
HflTtQUmim4UZfbREJCRQ4+nsc3D2YEW55XMqLczSg7WA0bo7TNUp9QUOVsPnc1p
`pragma protect end_protected

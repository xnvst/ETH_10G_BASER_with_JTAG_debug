// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:37 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZSeuYfiHGDaoDTnHD6jp9ogkiD+p3RyEl2RsFutlFJcv0MhssOo2pL7uN2+TWnA1
OdsC7Hmqzn0GRvazk0KyG88GLwVLLIg5tahFYqc3By32MSuUoH0BoaWqzlZN8Wx3
WTdvYChbJMTI0dZcAuHZJNA6a+Sl8lf0O0iDrrfqAyE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5984)
Bi2iIR8Q3mZKqHbhXzc2qzED0WOsVyUiolXpCnpEf8me6LXsFbzZ+d88O/hve4y8
1QLsvTI447jwppOx/Q8VCDR3OPQTmpdEu5CTGXf/e81BqVt3rwvWb68HbJH8a7J4
/9yiMhLpvu4ZSGite1eZWfILXRTSRffUMsHc5XI2LZfyZF9OXbW6OIHdt2bv2/FY
j2h1pDtus735Gqkm3jbkjrVjdue/5JoRQ4biCaqlTMxgOc9nQcn76EwgIptlChc/
NelbHgy/husWBr5iyVHQr9IKO8wa0oLw5ZkBzbd21qaPTfEbTsEflG19wTO2k3Kb
u5ojKqest4/FrsNTFH3eo/lW1Nn9g2FuppG6/FaFEcvAxB580ZZtCp1Nn831vhtu
Tb6oUXhDgOT/BECYhxzQHALYHnYh5oaMYN8kzEewU/XhcI0GQtRZBD63dvmR44tN
T51tLbed6PM8IzOTJ1Oi9ia14CDveUFoM+pA4UbPvU9syypxtYulsezv0x3ot2vs
4bQmLLuk0XiU/3XqMd00ASo25QyLjgrYWMxWuN4KTlI+dw2gemvDU43Q+AKTc3Rd
6FZP1KyuG8v2ELK2ryzfn0M3SO5qsZSh88ud4iOz+/mcXDtBSYklMjpYjA61enpO
VhiKsMVsSO1rjrbyaj43j0hAlryjxEEUpi+HPq3tL0FnmY3aL6VNB3qL/kkGbILW
JpZXd4geFBf4ErzVLB+fhx+tS+UG+KfruGKFvgNAvVhpyJOFk9juk29owO3deTXf
zccn0TeGVnF3Wf1pCbHbR6APfw2i20yp1NlgzApTm1W5AxpE3VCPDaX33YJLFF1y
LCrACa9zWioPHf3Oy7SRWcOlOFcqJipyONtc6B4cYMWUzTYcXFHK1OTYJpk9xHxJ
L0/3hsAB3RBpp2jL617LFWR2BUyfRtGgqmlC8yCGzEbpV2y+ZetXVn1gVKhAlmpn
JvQEGRUBWVgXTyEmlyZ3rq+XrDqruFT0wlXdE+biQ+y7DVEIwui8potHx9OGx6Hl
EtNJiWPilTpLg7ul82i9byQxz+fVXaUMC7TCMev0CenaI1VFEJqiHpNYi6585w1f
5j1ZsXZEcqjzx1aOiKEXkCCcaWWz8DNUgHm5K2vJ0TPbnMEpX0DOb1U9zWkVdGPi
wJcllWvfmrhn8nxnO3bv0mBOhivnwluhU+Dk79lQYdZ/EGge9iVj8cx8rKF4LJGD
SBAcLU0ZXhDfRM2EQLJUqlp1ADfGZijkvS+nDAAHoV8kEyyD2EVVYz+nPKckJddz
/YVPrvwoV1rqDafKxCicQa7wTcHB/ASEEybU2t3PIU2V5zOBIzgi8SWCSWuulryk
3S0W6vX0oM3G60Du8rqhnH2qtLakhsikkyu40l5RoPkNzp3qt8IC7siy73VHjvGR
oP6ziTrxG1EeDqN1SpvKTu+a0phSwDKZz6SVJwCs7YQGjsQlgNia0uZmXRuQOA52
9BG/QQI+vko7CnEDJnzXK9vmm7bombymg4se6BhHF6j3kl2n3g48PIN7EXdQZ4ts
8iwC907RWYk2LiOdflRz0cBtG//xriP8virJoXAXbV1U5xvoaWlsqxoVnFH5fjrh
ZfJaJfPKKCSlf1I4Wx27J+22jgKKgHj7j8guD4/ueT9a0oHzCmo5sAsC19+VzofD
YRIpx3gWpf4XBrHrwyryinrPX6CQNemUQ0JB0vLPLJ50ixXmxv3m9yrS3mV2Aa0l
v1Q13c64ftVCUsWNn/rFovzIVjZwohW3xql94eTC4ovMnyzdwjCXj+URnu338jn8
k+j7hWp7ymuTvhDyd5wJhyVC3/PFAQmAvzIe3l7S65epFmlgzLjoSHwRt/aps9q5
Y6rZJFh+oF0Q/bheJ+wqDN4wP0TNG9rep7BjjR4YctoXVldIzDvIk5GBNh8xJQ6B
jwTsMwBENNXut+Rfg53KdpmxRkWL0iTNQhGQ5v/i4d2/v5TjNfmVT8Mjulw/G1SQ
0zSZsoUbQc9kfF3pAONiK7KRZraxm2Wqy/NwSnq/WzdkoVyyqI93cBvK/JOhDXki
K9apS6+w5PijrpVCSyIiripd+tCJW2Ywnp7AQ2R0NYZAiWiDxNvCAVnyRQqIbDYs
0zQV6402Dpn/3GouUZIh2ZxXo+1ayj8f8l2qRmMtmr3wSDHQvFw/iweEEBwPLUX1
Fz2P+xbI1yEaGVke6ShzDniqLQBSmUKHha6Y6GhpUPifuBMm6IdKFQ/DKPfWkkrY
W3hmVjsSiMww99ZVzI17mZHsaigwFfHo6KKZFSTG9n8Ql2mK/NfgW8V2iwfq6DKy
3VS4R4ql8hKylVmBP3robSHE6Jqtw8m5ojiRJ869Pz658b0HqOQHSoo+pkTB0MI/
SjttHUJAZC9iuA+1Cw+X/DGVDXycDQzyI3uYo+Fj6rQeoJfEqwr7Mxnbyf9NYkTW
v3va/q9dBQE7DbHFlPT/DQ+muATt7acSAaDYwptj3JUudE+C9uMfiYIybqLqkBFM
2xRTkgSWB1Ww0oy3RguVaEj0lfKHvKKnBD9aGJT5J50evWt77y0QpsBOIXkTtlkb
lvVMnqJzZPu63fd2wVvXlQB+rt5TckkdSN4kPnKhzY7g0TyazHqNPEdj5sEP0J2+
7OAQoaRjPPNkMVT7/Q9ddgt/WmwnQ/erUozhw8kW4+/WcmtVrDaKwRAg66rnI1wj
m5GrKH9aT2+XM1XTqBc/FBFcUp5sGAa78QdIxsuJPjmtyCZ1FdsvEAFtRP6VY9lD
0lrTVFqCfDzQjrOvhawz2r59qfaVnsWZ26x+2iYUo3BgP38XrlbFHa9sdjXzpHpD
e6hw5rk7SNaFdFkc3GAfTUImawvWNM+Bv4m+AruH5yITN5BqKGdz3no9rKK6f+Ue
5pXkEoFsIXFGrs5fNiiaicY1N7fcRMnKwKLrJarkGz4JqIqOVvVwUHvr7d84DXCh
V9zel/JTD3ZMwhhTocmL1LuTalHhC8ugl3db+UbmrnB5PqhyoolPp39DuwIlNHKE
8PLwx2Kufs8tfDuIjR9msRj6w4ps6mmi7ynnvQrnbn5m0TNFTxqzNiww5cIBuaFl
7jLsAGg8nSbh5lRG+ZqX2uP+9OYCe9YSTIRQu40KjhtRD9XW4z+349hztqscTlB5
NtCTWpNJj/nHfZ0fXEE56Cv/AmvdssQIvNWsFnwZ6sJL7z4qfV5Nm9JRJnItXm1Q
1WZxPh9IADMrl03dU1T3bhBWoeenhbcFQhHLpgrBtLaaS8c1OKJTUWi8uskeoSTG
4oXYuOJ3SWGZo74LbxauFk7NS/Y7W3vxEmF4ct2AErayGaCh2BUsCjdIeKXrso8H
zk1ED2dpBQCG0pJxSOBPMKNbVpoiY3K5Wem+61Iai2zIxS2qs2PLiv3ZAbzWm7lL
/Uxo1oYSdOYdJFZpXUpuiNA6egnBm8fEkdmHrSMAmVj4o7jVtb3D7l1Fd8u3Uuu+
AO2LwnSRD1OZl36rrOKZt9fs/XNdGtTFAsEfiYyibDvzF6uZHjmHOnAlMrxwkcvh
rB8h1pcJJ4ay96i/ZP6jglLvNzg3DGJWXXRCvGzw0gmNMFpnoJ8mGp25viGsNzm+
vjMBkzJfneUSRjboiPjxYzZeChhLarlDCTWnDfJR/XHrCYzyqJQI6b+XOUEg4/BX
Xsk1k2+FWJxWlVrkdsOX2oGOayD1a8lA/Pu2T43WaufJGeMS5wqJSZKnofssC7hF
o5ajb9rFEbX98wfDuyFJtLPHJUwhHC22ETaIzakAIUTxCrRrCfXMa6f5wFCOvrzT
NV5FoFIzb7bLLR5FH03cfIPDrRFVulMvuzBUXD7uoGeSerEcluo6YYCmF/obG1Xs
rLHcKlnT8bil3zyk5onfDVE1NylxzE/+eqmNAoVEySIfLoXxfhZ1KGxqfv5Ylrh3
9mzVYlKio14r/nBoiyDXzZF4RN0y2t3P2Aat3zHCHBVs7b3kjUBjvKAqF/WAJFBd
8gLIwFZyoaJCGz6juiE+MqsrP038EHaasO3sSR0vjpvviIDo8fjeQPdmU4I9Ny0+
7LNfpcs7N+VUuMG+pH47Hn0ClmMkkUxOJjkyNMecZemo98KH3rozwxPWPsBj68gH
9IryhDCbye08Lmo9LLCKwpu2e5eY41Juybtx7JtRq1uFYf6czw5GIzDjvUPWUujo
YJhNVyhHpgkVRvaq1NFKVoqzYfZxPAJsTSWzfylYCvTQzJZvOv16TEE9eYTwtVym
+6dTZqfcZqDlKpW45uHK/CHazHiYD18FbdJihSXIqCKIDvpLZNmJ4pM96jsmwHG7
zp8yLHKvvgA/uB3BZpHFf60xvCoBzMzN2ypXG4OsKm0eBrOisBaWArYrfw8p1yO3
76F320COTKgFEBS6ODcQY082EdRf8Kxx5Subej8NtwULQmOY30WSV6T3H0G9xkpg
9WSwzGOE44m/wx9d/q4fBwyJRN+wAQOTNfISMcL98MA5SVlTs+oXH5lQ3yjaReLz
vC0tTzlipTHWB8mls00uGr7gtI/8LCyHbQHgRVD1/GGhFZjACm1rNQaovK6oPu9V
i/9MZcHcjHrsvuR7IDG+U9N98BE0OD7irukb6i3JmeGBdAxj6kdwiFJCNm52FLXH
nDBleSrR9/T7JDNgKD866HyDyvkoCKu/GmfXHtrn3MzKLlmDnvrKIDIrmTfxTe0e
0n7PwHL+X6c9dQJokFHu9eqrb5jNAxI0SepD0k/MSnTequOdQlYxQi8JJ/Tsutbg
bqYTE+X1SCllUk5IIYAXLLBZBxSpZ6BOvu64CPryluABh79i1CwjMf6eUZUfTlBo
1xJ9A8ayj5DNgGvQsK97pLs7to2ZgSoEpEpkJ6ZCiupOVmHn/0DCg+K75A+hdm6l
F49AyRZkD/fE82Qa+JFQjYnLjWkVFPeadNOpkQ4/bRxxi6uZ/31g/yB1eU/YbZQp
DuBdcyoLZSfgG7HJutKBa1OyY1XR9PgKNT9ZT9Ab1j6mYkB6EKvvsie6KixKiNY2
MzSYGO2I5zHWkSf1n8OLfJiWitfd+Fs/Fx1WdzR7kBgbHY5gLxZkTFtEzYPGdDPl
XTRnYMYJxiF42OdF3srA+RzEFCn9FofONGTlfZedfcZhh+8ycLAlwQqxYZkPPcOG
TuWMFVzfqBAQrFYZyNVdzRRPSOGsP5+lSvP4eO6wBotdK6SgSnvCXDb0YHCacJKS
pDZ2b1lI6kKh2s1vfgMxLAKiuBJc4eHFq8+m/j2HM5M+kd1lukuL8EQnLAbpuRrS
uPtSAgrn9VyISREMXOFN/qyOGC48uz1Hl35OXd3FgGXaInLm2MyfEQM/3wENbprZ
IoJR2dHpTzXo3TpSJnMKKJPYCS+uYbadtFxUrVqsurZT3c8wYSDJwjoZ7FRmfLcF
vD+Ho2t97kZ8zQ0Y2ZdKuZyZgUGUlY9POYGzQn1cvfGbBKlCl73DFFzYh2FSNNDz
jNBDMCr6JGIZXzGJgINOghLB1gkon/rvZoH42GN3RpbqIUVliSNg0D+0qVtuD8my
LpxInW6FrJ6MPn+yXHL3fNdDPGO1OGMkZ0kWNZJ8nfYe/+J3cnRXtvNTiG1848tw
alLkdcrAFm54OAaHAgGwBjKEKW3IgHpCq7nknBzzjTB8Ja9qPtFSrSdZpfjkOrPP
Qc09qEkXa0SM1M1fVp4IueBD065Ae8Gut1M9JcYy9b6oYRCB+mx+VlG5USxr+KPp
/30Yf5Lq3Ht0SRlxHGRuInDpSTglM3ZpXSIbhBQ7/VkMtKakuFzDqSDcK3FrVD/Q
S3KKOqEWNB40JRqsdrlRyZd+RqqNIsYZBGoRDSSYB2qQjlg/pXVTI47/9wXmqNTd
wFpD7+ymcWQTWKkkfsjbHoMZaGJNren0oTw4z9IZxddbrHV9jdcaoDVIp8nDjWNF
j+BGq1kk+jKRYgp6ttg5cRY9sNIpqS3mFczKjy4yU30qONf3nIai7AcEt+ou8I1o
x37nt5ePP+qznLHarmSOdFtb7ddy6bx4lpewT38ir6FQIz5eew9Aly5S1AVpPX5Q
/o9u5nEWM1xgkYdvuixHHEM+tRDr4WWmpqslqP82c1cnCvOoZEFDyrkl1HCjVftW
48Z3OYVs2wQOOauM1ysy/RVr2wunB39iFoD0d4PQ8vsEWgeniEhqAsWgKCiDtFas
6DRuJLLi/xJMxzCk0dmUtSrSCaR6+KUy3DllAoENLHBWzYKbQhYCu26JhR0VTWtU
B4G/qtMU2/KUut6tznj1SxH6fpfguZ1Z5akQY97XOYVQPbmT5ZYOb2rH5ivFDTLg
NxRUfKZfQppzP7HmTSHoDH4LcZIhffR0Wy5xySQFmc+gnAGUy4O/tX+5bnH5KFfj
LM5DmgTEK+T6aVSzorRAeAI4lwo/8/fcYkuBYvr2xULvJRpxrDViLxcIcZzooLGn
xstOCsQEVOiVJ/yNx+J077yA8mR74AnHBdxeGc3pghUqVbAHFUQp1WeYdbzOT1OH
Xz42kAuji96Hpf2Z8GailqjQAi21na5rS40EgMDHO4fxiqX+JmX6V2r4pWGXmDN0
pfRt/S8UhA5txcErYHc13+NIBm2oR1Znam6psAnyKKE6Fs3bGbZzX93TubmOc9Kt
XvR6fhsxD3DiprmtnifzyNifWCcNYKSqPu3ZP6q7bQVrTwVn8x4zP4GL6p1jms6r
9tP7sgOihef5RIYZB615Gg7xkofnXaaYT5CPMCTh9TLwHsRPhvjYvd7VaINVbC1j
B9jiIjOwcDnqzQ1U557G3cQowEXjMwYEr0V/ZvHZOWQLO4TXxaSdk84KjYNcZ4B7
N8Ce6wbOv2GTctat4TEx0Bf/JhcceOyggQRffuVCXrs/Ke3lB63txKleC4jNlgOl
pY8Cj/YN6x1Y5Gzelfg//1T3kCmMnfUxFlviqvXa/SGG8jx63fJz/ltCiLxAfeVP
B3lGhOB/jtOqJLbLWVYEzX3GLQnQVcZxHC1/m67NMbjAA0K5kQvXwSgRAm/JtCsR
RAxeJjN4G1zRXM6CugjI2HCw32SK1nJPJ/6Y9SV4LtzP4timk3Fm6fljxEWGObNq
D1lAXvUd6gn8p5ebqQPpkn062dCYXO4qY8A1lhVMY45n0x6VMZvl8HvNYYqJBslW
DFHuMvUjtIg6+0uZMRNI8LPpsxuLehZE50OJqIDApKJbxoQmEmEU34oBOvPWvmmE
xsg6+CPaJ7a9c7CqxN8SgLXM5eF9u+hKa1geQpTgu+N5CRqdPveUXm9gPaKaHQxW
B5pR7SQ/xZCsyRQZK2ciZ2PMEo4qkS/Yz8rQdAE3qaxSGaLyjM+pOCTPFpZFhXD7
C3KNv4EzMk4udOA6WDkNdjvG7qn6Zg7cXee+twV5WTEwQCRnv74CsRrYTUGQRo1F
pjC5Nb9A3HbMw9sEI11+0dYPiIAnxowi0TS1g/LfbImmN3EePhG17/l9zhuelmo0
7kPAtLxa2Qd4Ul8uCkwCRq3za39BKm1dgM/NEP9rBFTbCwSM3STEhauN3SZoYA0H
Vu12nqkfDdVFKuICHqV3B5J+CQ6MKE3kyat/yJulqa8FryZGALjOXaWm56uAwJZq
heMp5nFZsmWG2bC9VreJyA2rA65/U7brnxSFMdoW0MI8anM/vn+XW9WvHKgu6+tg
PFIcX/9o1pNcWL4JjrQNHWC5rs3y4IBd/TAcBQ2egWUg2Doy1+yEd+3GBMHDG6HR
0uER0exlRG+hjp+YtFRmTHyaqSnPzvT2pTraeN+W0Q1AIffb7niRmIT0v/d67nux
TKN520vW7t3FQ5xA3hvylxtEpwcZqMyfrc3KeRzNbOWIo0BxF2xHC4mC81syo6NC
irIXQIuG9zO12mL9Q/33VpmE6YsBmM09a/pByWkaiUymqJsPpm42I9YW3pM7fkJY
ka4wS+E4KmGj3QKVfyyqkEsxJdwfpf6L+2SG6RJF5YgSg1IV3yDK+cjR2ELl4hxq
BwqQ17PTv9gjGKwOXP/4a1/rf7cttRkhiVEzOUoyoRo=
`pragma protect end_protected

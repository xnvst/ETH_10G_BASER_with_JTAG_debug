// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ZSgVcPkmF7p9woTtCkrI/y3xY/u+qvJQ+0XqDhpK1kqsPWof8fstJDZaui8J8m9VdJgM4wnoIpz+
0Ai7nMnlQf5Cy5/fZsDib3pWFz4RwkkgTWKvQoC2ePnnWYsB0Cdo4/Haq56lg5Sm3/KVj9A+npMR
7ugFb0zqPmI5DIn5xGyQU/YnMXlIg3B/EFv0RuzUbrgiMjT1PFk+y5uQDGgnfLakwFfH7B2jetR+
01f8CEtMb+U5PSHSyIGF1hg7RB3xk2AHUuk05PM/nVdWIVMriOf8hxiUoB9PQ5inB/PNAwUNWn7t
fYHwQDdJMdIZUon2hBeWLBUYXOOqI257JnuZbA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
8WjybXO9K2VxRIXUTsO7SL/wIV7HVOdaHrfBJZTuu5vtu/3GvTx2o8mBsVjOb6R3Zv8I+2IyAubE
xFEpGTLrZ7Iu+N+Vg2voHtRh1h3VSXwNYi4tHwAlKkbDPoQllEOJU7e67UpKJY0XuDuFv0yoTb1b
IAuA63zmrJJnVo/X0aLaO1YkFqjEBexB/EDtZHZYjdWFwbZvzpRfFpdhqH+qm6IWkYKcqudnu4cs
7ywghIrGeh2tVXMWRyI3/LUwh2Cuh04i7SuISLcWQxSaQ9pKufMR6S/JjnI22vqEQKtB9ysKpKa4
/XZPhkcBveCmnR/b9grR4VjdNDwQwTQSx0dU6QuTNY24H/QxFGX+WVM2p/M3Kac8Saab6y+4SooO
t+FPjdfUEg9nNQXF+yqe/ziM2S9q2Orq+QnE5n1skDcqF4JKwWKWbQJ6G+GAxtxqUPRwKBLUBYDI
M4FAi7DLXILusUIQZpBaA8uJtwkswcjX2cLuA98ygDaFR2onVj5HNBBdBg9WB0Ik0xfqkoKtAFKo
wnrb0QRpOz7Vyc0uPlGi/Jr8Sb1bqAWYHL+OYFGjNdbtAMeJyurhePjFUi9FRDdhG2FI0VjolPGQ
feq/Pxda3dKcDDa+WqvOgLgQeylx9nV6qbXz5W/Om1L9bTjCsvZoSe2Q3EoA5PPxfN5t3taYyveB
CBF4KLsDn073hy9Z+ZN21m/CzxWn8JDPIq6+2++VP1g5iETxTsck2QHaJmHnY/v9e5s9emfJHfG8
vDKS4831M/DVMpqur52IWx5RI03g7UjOW9JxFrP7qP4LY1wdAtrSznOdGgiHhESMS0wMYF96O+U5
T/sSSUDM3ZO//YquzPv0wK+yWlaxGxZ6z98G8sebp/UXbuAvQTjskrv1XEw8DMpQTgOny7v8hRFF
hJ0K5PPJ6bSMVqYGsJfJw+3xdjpOmxVnGLkUO0e7UpZ8uAJziUdfSZERyrQu/PlONIdjDZw+jLKO
DOAz3IJmEeNATVYYRKrBaApt2ENNy8vUwnQ25rSIRDb6liHYUoznQSZqLd7AOM80pli/X+tFjwzZ
OfiBBYmlfmt7terwu9KIZewrXyjK4xDdNoaTUGg4nuwfd5kk9F/MKN8n/nYJX0atefIuaA169CmC
D3bkMzvJTRHo4PlboZ/eANzYl6GKBZbtJAlKbjxIs4W5Gc7GarEwq5UiClIv/Hvwjig/vv3OHoyQ
hOfHRjgfN7Hznu/+5IuMxSt34dxlklyjlXK2W4T6crAOfDykI7QX15EnlKAdxn5bguEW6Lxrjddd
sE3afPj9VfkkEht2a+FscU/4QBe1fk+ke2T/yjAc9qGZnPjP0Uq23HlwT4sattYGpRZovuuanNLl
tmkbYAeKN0I4ql3aR6vV+WX32uMq+4YAiclZMua8VKRlDkaMLmugJOka/IhWRDZF1rXMlqLKC3xm
n2Zf0kRutCY+CVEf0htEws/L1hSHbcj2wEgyMFdy10WUhC64je3dCoGJumIUFrTFLGhD51gZpzzE
w6xSCD0FiB3bSafyxg+C6j3nN2BXidCkNpvgxweCGXNb94s4gWgT4fwUcLyiYn2n39+IX9fOoce1
Ed3peE6YheNYODf3hp88aGB1hA7vPKNIuuUWwd4TrvtR5XkaeOUY8wf0M+f34hIeK7iEzhiakO4d
FpvbA7KkDgvtmV7zFUxovcLG+f4WMsmIPY+8I9MkFHDv2+8bnrJDW81WWvzOEtx5oPBZCUpFkugO
yYDzZCY8DRjtZVr/5Im5HPjDwIMqL4HO06u/Y7Xn/8Tg+q2Qd9LX7V3LHtCERWjnfxsbep9T2TaA
UQrL5j2EaqM9DsZ0y/ONHxRuoWv27Vs6JovK9he53/J5Rp5NzJeUBY9jPDN1jiuOSPqLFrdyhRNa
7cpg0cGfiN5cuJxR/b3KCSSsMSYaJt5CEXq5CH9QshcVEfGs8eoY7MEDHy66Cq8+d9SOA8Nte0O3
uj4JDAfLgE9oykf9Ersghc0MwWWe2pkmcXiZoMRndUmVmRsfuc4joq1ae3af2DplA6+abnmZVGhY
cRqrFXYuwL/9Qfp090wBM9itTEsV4adNmNjq1D5mxQt78x5UnsgCvAv+ARTEwnyE1PtfFPZYZKWt
vsjutfYMcy9gizDvFpeRBdraQvoIyougPcVo/luE/LYNnxCP6qJ3jrSfNYvfy8mybyVy1QNsc/3J
sEc4+ZbtD+V85JyCQNp+/nUFYvGBqq2lnE02xSMFGjmWOMXp+KZn7vEFg9c+CVR9fMJSj4E43wD7
gMycN2jtcHvTJ0s6YUqZX+rQvktVkM/sgf3ZG+itHCsvP5kGnM/7lqxry3t4B7VtYoGs9lAhZoxc
irUFeqIBMEJ3ZFPiHbFUahDhe+kGrwhHt1xOh5G8cxDmYxgVW/hQ9HTwDyZD88pel7DTze34q6/Y
L4zlgHwr3F6OUpgzP8rFUW+0nt822czqigByEmtAQuHlKb0cmP5w67C2A1gaFOJlqS/l6htfawSp
K2b03PmLbQnwrl7S5uXXVh68+4LIBp6W2s6WahOA0//0KVGulhMGkMxWedGm1/8ajjArRV4gZ9+/
YU+gdH0M7J91Udpu6cWbpF8F0nr4eRSjDioeLagnyVr2uc2dpYXu+OSZokXgXks0VCHEs9ou3HHs
8bK36O3SM5K/lTI9PYtgx/GMy/prX39Cemx/uv4PhssXSBUmyMZf7jjGGRa4ZbsLf2e8guhHoTXY
y+Da+qRiaEBMc12y3EhXtloNnBjVZ7gZc/ZqUhEFY8raDjA5UPxT94c/XJa9zVEs+tRp3qv3aF9V
lq1ftrqNC8/mTAsLd4OKLSTzja45LZddrGpXM2HplfuIkvuxRCcRyXwRvd6CvCR0jx06n0jVmVgd
hIajKDXW4ZmzXy0mwYrE1C9xRMvwN+nhEqSbp58dwk+B6sqHEaB1Ubwq0ZcFSXEy5AGvJ77Zj9vY
th8bAEx0UEptkEl/+8lmDHGLgBnsjulnvH1qA4jhoy14M9BxoSfEGS5tlnf8v7PuWhgZmUBaz6ih
C5dGJ4Yb1fz1ya7u/2Vbe1xDKdLBptq6Q9iXhw/Wve6BXTIS0p5042q9TH6ZNcgJ2jPl5OUPDDWL
WOQNHeLLloWwD4idRNVHFYU5ehO0e2mTGnEVsu233G5ylTwqRxC4x5xQ0k5JjodP63FDw5aRtWlU
zFB908HwU2ts4nHDj3dAeBLgAcA4f5GXsP5IYXuivCq8yC66pM9PbCeHUYILUmqE96WgcLAXqlgx
Z1ccY+PyPi3X48a/pZ7TRP36mZ4aisVLVi412HKaAEtiHQ+uC/3tnwE66M/kEvUe6WBTrVBfFMtH
LxpAbtcFUSPTuy1tAj6BeXQ/6OZf5x7Va1anl07wZ1KTA89WKnoIhv93zK+mRXzyNF0T2mbHQZuX
SviZ2qlhX41jThQSPTGddQZb2V35yYsgZpJTxehib3HcdD+XnosOHQBLECKXaIHFoKtlbPGOn1z4
+HngguKTQM4TXAr8gaXWSKB2/BZANNzJ4T5SNlzQsvXN4vAfioWLEaBqrqfj/SFlVgHMVCND8rYP
R5gq8rxM6XdB1vy4UNWJNgQM5Iv8Mbniz27MLBv8dRTZsM8kQqpjNo2I94AtqNmpXY+rNzRXmepg
LsR1qS6YUsSP/umr957aupKSiMNjskUUyEDBcxfr7PvKWl5F/D5pbyxJXgAXWlHrQFYjPOe/z+AY
3VcqzyqTsSBFq4aU60zLGExfBMDVgGBxrfIc5ZrmvfkxjGrgRyPZlx7wCCEZCN7xcwL9RSkaVE+9
b4wSiywhKkZF5gV0CkJiIe5IK3dWmB49aT0ySA3hl4g9jC8zt/EbILfm/YevaUfKj1vPSFQuRq/L
GaUa0Dk5yPhuCw44TKmzGt2kP1cM/vSCLktkb3Qsj5rEPRuxb/hQL//Kte2NWOIxjn4mLM0xifLt
WSxjGJcbHPRaxF/dA3kJJBDIc5qHTyKpBbw50uXuXM7TsKZuYuqRoq1z8s1APYTlUybMKpo3UCkX
snZWyhfz3a42luqW8FC8LH7rI5wNHUhGIMyEV5i0QilEI3wiOr6nvzFmK2xf0CA0GXIC6tjEPsTx
9F+1gbFKTi5aWi3fkwdgdAOMTKcDvy0Wu6xgx30ICxgWuUdjEzXkbdFfQOhVINyGsMtSJck4MqBK
86+VM4kPJes2Ab6z7Wz8B0XZgNqg71oJ0RoiFaEQe/Y+RBAvwaoV0m9pxe5JaUSTTsdIi8RImzm8
dsIAgzWwx70hTDnxInQnqUB0W87yvq7k/3TGl9Znv7SGx6xYzWY0wfM/GKwlTUGTh5ySNuOFEja4
vGJcbKLV13SFL3IS/XJg1K0Em/jJC6EkOUVcYWBGwS3gR2nwCgQTuCbVzfmhIc3hfdEozPUXzWhq
uZiZj+F6f1WHI3ZW+xnJMWrlK1/jWUvrjjIPdYnKOSc977YVShTHGjIzZsGCTjUEAc7wwrilOMoX
y2maHfS992QtJhyzCe1e2gwtKzmsI/Jl/SJ1Ek2IVYq+SI4CHmuq6/60QkzTz9PU+lnbTDJJDq+F
/8A853DfeP7PjDONo+0/oMGCBO5iS6WN9Kz1qjaO7YhQD7SJtyIIYeEt1mMgwFVc650LQ3Ym61au
XreDRNLpsGFfJfDPGew+eQraXdB3zhazbkFACLVPtHlKg0xrJKQI6LEfLEa0BLDRxi0zGG4KudbL
/8XxpxZ26xzQtb9KOpKmsn5mF8C/XI6GT6F12Myvru58JxRoFT4WeZl9UX7ys5k6NG1FNVxK5+gc
nSrIXwLaTZgkjz3YUe9IE0aUpIZ/9tXpMhYa6b5SXFDJrJMwvAs8XGac0Z8b10IsqxX8m+uDkr3n
+p6bpNFiEfSyn/viP/1dJENb5uoscv7MPyUucQJZ3wF3AJcougBJaGObcgCVYkxvY+x7GaSbrzvp
qPZf00MI39f+uep0OKHJaj9/NNOcylwrodFs/u46BOlk4G26pogMKKoKLC47O2drNxH68exqUu4Q
UTw++j2NYaVL8XOMB74CHLdbdK6mq5Rq2dZDAVk8OnR1h4z5omcE+0aQIXtGHApNjlcgO6BO4pJM
ovGBNIm8+saonjF2IYvU4h/K4JNs609XG0Fv0nSTWnzU/Oqd+mKKOb1CKRJAxvvyYhIQouhmh87H
HcgzrGtsAmZcfG+DKH8T3Ppy6zJt4tB6w6pBO3UJwNUyK3mBsyTFdoCxwLoI2dJ82dskoptdHIfi
ijZuie98Hc78hdWm17uQecWqAPfENzK3mJUF9RQ3CCPs8HNNiydTTvtOg3l1nKW2SgHElNaI06NS
wDthptC3X11zve1KBuXp9BwyhplepShM+rcpqb8tvp/+cjyEatpaQBa0nIM9HeoqDs9KDlxc1oMN
+xo5N1lgp3DEiTa5Lv7t+QbC9LwB+gyUWOFXNJsOckKaQrLWCne+H01nsY2bNeeIyNpcU/IPZ/2q
nDQ1uNRkCR9PSk0TU/jxwxCXuBBjEfCqu4+m8w0DRdL59zLezvYrMYo8VR7yCWJHGBYDNH6nzopX
KzFdBhQuziz+UJ2ff077vcJ8gTulbCi/A1v6MXrLK9Dt1M9qwOVD9or/h32OQakYuF6Cidmt4vVz
ILuaVQJIX24s8IeQ2Gcqx9EGh9eXKbAsWEu3aTWNLqggKYegSXV3PIgHXFX5zG+xGxDI77bfrOGh
ryZhztpzhJX6ZHK7ulU84hGZOgbNL9ogoNVUAv8gDGJL2nEMREwLw665ZfPaJb9d5tyQVNv0x3ty
+fQrbVbpPZNl3r63E2WPc/clDwF0MW2SvS3MvJ6lta9Fl81bNReiaJMcW/uuR/DyGbsSCQzH/Ny1
o5UP1WsCsusWWwdLOziZuq3l4hv1yTRXAajxRHke+e5gHKpN40K7IfvJqjDZ1l24MFkySqKKwljM
UCMwhhLbxVfcmUPSXmO4/biynWQ/kKFK6F6nODGwKc/gWE0k7akb17R0mzgYaZP0MHMc1iLUdnmx
iVY2iW28DO9JLjH/HcK5D+wYeJbTPK0kUl2apBFQe4g/VkeJQZUxmeyW7ni7PzzRfUd5Swywme9G
mXt+YFpkJ8+S9auQ1YbIm2022lbp3WtvwWJW0BrmauyiT+NhZTWJhDDqIPolN6ZgU52KlIPT97wa
/czwIAEMmqGr4dV26AgitfYZSeyQh77qDSjDktHMuzpTtTTE/zsEXN1bwFCWg0S05CQczES5tfCM
NoSTf3zNBdreLJz5B/ts2KGx4C8lokZe1h/f+iKtoYRuPGTPsRln9dckLsM6RmHd/NrhZzuf7/U7
d/3z9cNssSz0u8LajT07ypr9dMzJhrAfFTZAzhpXkMGPVMHVAUKcnNLLaXsZO+fsd25ZgA3+3ehD
pu9RiW9oyUOGMkGFQuYtzBRIumuh/FQL/fSEHirQpQ0gEbOmTiDnyXYc24yZJA9TwJxby2xFejdd
knQRDNX4toNmLz7zhiR0E0bwRdTFJJu9TdyX4ewBt1KUX1wh1GQnIs0cnvsHQOOuWr0tHdT6049w
LZIlUDyCZlEIAqaK06TqStFHnFw9tdpkeMd4l71ktyxo0Vj3+3uBJMAzVK1slPgcSNNrAIgWqpMB
Sg==
`pragma protect end_protected

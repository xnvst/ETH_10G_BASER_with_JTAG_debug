// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:34 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MlJK/POaQEkPD0ZxSJVSJ29pL8rvTfflsSJ+85ku3Qk09+z/R8v3Uwq6YSbGgTwo
JsCIXU9F4nw13Q2W5q1QzlUWPJv7RisqczNqLLiyjVv3qfcawiiCUSYFOpf5vtys
e3wyPQXRBsma8xWBXIsVsN5HH5llR10vtBjIq4kF+bo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5168)
2EpFYq5qiBiEw0axrcymzyu8osZnc3LkXCHepHbpMBv8a7pfD0FIEauuxh12QZQO
lmYIkGyOCqePqCkGgqx0ffHq2vbCOCIPIQzQM56h/bFdIz2PizHjXM1IawmrH9ys
wiVFpTU8Fzhey7ELEFjA3i4NfbUUH2Zfzl0nZQcoZVxiy/Qoq/UAiPbwat/cBahp
uHAItCBTdmnufx7QEaHCGhIlFqOFR9BOwKDMgDnlfoQtuq+uYRG2a0hc0TUwtSQw
G0ICIA8/Lfb+gJUlg5yNFk+lzUShtRpje2dnRc375HZK6Bp6ejSxZlGiZ4PIdW1p
A/n5ESd7huMNxiGvweIebyJ9DLQHMJHClbIwHq1X22ItTrKrdZSSbR3twZmtCc/f
vhAfWltGlBiUlqZ6u7rDFXciT6ZT7Jc39ifYuIHBp54yFAtMIw5AUH3+LEJpErr5
q3dy1fcD9R0Ulp4/WUi/IKit0CL1zL2zbmpKBPETzansH25t54XDp4GoJXOVOZCW
NvPpWz56SWMJdV5c+t9s6KHqYVDmyyiPGzPgLm9nmVd0T1cik+yyLkhVBEKE0BU2
qcEJ75IWWPXrhkmwM1GbSUJloZbhKyCAbq7FZsIei3304N7H4On+BTjHDVFJiB5d
0w0u3hzfZB74qKpPgvHHyplXNxlyE8s1t/e02yy9085O1IDtgOMRW7sGobaJyQfy
ZgTsDz17o7iaZRh07dKeFHVnyAEpHuUu9HwOpx5a9tjRfkI3zOEmW+jSIsivFgKh
nQI2HHpulQqWgeEMRDg5Weg5jQzO/MKJ42FfS4n1tYCLb4bmaOfC1I2ZHrXT/LBA
RwdJDE7xF9205pkgQ0o7PusciQF0ia7T11UZt0yb0qjzJ91ZezxqECaG6pKUTvw/
OlKjNJTs8ust/YdAHju2zRr08QBc5CnBa7PqBGxQhwiT9qkgklLjgdKPq7B2ltA1
1ry+oKxV14SAwuCnYNTMiATcHYl69ezgBP1310NKn9QbLhxQfBpwsqLEgNOkyIEo
Ta15UmfFmglkhS8fRrPjkee4Z3FQq05DwUCVCtodN5hU6vvGJ9kyDg1aT55VrVVn
Dttux3uBJcr4yIeu/LmKJfLWDZk//GVVFklIQ6gWTOdQQ7GN9OYULXWA2Vb1ha8L
XvnI0UeT+RSdog3Zthg5huKIXl3ajA1ZfoIDv8If/eOj4SOCl22vMvsAvreAlU7V
cnVRuyatPXUJE3EU7p9I1Ri81XK0aDq2UKVmXECCG9Bj2x3OibDtdYL76Wen5XMI
fwJFUDAgSJ+udJP0vENhLC7aes9hrEsd7wZdYGJhAoIc0yIrRxOpXDaNZlh0Mn2H
DvrINs2qJjX2n6E8bAnNSMHYTBVDj5pc6XyL+Vr4gBE/1p9URyYRdqiFEQKwOAPx
L1p0+r4t7I0znJ7Od0MzV0EGp25kK/kwlGfBhUzz7BoDkWl1Qbmg8UASMFW3hlKb
fo5gpj3qpIgCUGsBQUbxsWh+KfCEjUQignkrS6KxfEANwws6+Rej0UvgO0N4poxL
PsrpKEe+vkdaGagITg0yF04QCC2hnprvXFgXypJIgbb2ALyo0kQ6TXXtNKZcUV/M
7FvK1aSTBFzS0is3kQKarmYBUoxv6Bo9WadNiE/ryuiYQbtDOeSv4cjEsmKTn467
N7SGZjHHPFKso5iYzDqPdq5jKPiLZl0U/O+IJk0BBG0CHMxx8by6es6YKS2k530q
ILcB8xoha2n1f8cFukxKs8zpzH0j/s68+jycsraP12Xak6Dmt4YLVCTdZmDZwFT9
PQatmXeBx9karoGZRSJzGAGG0XkcuE51wQjo8I3nvMjV6hN2T8/Ck1ETKG7AEyG2
ZisQ06kI1oJ52A8IYKYLKfEgLucF7bhcZrd2eoMfSkinN6gpFzzyW+ZbLFfi9R0z
MPJFyjC5PDXLVIu3qvPQPn/Xs0jxZV/dTDapI8+1oW34yVhS6IZIFP3I0ucnRoAQ
IvorYG/Y8UdCP21+7KIM9W2tCmWwfVToWgN3LIz/EO2S/VoW7n/iSpNvxMK2Cy6I
7uHAhGw9ZumegQk4Law/2iAKXL6AT/c+TDWgfVwFYLx542qqcZoh/6CXkxXrQMqa
JiVzRsxLGNGfIb8RuqTZayo6IRU5rrOBVBRK1lvmIJ6BBHBu4kvdLe21s7bqd2R2
bWWA2VFMhU96otuc1X+OODlsC6+PjVtHp3fxXbdNBHqLhMKmxRnSAszKtCmvothg
x80ZEXezDLnLsiEEWRsOH44kT3u6/96TO9YLyYrS62Aov9xmJQdtxDNrig8c5OCJ
k3W1NLwvYJAc+fhp6jZPXEi6fG1j4TeZRDpqLuz2bsqcLyOALwiYiPF9R4m1KViN
eYPXG3vfYT3YF9mmz408O9v7sbanNBpieXYDawEUiP74j7y2AUbOKBYk9zUU85KS
t7HJ3sqnjGRMJTAOb+YzsaoSa6/AEMu2UlPW4Zd9ySgx9MXrspZVWO9ooI+9jXKc
9RMwmgaQI5NDn7UpLthvK16L+MiQZJq7LTITFdmRrmoFIWIur+zoIeRI7qnLX44w
d96wcbfBeUZyhuZdojGXk6YLjQBXMeqrxKG3YMR1+02Oc+fmcCNm/IaZzw5Qht0a
mN/sjBu1fdFYEqoA3LanPdmi+1WT1EnsYgo6Y6eXiGGENd0qdBIeRMls7BHEGOg5
cIlmOIeRAh+DNhb/ESStti5BHoqVyzES5s7J7AskmHikEGr6TaPi1Cxby+KXhR9M
G8jPLTspcGCk8z9pu8fnl8x/orYdIt3UakiJ/WUGeoLZrktQdW8kK7Q0SYZdidpT
zyyxf89qgbLZ7ky1xxAIzLosUiFhnFW9qDhFcFQSRro4f+0erVVDJ3MiB0r1q8Hd
v/3VXbzX/kE3hP9pk1ubd0OsEOok9PYA0L/Tss5DYy3tWba+qOyxotwhKSJq8un6
Lfv5R2QPJiS9FmHPRh6AHWldt9Lf0qw34xu05uMz85p8GMszZPGVYi3b3m0YRWya
PjWEb/3liYF8KkEDY3M0MaQAVuJ6Xgim13i1+VIIxQWfouXSFondXX1rdIKJ/WU4
QR1nvTbUycAyH0m3Mn82BNZVx2XB6ZrCUjM1R7hsL6ofCpntQSIP1LR1ASlym5Ck
UZf7AxjbBg4enNZ7ZFhh1kma+IL9LLnyyG99lhuUc3Jqv2w8QDY928LlZ/Y9hdRB
lXlm5rf5HbdEsTeANc4rhlb48NXV7IjnAgm8Q0ZY8gvzfp4Ht2PwcwgRbLHLvYXF
rJW8IF659/HPWZIg54En3QTVkSPpjrbGRaq9MZ0aL2WHQsSRCr9KPLQ/TJpyRlia
kqVCue2tvlNOm7K1BTp3MTE80X99u0QKHJsNZAlE20OhCmw0jHopgNiTCVcFm7XJ
G0HNmE0OLDu8WfRqHEngAAvq7tROHh4m6GsW0u6olfvKC5+lu+Oj8ksG2P1qmJ1Q
hkGQrN+oWhwBMKu8sT8Z8AnZqf9xJY+v5zzYk+l9oHkSfWQ7xytokqrzgt2u/uaY
gSdLqJceCel9GgSwxImzbd2f+SCxQvgJVHCQ1Ndigkji1wqfKvj1Y3RaaSxvv2NN
E7BCusIB6xFYbFiI3N5q1eRSBJXUrGvTS8j6rNGDI+C8uF9D6CAUg6JsHjw95MKp
TC0buJgdO+x2cXq8QMMdjL94NPhlGLTM8dWyKzogbXdRTXYkIqVpALJri1F8ckUR
1VECf8IJopR4alYzTXrkqqBILY4sECRJhJ3BktCwCls4VhwfJMXZI38z3bi3WvLt
FPMXvFx+G77hypZo/MuQKe8VKXTSvrLoOdnPgW7rTjAPlO2UnQBruMbrXt83CLBB
C/2yYK36yUF1fGVPkcEULO1Nhu2hSYVh5bGkTRfM7v8T32E66rlELV69xNPNsgTH
xfgcwCjuSIKHUcQrbwJBW7U/gB4G5x6bni+KdaOSYrUYwVBOo3sh/7mmJjG+HeIV
PTrlDbF+jAamjB3Evn40ojwkwVtdHt7cTgN+FzrAPKPCcqWZkXqqb0E7stxtJ+ju
Dhhp2fclHLgI1O4Hp0eBuoZNazR4WO3kDCWtPhTdNqIQgmGCqFpfDj2y0lpN4kkb
U8ecf3cb0+RsOX5xFybbQ1Y21KATggtca/saIH6TEUctoRbNIirj710DKTyCkcZG
l/JH+ghfqnij0A7BZtyHaZ3fgWV8WkeL4IV7mbr8HoFtTBl99J/p8vWj0Y6SPO/P
EKZfvYPnt4dxKAwMx+H5vjbifFRoE9jdqUHfmNCWDhbVnkRAF5bj3HfQBQim8saJ
ips5hR0RthfkfkOs8gkPnWsxfdoIRlTi97aE8nqVdlqCMK+FAFXrwFbiaytWBiGZ
Tf1hNlAbF7ie1jg9YEbVEU9UppUDsN7VSALlfBXecwXsA78yglePh+GvjVTYkCi8
GG1oCJLzJUwqkQqKxDaGeTOc2ZmUZCrE3a7L+Y861I72rHcH1RiMZb0zc4oNKGxY
fII82mSAtw8sBgUjXCiBnosyXH36qtiWzsGwwIHT+EujCBMmXpY8Y3rDJsOa04Xe
pGSOMUcibcx3EK1BW6+eBUL6CLDqHCslDg/Gdt0vtY5syh+X4vwoLXJAAh4eRmCx
hGEaR4BofUPw8aKy4ft+6RbM//2OWrwgQsxt3oKCdtTAhxwplS5neCdVl9NwFBqH
DZa8t8KnqmEXliuElW0JdZCTMX/vz0jAHUJc0/A7OrbEhZPMSUor2g78xHsKkmj8
0xCz3UtlvJuQxfOAlH5C2EQRuIPCp5IQoDHhQJQK4FU7fFOB7MFTYEwkeHlMZPiP
Ah4+1msx8qEOuAbQLzCMBJ/hYwoAYO2XFFqrXu2xnyLVhGGN3gNyK64OXwgswRDP
S984iUw1RwHb4UX3bY4I/KH4vbJbom+eykft6OZnYT6ifMzr5OnpXyHx+09CcLBQ
tonmWulXfBwf+LVJe60Hjwg+C/KPHH0gtKjZeANMkMB+VX6dWRCJhf3PQN7syzwd
FTGVN3IAtrxkX2dqLWsvklCU5P1OvqYH4nX/1SkEjj3Ge3DN/ePkqelsUHsMRGP1
O/hbkQt6KqA0WzfeiWxJFgTJd6kHiBAfiyPmAV60spMAizwG5H9ZHGuKxrYjdr15
yonmqcybifxxen5pbABalFcPNjWnjG5HSQKjQcp4+3wqN1KGwQyO7ORQ2k3LH2aB
HDeRekZ+KsVQgiHkJTNqIv3vGjOeyeSfSvJTTqrbyvrlQEFySYCgnK+3Zv7KtnAc
ghoQ3kE3LJ5yNz4QkgvypG5b87I17gYBVIyLi/phIhdVQ72jCuFQos2E+AYrS+dp
+5hZ39oqDinxRXxsfUtLcuD25GeDC+ChIRRQWP7fQ3DGQAAGA11gkH2ZqxYEO2Cp
t5b5ZfY1VBMfMgWnLnJO9bhQWI9B0r9iZNElgwRqCSpAuIWwYM7Oz28Juf//vLRp
zP0Yipy0dN2S/W3XkZ+QuwcdGzKhxw2XHtlZILak+koqLrtqkMWHQuq9j7K6dJBQ
0sc3JxTGO2TP85/DvHHNeniruHiZa4ZdxEGePX+L8Xk1m0bcTtExTm9Ait+qhj3r
Vk2Pn8nvj3bVwKerdRyeJLVnO6ShrjxKphzM0Z4Lj56n9sg0eUIHUPI6lmfQoCUp
3Hc+cqgVDovyZd8HgL0OWU2Zr2wGK7zM5XhUj478A6Wawl1gBmQIT89UOfEfywXn
K+xTbHlaAAo5iSR3R3ZjAXLax54PbRlKCOaYKw0IQPXsa6ndjBlvsJGBZOeVjrcB
VDn869TKU8AGQpU7zJGZdkccgitq9VfROcbDKzZVV6wAZyVJ80TUcIcT1oHhAt9+
FxwkzbpRR0VlU6lv9bnVpp8SlM8Sn750a4ScOFapfop/orCSW6gry9ZAhNIWG5Bl
AW3N1norFsbM2bHB52gFU9ZU+790csP0M/HPnkbtVap+TYXAaIZYe7svFLXcmKLZ
I4F7ZGXoJ8VLxi3XbdW7GRnjOf6yCOaV05AnfIjvT1BIC+DMNNy2y9rglu0aa9Vf
l9j55NO2aUIIsXAK3BAsHBvSK17XAuzVIfJFaHI63zdEnOq7fnKPXq0Do0SKIafM
tf4sMddR9lUBeLNf6meIIxrnH0SlxE/E/EqQ7F3itQ0i8NnTuBa9GjGFWP6l1duI
eHG3cRshIjq78zKYzClJdk5UceLkMdOiYazxxR8yxlM3ekqglEJcWWdN7BZNe5Z0
G2MPAWJpzszCTe5NgkinUQOUwAHtgfBngxhL6KuOLEow+VjvMRBE9zIoC1H4a/2+
/wUy0EWz7/t7dyJCi+vLIRK7KurDwm6v1z8VSmBCtqJfxdSjxLXlgSK301BFl5DU
f/V//GGBPU3s7UTHEtlbLgoZ3DV6rlNmIIz7anqjlSUPDNgl1nSYt7BDhhX50VTX
hzyBwpx3wq8etr5sJriaI9DONoL9E2kJs0ZXoFQrIed5XC5ltVdjSowtaphKGsa5
PD6jkqDzSj5he/DWFlD+i8HPI5YgHSXXbTBem3MC8EBLhDIbYdM7OmXPLCDFK621
8UBF6DqaHQ0mtVQor6HYGgtTxk/o/RbE3bX9llpGcEpTLhnvPctjlRrw4Wvma9lp
tBGom9VwnihsLqfSn2RmGQfx/P+PkwL2IfRNIrPT8scLpjVRAM/dEevbofUfZ44F
4sH2PwOq+BGghGpEMcPNlNfZLlt+U+8KJ8Z4H87q9p/yn8uA7dKxSnd/2+vL+IuD
cn2/087CcdSz7yn4Qhtw1N5IP0trqHkAsnH52K7qL46GYeqoMZTQgSfgkuEZWhw4
552un2FKXhZ3XbrqYiEGrVyLx5mzJytRvqvJgHbjmuLsPQeC4sHnblWQ6gmkzTeC
LxUHd8puCLfxHOpcmnIEWa+QN+EN2mwA69mqzg4B3yQ=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:42 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BT9jE5elqFJuuh9Ft9o0Sd5w/P6J8aPI05VvIimK+zjwhl4jtHNLyGYJnzXl5xjP
Y2TzNq/evT2A7zS2OggTUByyWcbgvz4V6IEkhAB12Iu4oiXsUSDL78hUIe88/qkV
NgeX/8rXdlQPiTYIk4CV91jTuSNmndEFKInMlI7lfVI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3168)
gi0KJOZC6oqLylXIPcmSUY/6nrnrhBFy7C+OxmmVFADQ642ofwCD9lSWQ8FKc2Ld
+6ZCurIJqhDdNges+Rc9HVySr7AGtLltkcrVLV2yuz22u2vEEH6CU9gXroPmYEKI
VOQgWxoX2dRBQB8WxqO+uL5IK/8dLjgU+ah3kG4M+jj7SSqVn50J1hPiH98uAAxr
thksKSgJQr+L3MVQ0BMAUOA2PnTa1gyORM8LA1tzzp4EHj7ooDrbXCFpipMo4u2O
9t7Kdfux7b7Tq/6K/KJ3NROzzY2zneifm0PwHIoKIPzbvkASE460d31gvr6zFZYr
xJ45Y7uFrlMc03chgPnjIOBNllWTP5qSXm0tMxXaZdQCzXZ78ecFn9FdsX0LTzKX
+BT2HoEWOX7Q4VbZKGfFm+w+8/yG7aFCwnnOKCTqSu1Lxx1FtPD6TwvbR5hmp9P2
6pbjuDzi8yYlPk9EMUfmOB3sDTDVMPlPzN/k8L7nPNIQ5OCl7g7rVwuoueXi39Wp
o9MxKq01gsyaJT7zRVgWIz7+Z6SmflVBp76PBCRogefse+mH6NObtEaug3Z8Ii+v
pp2LrXn5oluvqC6iCzyNV+JY/+2wbx53xNazJg8nthiXpAkeNS3dyGoblsvUn+Wo
quXcDs2HCQ6lnoLjGOc4aIzdKtPZOz+YfF0nNxzfOVaXm2I3lu9UnGUU4QptS1cQ
i//i0mdvh377khBVDP5pwSSy48tPkswdJ04XAaXjV9WxtSiTcdcThXc+RSYT3KnP
4095YFpTtg7A0ZXW7NjxkjQxEDaudeb3UcBYr1VT1y1FQQ6xfZvU74OlOXci99oB
/xPMmrp5wwVRCU5+AFTBNnu3NyB5Hnx/LXg4v6XTJZ3Y4G9se2YeffGShFSD1H4K
prxd5gY33TpRcg/IMTyUc92kaqneH41DNvrtu5jPSozIPCNkKj06CgN+NCsUuzNA
bgWUZx3tNN7Kvfi64o7/jiIlNlDidrKxWVwPwKUNs4uNN4x/a7YRQChhjaRtOb29
zBfKpXC11hkhZMeMAbsTGABQeyACyHwWgt6tcJXyZFgqm9+3fVxXRO0e6ZQhWZgf
3BDpIdKx2B2mhdNkyIMoqoNRHOrx+UlRVOuJVrZZBnh5b9SgaQ2woGiYeZFr78GN
tt/rmiYSZwVALG5zIyYomtLcAoWA27qim/PTLt7QEV4i+hMmDG7dVrrBCPU9t6Bc
WRRhogNFw3RFRnNpquvOgMj2OQRdDp9byLtoUMjlXgfB+///zP88yeWNEQ6guSTv
xDRU9/DwQEIFCLmnhHD0M0LWZf7bK+QyFU9+rALnEkQxsiUJABe/oQ0ZBA4tMBol
vaAWdfGw4xd0XvjXbYvdtJoJ21IBJFwDfSnRvf4uqMN/XXzcVrx/TElclTol98Pb
pp1TKKVnThoLw7mtWFih+bLxPtcfl11ESAbwq50RT5AelOJxgI4ZucOnbLoM8AzV
/B0xOk92SuAFEJGSnJvSzulwPUF5llyHJMLwyAJ3kn0AcL9t0aMQcTZaOt5eh16g
4uaMdhpIrmOjfGF48vaVJ8Pr5OgCcin780ytlYQ2OE3Nw6MjZm3AsYLv5zXGMisZ
3BjRMuatK5+pLMd0dCzzwvP5icqIxNfThazJYcs4bADwQQnAZdNullK76YLlDIRk
EsbIB9PqpGlnt0cBu4Rbjd7jhfW+B5l/ffM4iVzPla233fmo+xwKntcilG9aFZdW
9phu7ggSYF+xRb5OJTOX5JYd9S+oRLwznG67RWFGKRfrPRt4QLx/hvGNLvnA7pvO
Z0aDu0Y25Vc5IBzIgPat5TNdkzxLGNh/w8e/WyIpGXU+eQL7/BPzxSiHIMiwkM+k
72IAsS29F40VN4FDf3e0aJLAWlyfWEZ5uNPaUrMZPSm+HEGBnQUjdeq+mNbC8LRY
WRMKwou1gKtEwo5Bqxs2NbLdPNPXkdh8WugaeNM0CWblLmJutmzKDQCM8h6YOaUH
ldIpAgyhXMbWZkN1Lpj+cnW6JWKBoaGjICGe5ek0thMgxvkrWVJWnVlxN2DcLj/O
aZaGWpfEU7hNUTDRRthrSizP8CA3Alnp2rdH9wm1GWb1J0Ds0ESh5dTjF4hbWIwF
MZGNbFjt88AtisngPzfg4p058vcj7xKl0XV4j1UpShd7erLvyMGx7PxOvZzZeKJV
1xb/XcK+IyES0o3tee7CICqebhdJInYad8YRWLQAiqB6B6Kfd+LEGTSLAhfNGIUG
tgTbdSpqQkhXdzScWXcNeOCJKapqtp1M0lVCIZAtjkjDYM+xzSTRKwb4ZPZ8QY6t
rAsYBbKQgAJzuVJvs8jZmKFujUHM1zkU1j1M4S7G4OiU5kmIq+bOEcSn2kLGs0qS
37jfpxP8rD9HbgY6M1VeZTZILQPmn3xKNRHQaXz2oN0WWFs4y7eyLiaNS3HOHiV9
gjihVGOoGlkUUziFjC9yERcB/uvV+qmT3Hn1l6P7+eXYnSZC4NEkJ9TddHCYBqY/
bV5wCg3BM3GeYz5R9dmjYZ6JqsMcwwDZxNDINzQj0UnpiIa24HYvE+H1NPBdGHuh
FyAmrbnbQFSgMi0u5cY510Qdhp3U1BsfsoxCKq3q91xE8FiqB1Vtyl+xjcBYeZpJ
wic798ihu7+Hk5ZBaWJg3zncu9uGCnPDc4DuoN+uz/p4u/msOBjBhl8MXIjEwn3n
mr6BS7R3YRzDVI2/hRYOGDr/4FmMLWBBzeeihrFAYZpD4h/Yrv3Arsd4kRlMYLUl
UcDkCiKj+kEmm1A6Qb7Ys73WJ53Es0HmzqxX0UmIS096TDhEF/Vsnym+HcZ/WAR3
Ny11uXYn1LcYjpTuHpcYFW+rTYdYXevYJfKhxuPNl5VIMlJKT8UbYjYEK9KOUpZy
jWj8fSEDEIcAlqCn0FyPxlOF0hxnaEXq+3N3Jp6WUwH4735KKEdRGDKhPpy4w4/D
4aQ0MVrkptN8StmjCcb+w6w80khsW4hEafRW6OlJVRuowxSUEOhc+lDqCiWHz/oG
ubAlLnMCWrGjL1V76Jj2BGx/7Rqxer1n5s3k70jVRv5iRCMnmA+ufOyJ+eX8w9+i
GEMDZqTXe3mYUlpsfAw7cy0s97jqnzF8UbebBiQ7xLcK2OCDkFwUt7Y0tYle1Wrc
5fz+Wjz99NKqaDJSgs0dMQAzoa7UkTU89qk3qAHGm+YYWQHBwzNnVsNNU33nPtrj
Z7tOVLY3ZE5ickarIChloXP6bapyDH/tYEOFYSVb7WXJX1bsoEYuTZnOaZhLqWOa
fEwpqdkirgyLYxpLlsRv9oRkRO/7rPRSLCVK2L2lImf1EEBZeTDRiLavXis8sgqt
9Dy4/IRNaw/Gus9t8hdmrtH3A5KH65+6ETg0IAeUgLqcyL+EoZWdzyGOFY49f0h8
lz9cnQ1ZCrEzNNPf5ONPDXxr8RVMJwMwsZ3PQP0t1BrKLVseXGNmMPKEh8qY93cp
nuODVcpczL+uyIT5bTcswB5ZCNKJXDej/+kdxTAcoyT99dEd363gA6wv93OGgFzK
TNbxxjqR2lNGclSeHUmMr7+X/cuuu1N3svbDRdpjFC0+nqEEFzeSRcDtMColPhPS
3GnvCyAa9spxJ9/fgiTHtkEUeId1T6k2cKRzPq/svvT6oYrETfWcywRBRw/iGG8T
nie7qjDIh5EpE5WWyQfwIhiV5c05ruu6aTgX4fSqDhO6p+fqllgudh6DWO6r5sG/
fvzMPIeOokD17pLOLqEmkszD1oaMTaYlh1N/s9mbhgwXsrMematSYC1OFaA0tGT4
qlJckwAIV2xM5dAsNawPe1SZq39smS2iAVn0kT98mMNyrUHFsZn5V215IfquLAUV
5t4vgbuqgsb95Xv7e+4szGVifpdf/UjQby1745af4c34IZ5g4TYk7pPR7Icz6hOe
RclZ/g0tIPzzvwL8ncvkbP+Vw9mQPJTM2l+QXpKoAQV6Fh9jYxkMx5yo0hierM3s
MBhrUT7gNa9r3LKxD7FYng9rwU5cvOdIJ2JgCd7/IVAuSUPKljiTt09TBGvJN14V
8gs9l26URT53LQswZEmhdDqlOj9ULLI800paI63BmTn/FFhi4afi+x3/M0EHBkSa
Bv3gi72sQcf6kW8pMOjmAZiPEszfZknc1sYfwCAfCZTo+vPagY1hlny50sPbzL8x
qJEavFFSvtdl55Me5uLnbLeIavrg6wpO65DhL1QSCaFnuevYGxF4D89IHYupvaiC
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:30 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F2QS3/As1Q2JI8Om4OatXPhr/lkOhp5+H8XazkvwuLZBlYtwGUuMXOIrrf1vTTIA
BTNJXp4VqnAdKcwDzYjpR5CkI8HnXaehPtlRxQaeczjyYcrtF1P2I6BKJ8LbL13Z
R4YQNENaG5T98KtSNDVR7smDuXCdIUNONQpUgYFj5Ds=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125600)
7Q5l4SIKxMjKzx3krQMoVZeFITLsp0VuhM4pYSFCDw0CxRJs2Qz8hr9E6qQ4F506
DtLVZ0T9LACnamSct1kuNOZJwBpKOg/PcH8t4NDOU3XDrg1N4ZIz/vPcAYoVsmKh
6CjWjZwlXHIuP4SEYwhvAa/ShI2BHGEp9oBD4yqFIowp0dd9XtbhOgGuipiwRCOP
+z4IqFcme5P0R/ZCFdkcyNX7bNc6G8s83F+eipqRNH9skgO4ApmbcX1fyI4P9rPN
g13OqegPGNip807a6yR1U0EWVqlCPIbMcZ85WXTC9gIX02TBVhykJ+tfvfiabTRC
qSgjFfL7ZRjSFcWTR7QJPc+k5GI4w6RJ7IqGbU4NKSoWquoqNEx2UEcgYZs4p1tj
GguTChy3+XDqlGpp8LqcmY5R7rxAAf9I475n8DF1i8B+g9dnu8xaKAFUimUj/19J
fvXpmbZ0xpSaUyLrNab1kxbsaPMHsA/nl8tZUDXWwo2P4AE4iURfWMK5F1GHvhNd
zAnaDM0buMOBzaStmjB7dDhWlCo4way+D0gNze7wKmDKXejml5Qx/3HXS+NVhfP5
xJfSZvAyhWf3FJ6zNVhOldjJym8iebn8yUt6itOkpIyZkMkzkzT56FaXjz10vyzD
B2R9hYrUqNwqWg644SENybse1X6yldI85MBvNfOgYsfhTIE4vb6dwBBl097+0/V5
sfxaPDZCu8BGcTCFHpHJ2DaJ1hxwUNkHVQfgGOatJifBSSxO9PDYgZIXawn/rZZt
wYT8phokVkCKiD3xbPEondslUrjs9AIjXMLxg4hmwIXzS1t/ZRtatIangCfO2oes
xU+Re9oJIQwPyqwYAr2wcHY667nSgki90QVFYt3qCN4qolv8C6aIXTKH/z40TTOw
GHR2g8jk8f6BTGEK6ObQLEEpOX5u2edJr6IJj/U2wt13u2YP+2EW4DwWmt7kCRgH
vqGDhRpImSi/m4+rHyWeWFm3kxvFVHT5+rtfhFAfjvMfxTvdBK+5vjljvpeT446o
g9sOcM4tT5KE3FHcjNq6oHTMRbfj5TwdLZf9GY8hK6SOGvG6nRZ17YinuMkwAUji
6Jy/RwCYT1Uh5KdXwz/Di0YyiXzF9qLfd3oPMwuW3nTCceUMa1tIsKEHmI3YN7NT
MBt0acDnt/uAbbHkJlYMPCFJHLNsLepO/USJpU/Ljvca+rt8TkBqKAefQpnF+398
Zl0CuXECMfDyXl7StXjT7pSVzRAFeGpquXJC1yX27XM0TheEVpAt+qm2G+sogguD
hlTDDSTonSYMEWkJl9c8Rnv6l6c85VCW0YrHplQxaHlXQrwvIc+9tAoqVtBECfni
FlbgYvR6cgZBkyVZnYWZL9eYpBsaHjnC/INiBsyGSsst4FOIlo1jAFxfbhdzivTa
kw1FG8pqhFQBR/yi3uMS99IV5qdmEDZtuzRc0j1rbtaKAwKn3gyssmDvvNKnY5en
gAG5jLuWpDUMAzRuRUrgEWiylbWCA/Au6hirrfuiUu3oWhF9vg0nKBRuN2jEIId4
uUvSfTGPe1ZFy590AL1pSUx+Aqn+imnQ77qkxUc8vjNciPWMKmTfXEw6GN4klBiy
S159eNp1lfZ9eIpCc3oqMtqP59xUTBpnuzSkqx3egbZFKpve2fbMghwc6CSv0NNv
NuO14t+mVxoVnHQByKzhrFse/uf5TpLGThOSRIcrL1GD/6xbBIwtbNL4nMZwB4Ke
bJ96HgWoJCbxzJvj7YbKrZSAuS+/5u/T4EJyIn4UmZ+9XyFDLpxaCdL05e+f/YY8
H7to/waCIDp8G3jXCFiTpU7a57sAv3CQhwNAZZgP7jisl/gVPd92FdlvrDyqQwUu
hhX/ovVzGjQH633LruHrV5h9EdgDFOBrIp2nnVRD2VpF7q5bRhUViW3Sk+Kf++Ay
V4pZ1kprL2vq4wi8EXhOsjQdSg0cxN5ugoD0ObcQjvsyZP8pQVbsBigq9UTOA+Bp
IAqf1RsEm59zKoyZaOc5CX90izA9YBkmhsywto8Un1sqkWq29fnThjGdYkLeby+z
vSF/9K9mN7SJsGfaI+j4UqGEF500yDNDJX6+C+gIHc6cSKLEvjWoaAcb8UO4Kg6J
4MGia9TeUkAvAowIO2EMOiER6DGSgAmJb75Xo2z7cjVESmA7ZaDr89tV4UVAM/It
1ulyVd5l+vcI2OnCkme7ICgSvkNTSfqo5p/wI0crtZguI0X8qfH30/Y7/XEbq/Lg
3nJkHspe5E1rUpYes4sg5X2K9kZMn+FyMBJ7+MIljpr24cI9FGEkplL0M6Tj3+8K
NuJ1u093qcsg9mTjYAc18tFdqhoX9EPw0CqYjGzUCKVWMh47sf/fg5fE7JIXRh3i
AJ8aDnrUnb6wa/ELpg3ZApThYlb2SxVPK8izcElsnPFP7HfEU3ELvkI6Xmz8hsWK
9NJO+bZxP2HVE7a50+c57z4sIe52nNQmMCKyCnLUOCjiRXgyLqQSWuwsHkGsWQlf
2rZ8CM9GfWeSJo6FldxTUNIe16HJvfn7ZY3IWs3TrhfPe6QMMkKgXrD7XucEW4j4
Dyy0sJ47/MP0qRxDYxOwWh5tgqHU1M0vi+r51Da7lqVKxqsCX5nSmiCsIVEw6cdM
XDOypzCIhNfWO+8xTpp+gaMBogkrOfqB6GfdRB6QIZnO9yt7SII5qxWve8DRT3z1
bMBor668lwcCN7cx1nRjBwXEWnstRGoeSya78hKDqD5vuXvTP2EX7Liv68AZPRfK
0e/ApS5tDfB54yipSSWDzZuy2ZucxC0FXaroKFWBKN+wS+WGr4nmCs4M3lkNSPNp
15OZDaQsOZ3SONjXdMS7QLeY3+F5SxsG3kymgDvYvnqswIfnzMNVxeV6bpmOWOhe
WRM46HwZKQUq44XZ7Jgv+DEQow676sY+6Xzr9yosEwM1y9ncMui8PnihjaoHXAkB
ncWbrQCuJBsT8/IsDSpvoE2nMuexkHjBCBcXYWDw/phAtFeNXA4LDCmG/wDiWgXe
D6KLlY4pRGLo0nllkLJzlvPYA1cw0k1mBeOnRprD+H/E2lfIOFh39gbFsr4EgJtL
VdzbcUZJxiMvwYiaj5ab6kVG/2clB6Q7d+xocZm1zO979N3I7PcdSfm3cpsw6MRN
cD1zfq5qTeodseTN8wOoam+Mt9dPLP9PnLhwz3If5GfFdW/305H8kdZQrsecZmgH
T06Z2FnqwsxBdoxlzIviFVBaCQMmx5rYNjH2O2qJQJvg0X+4GYnqnMVmv30vjHsG
iukv06A+zq5EnzLl/Krs4YSrxDSo7Rbv5mq0bMKobRZiZK8bJGmqRoo7rl6WftHN
NhUYzdBert2Q4jhip0p5ATOAhAl367wNcdauAHv/6n4gdNxQCA0OxxVWeWpg8ta1
iK3Ly4fQHkhLpS5Y/ubabDtNOEl9WtYdKSuS9TciKPrRCVzAbkGs6X1UynbimcSK
eIyEwpcrIWKOKKxvuJQALzVge6IUOjZSbyBXFMQWyuYKKa2vK+5OXhz3DzKQorR4
hPxIwg77maIXrNHwGOE/WaR3CD7GlCHVAGZuaAk0jAgl2hPTI17SipJLG4sfXonF
feHk7V8UGGLHaedBr1Y9QkK08EqHzD7s+dREV9Xafh/5D+uXtUupNSZhwIBZMG65
+YCqmESy56SvC3WjI53iwqJ1wGbBEbpu47lze4tp8b6+mTiT8eJ47FXbmBsBpJfC
tLUI//ctX7VlRUvgyl0SVBdF8m22JOUqT/9ETXoay5Gg/LSD02yNyco02OTsFFxi
QH5tvRjYEEeUhJFI03FaiOIcBv4bSsaEW/LsmMc0ETU+0Ra1OMYuLN9M0ggXgaRP
bmlUbiFClAAcOS+L2ur7w+uMHlxFLlknrX0l6b4ufQQ87zZBS1MIB1t+krEgv7CL
NboKQAl00us00fMvawBWWm0H2Cza+LP3da0ShYAwko/IbWyA5SU9y2c5//whA4EU
QZ9UXnjObvKIsTP2ugsMqVOcm2HUPHZvk1NjUY8Vxw3z4ZoBZns5HN2yWTB8yhUv
j/h6b1rK1r8maYbQzDIr/XFlNiMdkcEDvevkxg1AmQxztZbA53N49HVoMVggYjy7
1/epP74I0bAgfe5uWuXBZB38q5KzAcMjlF3vLvMvX+1oqWztpWxwgzQVunQwE86K
8AzR7puDPJZ/FSDqgQ1DNpubl3ZHsVWP0ndgqKreYoc2NQ+zvQu8PJmqk35zf3Eb
cbidLH32jDjPIqTrxGLyAXqxPLMQImsgYQTdgB7e0/BOJc0R2y+CvE3OV7fvRJy/
njHHUq6ZLnk8g0/qsx3Ws1eARyCn7orIEGgu+8EIpb7hSuXru6ugT8UNG16ngo90
IkBS9J9MnHcgPAX5T6iJiPF93v7bmeMLer/sgCMIHIq6h3MWW8VH3ondJGp9pcbE
CqcVyHsWUxqsiczQk9v1Eh+ez2zHVrc+Fzse98rSAs8xyA90ufPsgxK6dhLIk+VL
AJ8hFQ61jfk4Xhx1rEh09O8aLeT0vMu0exWcx4/K0/Y220svc0bvkhmoGIfOBBnx
qLq3NlOe3cKSAd0hJv47wQzjtAy80+KGtp4EGpHgVogGCG9wIpK+J8skb1QKB2VX
DsMA1pdn+239qKwn3sAMeIG2Z2FcBUGgrkxbnm91IAZYtGLufApo8GT68rw3FEvr
Pmnbnyqh+3Iugv+fXxOjuTD6j8H4up4IU1jHEdi5IkxKkcy/CxZodqYJ3Rh2eyNQ
P/2148sbgZjLX58o5GC5KqCAceRLEOCIIXO+2jn9zMrth81aiZn2ZdMDjrpxo7Kx
yenoo7MjUDW/PWSH1LVZP6GQ/C0rpNSRL6/jRnYwvNNoPNFa3dOEIetjXmdyxTVS
hHqnCZin3SwUdQ30dAr7neyjmaKoBBxNmXk2vPeZE3sNzTLK3A4ZwZAc5KEwRb8E
LApa7zNTAI9lwNkSd57d4Q5RjpEDGOy6SaAgC11OIms1+wvVj0em+ezeemVJI1Gz
tYW8aTbQszVAEonZfqlF2z5Le7WaK89bttG0fuya2UKgjucQy6r+VJd6DU8GdA0Q
hCp5OB1Jqt/rUS1Kv8/4DSiP5lpMbEGYJ26sBp0PVqXGZ/s3w1V005Fcl1L7ygbp
Xwz+kOWPzLPkBCVA57hsCUnCdIfj7Evqqeeso4aRKtYUSofGaBop/DiheRK0Lfh6
/y1jhpjzfh/mVk95iOLxcAGSpsPY1d0b7b6kXg0v0g8HcoJkJL2PyZ+Pfdwfbd6d
vdZp0hVC+TQMhL8YIpuv4Rdo5VMEEyyLDBYTUTAm3xbfO2pHdoJ7H8id65iji5Ab
JEF32NodYWVQTYqGolGmP2ciS3xlPAnCZUb7CIaE5B9HVcxP78RZvBG8+UtwH/Lf
RhKaPje3wZ8ekLlrTwx4/CMUQWy3w29kvy9wsR2aBf0Fy+z+qeSIX8KF8wI5pt70
+JLoDyuuggh5mzK88RMMjbzCjWkATY/Ew3aHz648yf9dr0/j3W5f7MO6T/cGN2cm
N5r6gxVN4fSvMt/FgX6lfuY9B+yRedJUAb1A/gq/LFG/U8pYbw5JpegyLxP3VXRi
ZBOXpWu0t9fs7uppToXnC6F8ROnxNibgNxdcY7+QT8eu9kAtOxjEVJeKcc37xrin
9lOKHf99nx96xtmAOhhsOouX1gmxtD1u4gJ+K0vKKLzKId8rrkzuI0eSoq2Z5Ftm
v6ABPhzWH8PzhsE8ZrbhBO6DheRstRiSWNg0KmC9WRItlQAy6yECG5ur7pAgJIK1
JN1zANvAIu4wurQIDQk9RaODyOSrLDdhVuX4QoFx6MfWLdQmfRSzPzD6KfmyHu7c
PCgmirIJZuSNxNpUuf3BYBpHNeaTjEZiDdXZdgH01IVyRTswfZKRTVA0RVt2tDmm
1W0f6Sle/Leczfo1OqRqPkeGcuv3x9OdyVRGhMKGQ//8eUqEkI6ls0NjKfcwRKNY
bmrFo3zvPKTRJ4EZ25zYi2G/7KRzxpbn4590nsqmMUFA55V+Q6+cOHD+08WQSAYi
+YOK1+AHjP+0Tg/EGV6GvYLIWpM+lRiysNvepFjvlckAJqWNWaOBXtfDVTnNHRWU
Lghb3NFi8TPWTs4qPQC3DGTMFA53E4VN1eaeaz9fZy1hTY1+8euj0uirjsYXsYEx
+bpS8cahb19mIxxAgOBSc0ejLuV3Ed4oIQRV1/FljW6dkqQl5YlG6nXpcT5JCOdp
XIwMRn3K2u8OE8SG91DqTewCOH1VlfiJSSzP9pAYQ/45aXAO+XZI1RBUrgj+ia5i
BCtABfbr5qe38VaIpS/AGGVJPCcEA9wOB3xST1oEgGQoELRJP2U1QiNRGbvTHDov
rgPnw84yXspKeNtn27kIZrIbvVGxwv8TGrQaW+En8jRMfSuaNQhuTuOOtNbB6n2K
UkDzo0zySNsPLJeQVLCII3eLWyoagwL446jiJx2P3YRdv2GZakGuXkAnjgbeAdZF
FO7cwxdtXDHl2dXOJr0WJ/oVDcP3g2Jr1xp2EsPoTZJDD/DdD81yV/yfIIHvd2Sg
gjLvVJa/pCHX4aQpIjca9f8q2Tf9QVLbfge+6zxAHD0nFNZAC+WT5kTPUGwrrsVD
b6TZEnN+RdopilN271N87Q3i/wBvFtKZY/LV3p0EwMEtkJmwEbN5D1G89cYk6XoM
wCwWwhnpZzA4YiPPKyXIbBZzoAiuI6/+AIKBEZCcQkuhAw09kjK1C0NTd24BFFF9
UTYx9Yz2CL+WwAtqfGYmMX040qDBxo/oy9cx8N6jsmnECm7NKtAyZ6pRlWKg771S
V6W/Tj4vzq7aWXgP2HD9IiOq67jEjafkLzYOOZno4O9+SvIizLDd4wOi02uLiGjn
iBHXdvLPUK9HAZw17xmKxo4Vfj2fwivWG0ytOEcq8dVhjTOj2MHHgdLod0QRKKd6
SLASClli2UqoCRONFqdArPXMc+9h4EnSGGNkVz2/XFx8XPDci2Y69h56qQpu/Hlx
hQfx7Ue7E4pQOVGamfQseg70AgiKZ+7oW4uFebwqT/i6BSgLqgDrcznScSRc1nxN
xGPt77PSSKesvOL1Bq7r8JdpdHLjekmGJgKqv2q9kJDSsyeS15aqoO74CITOmrSn
FlNBg/PvwK27F4wugY8phiaKG18/KGaoH+cugcvSpLgxo2gbpxFAX1Y5YELRhbkB
yfELaKZ0y+aIyVlbNQTHu/zqSeXHiDYk+mFUsYcn/scAMhJkxx1o/k8741YVNM+A
qK5KxkeLLu9HoGO7g0jD5otbQNjCLpAz7aHWCQAnGDNW3Xxw4/5Uus6YyJmtRxiB
dBISBA6K93IWnntoafeU4Kmep7WIx7pQ0V4Hwueg5k4IrdkYL7wxgnqj2YMF6Lsv
+UhQPEwAo3Vov1FRct/nsk86oaYhjiAmSHGk5PkcXqZwu3Q96SaiT+/0c2cyAq9o
N3728oJ/DZgoxHo0mpJaElaIyQWlnEUINDw3V1ngcOuA9EW8491rIChEj797+aYq
ZT1Tngr7umONIKkbt71287nOXrWy0N0jI/x3atNTvQs08u+8sfPAB4r3Z7gst6ZV
gtYU3joDqbTSmjLks1Pvj0gjk0dnWPo+HUDtSsCr4yW9Kdc6Z/jGQZqdw0dIp4g5
T5tHz4oTDeoGOVccjmJ2WhIz4/VWU4+gniG7OToAcMytS9jp0kUxN9DUDKqh2XDo
OrPVPoMJcl0qki2kRuKF8ez1bq3OVH1fh3DHxAWmdWDZqeQ+aILKCdJJh3v5aa0x
KOL9m2y10jejsSZMakaPYlr8eRgdU4cvtQntYckqJnAVWdUqXf3nyJR29BdaZY6V
+W+G+WRfQlEAqBdZovl+lrJlO6hJKbsP3UubAiBayo0OD9uP/P6UX93fB/2yFtpq
yJ0hs/MtTTH2j5VETWgfYZpadzofJVxV31Mk7U8B7dBUKfgtXfSd1ZvSYxTW3H+F
d1y3fG8yt4VsjBS1F0UnQxOraJBCG6UnMc7Ll1NqiDg25A/E/JkMofslNtlhDuPZ
/Lqx6uuFlY6EwnOsQnAPwutzi3Xdt3XE8MxwZI5i99J13BPwghhSz1ZCjUPmelzJ
3zZwSlA4fMLyYtgYrJbLTBwGyN54fI8+R/rtL9IpCzqFSlYcVnNZdxpxZQeekotf
bFpBiHxd59gOJkIhgHkeaLNHuVDAu1GPWM0aNmguFM124wMIW2lFYrcw00R1B/R0
IAUfYs64yzwtz2V0C3nbzmYfZ0+w2AlgFmG73PhTXVL4SmzLD4P23AzVO3OdMdhG
PEUKlOzEbomsMH6JJoK+4LJtIIB909l1g/MOgG6JoGQgIntI18meG1CVsiZoV5nX
enduS0nLX5AY+WXGGFozg/V7lB3zO145yKu5Lir9QkCYwp8B4xfmWBFYS8Ef0OUw
C4o62BtjUtR4hJOpGfBOOsosbIebPd8QkAydKMcO5MIPSnyNveMWOeZVMBEYFpuy
u+hNldW3w2IF4beV0Er3BRvZ5v5MYzZiZkoMREgaZMlDUyL1PQnaNcbBhvJ20cC/
sT7NFX2UewRbs+Ri3c0mZgQEFvE413nyW665M9VLjhGMiaAUW8ULCZfQPM/strw1
G/ipfhYz20fs6lwTk+NHsw3GEaRpYyxHteMJ9+75/GEXBc155LD/SvGan+ppB7Ha
Z+D4Lqgas85S9plHV8mlqT+r8HzruFMWogVw8mp+7SCFV/5faoTdjm0oUCIFFkLf
zgalH38e1+5vJoCspnow73sjnVXki18Hge2LTdOGxQa1wxbbD4QdKqZpGTPSEAIk
Ps+XXn0TBoox0cpXboAAFBhK+sqhKbZ/yLVt1ItCRmw2ZD4r/ki6oOP9KhPhmwbv
zhfjUoXF96R55uA/WTCpjVZshi+SA96LHOzeGr3vK4u+Gm3JoeDSK0xsi+59nfhH
5IsNNyZN6D8JwoIyACQR8xKz3FjPvCDW7XCm9+OxfUbeKJ/Gkmr/BGzQftUTi9cl
8SC1rMSMNAedoMMlDBencrZrKNtUsgRUfzn21xe17/zw12d0S7eAMcRilx4vUWjU
BwH/t83atVAvhSzBOrrRB6ZGs4CFo/M/UHQDH83nSYVgMWdJYaIsQAMDSiRjgJVE
kevzuYqf9T7/m7P3EO3ga1JFgUHgfrdCWBf5WHsp7JOGhlKEJW//dRLH4No2ZSlu
s9xIss3f8XnS1gd8bK1Dmu0TPh3IJ1lpA3ETr0hFBx49SvHpFx+fhkm6UJMSWGio
snUJAU/RBTAf7a8tz93b/U55n0nckftwBWeQpvgKtyPTgt2GBCih77hcQLbEp7Mf
Hntp6Y1/8ILUV6SYu1VpmAJzBvzy+cN8D2tZ28bshyxrXe1ju6CtPXHtFj1+Czla
ewWSKaoHZYJ2cbEH0LYgc44KWssmsdxZmDZqDLQp5Y3X38ldtB2RWXmKerN3g8c7
jpeFiV8mcv2cIwWqbJZZNWoDLhthVJOx8cwyNh4hQo8IyqYk+IL0hoVfVW6umjMu
N73v8J68hksjACwLikl0ajRPdVLJSWqeKZmxOR56dE53GzDXqO/dSLji8VYNitlc
eMcf9tvRiyWdI7NPHdFDMYMX574C/TwjoIj3LwIpuY15j53Wt+KC6DHEN4mcCiLA
uU9VUySBu1I9cXZxBrjjiiUtBVMWmBHZKdZsduILNnJ1P492rZmjsgXkukQf3Zl6
yrU7dfDJB7E7wg5CdCZGrbr0VqoLtbTfuQ/t1KelRI0JYe+t3YqvLXxIqrWA3qFY
6HcmQrS9rHcCC4Blx7Pz0yiYG6sMYyS0x+mgBprUORlP+pTBrNLH2430BSuvI8gN
t9mxCMBOzyz257DQhqJDiPIVdG5GCDfcmOyF5bQSKS6aOechU7/23YQAC5ACu3JW
1BBXxZOKe3splFUXpniDKGfdG/F6/j92ezboGo8Xd5f3nn2h6Vt1Fc8jBNdNQTFU
lbLOXyXUsS3UT0BXlDxyGGlbaTfbZGb6FEkOMqMNoex8U99pWZMzgGvcrnTVksGy
slumT9LGYPWEetRdinjRSXToyqGbRVCYaeED9M7ZbN3QVmY1ez33y7B4LykqhIqf
Q3YhICFLQeHY8TUo1ta9YZW4BgKtdijIVmhngXeWf5Y8fGrj8z5V3AVH4FbihEfj
FiIYk+b9MAkxm0fEDTESv/9Idse5ZFAmwBbRt4XDkcAVr4YQwQgGrztx2kDOZCu7
KqVuPrw6W04EHN0ltyLFIIPmNCGPkyd1YCLR9FkxWMecT9zN1BtR/cPUgIlluqBd
+caTjRdeGXezz1tBjWO04ATDEe7ZHTkzlJJ87+WSs5utfroTR1rOnC/HuqJFadem
/sws8pXzHEsUVy1E5DYE7+9FVNOpqW4qwckJUZDfSeHrvr5hS5C/wjayE11UfH8L
PxlijeyVFRoYJiurip5Lj1CB6/7JZfFd1xsMOUszSFF50rQiWAcEVB/gBEq4JIil
e2wVUPxH54LjSA0wP12yBU9HfIonLl2eCjNHTg88VVxMMSEXznWhyrqh1xU3vXDv
FqW1hP4eOXeQIb1exPcmTyllupkTvtrOCkafaNBZgY86l83y7eAbo1DEfx/6TBh2
a52b+w6M/7aUUe7yLawVuYRDXpwkYaxUONpNVtOQUMzS7LdAuIa+5JMs/sLELH00
PYU+pR7UiDOsyDAxzoYQRBwHS59tlgNNPelJYZDa/uay8ePDqtv0FtT5OP1+MaoN
RVyZD9BxAYHtmFKv6oy8/g3o6NrnXqto87oTR/wFxkP7T14b8n7IVoXLdG6DzN8u
Q7xG7NBcdR6TYMpdYPXjgLkIUWFm6jZdxmePxpUuikY/dOq8a2MolCpVqNbP2ait
dIiO4bllVXV/G1BXmOPo0Qg5oTRUuj517Ed0RguC10RNVwem5bWikKps0cB+xcKJ
N0OUaMLrlfmpUkIRSNH8LAXv37ZISKmxDUDqDgT9NgYXcnCHZZtFu2czQS6VUIoC
AIY3ruu/SgN/ZiKuV0Ekx5PJuguHnhQLfqBksZxEMdKvLLAirREWSk3CW1uVa+Rg
0GxfD+RJnNEnp1/BzO1hz6wxMJWZIxmdTNjG8R0Zo916IMg3OCVS5bCXV3IdcALR
/pZeMJ3ZPTtjH6fSUxGLR4FT+rq1aT47tGXUUYb1TKHyCK3+jUIJ7hoJDFi7MrJU
r9m5U6blcLiwWmaVQOqXvEPNj1Mj4SSW51r4gmmPDBmvebLUx+wEGR7e7hUcqOKn
Y4Xk8fUMI5LmxPTqenw2TaCQ24W/+Ykm8+549jovfh7LlRY87lnldzKW2zST0Onk
023buJ9i0NEZSrv1G+1ixsCbz7GJrrUfAOYzHIbZYobLtb825t8aSkGNnTN3xwWk
24IwutCjXBI8zfUhzlMYcpOuyGxOzcSwoiH7c7m3mpH03io7QWKLaGwTPQv8rxtj
9TIVHbipnzUiozQntjaKZKOv9B3ASwNUZxP/i+J2aLdQiwqDuHSzcmjz3BRYJrOg
R21SozgvzDUIVfziPHHpsiQWAVno+Uw2vpz1nJwcwGnh9zt0wB8HjckajNu/t7eK
MsR5jKNssmBZD+9D0SXbCjdqlW353s0FSHUvD1jokJDMKCdbFzIdt/d0sd2VAE3x
DRPdjBrcSOgYgyO6xVoX/GuOfCss9By0hlkRWn4sdsNSqlS3L4JqqEnlxjZjPVmt
dG99rZalXVosuKlc1G1ZIoxFKpzVw+s2KWcKiHIvgpXbjNXq7j4ved9bxuiRVQbS
0xKGKZckGpMqYwviJ7DmTo5/uZKG1SL0p9XYLX36jdUM8gXnt3gBJWXFv+Brjsrw
ohC4d7ebhOB7OCoFEmB/IOTwIyWFd+wbLmAvmNgnMZapGssWG6G+mEhUknFTD/5i
VlI874e+7kv5X4WSTG7F3dA4lnTzOqXypAijJr2dmq61ROuHrQKeWpLWiTFiO+RH
8OTVhNzLcQk0jEcnxh4kkrrTgJDQho34zuesRKu1+1Z9qoY4DxqnmkZ5RHajRtmi
0GTpn0VtSlM7gVsa2R26WQt9m6Z1Mkr+d4YCBGIBHI8GPj+PL45KdLJCrWP4h2NN
qudMApHkVt9C/bJpinMnpBHUS7c97WlMJOx7XioEBJsYwrXccbfEVsw+y4jKQ+IH
kPtEgsjpB/Y3QFtwl+J4mM4tQ4Ab6nlraP0EF4rUxBexc1MEHEkAZloBMbt2kKl5
l2H0KwPwUbluTJ3f0wOr/A7FtJtOjQ0lDHSSXuOADuLeJ/2uuoP0HVci9SMMyplf
p9Fsu7PxfDEve+ssb+PV4A/QpUIxRCjG/T971l2lDkInJh/lQ2cJ9DtFH6DGcxgd
Wzuwjrox+Og/OEToSnF3+4gEHcEqZEwxWGAjjayn21+w5gCZl0PusVXbJp9VyGJn
HPG6OhI1/UcSBIbRrGPhD6crbjva4FnAH9S3lVQf7k+iwvxrl8+BL+V/LIzG/m9e
7wv1t7e94V39RR2ni2IuXQtmXy6amgnOWSIfcx2sNV2b7mGItdXC1fB7mzRJs1Sy
QjRxXfv4TlnG6jsTXl9rkGKKnp1ZJw42l8db22nzb4CtHAgXShZF5KNLJDIwdtkq
Gu0swCYFPfcKtjHumjer/Du4v6dKQbTT6Ld/ztt0qSwAvTkdAxC7o15M25jVsAO3
BfbUZWMx+9dWLTGs3GUa5gKNd387Gzgn1fVLNCckfjI51FVo37nVZaShxa7pi0h1
ym9jsQ2auDGwZp0r2dYaJMeYVRB7Rn+aVsfc5RlDX6o3ZknIn/M9O2OjWTct9Giv
+G025wlPPVepbAxaOu4aWcH6cFa+Se3R98qlKSJD7PbuaPDsbLJBFDv1gxqz1ZMr
l0lVDOXepup3RH0D/UB+vQBVgd8jFm620Oo99gT3Bcd3VldWrDQjdniN8bqm2jKG
v66IEokp/jg2R7FPZXQYMO7h0tD1+sMNbhX4os12zbM9kXkO3OGC7cEnNNawbrAH
tuMxTCPd6jGsUGnwQQXYcZgAhzAJqYVfGDBwBTfeTCMtL8ZsB9qI720dFzHrhQSA
sP17Pr4X7uOGrwkdvigA0K2n6bE6jwFZWR2mxNPD8hL0dgWLE4PN6YBKwQuuTmST
wiQ/DWj4SYlFmXWWXVaI+KG9FyjIT5K//do7vVOwsz5nKxlUwrocsGABmirpiAkq
XCnX0VLX2WEBDODD30ced7PyXGSeSUfeLA8jdyUgOK2ao/4A6BMJQxNPkugEOm4l
GAVv6nmSB946UAtcBBIRrv2O45pL4SJQpZHpcWDNQtJV5gR8buuBcCojcLJU45Jb
t8sbu/2UIfhZFbwT+CeoLsQesiOStxTOQGEAM/wooUjeBaRY2QRdidcPlKtcVnkf
oBC7AjspphTHX9FXK+e6ZeFDykeX+Pf2CbiqS5Yb+8AQ8WwGgzco6Gj4mS8zssjc
QW8ETvGTyeC4THzt2gd8S+jK5WBcR/H42ezRieVib+EK7Z4ubJ8MXrKIvyGDR6tZ
uMeTh0lRfV8LDIaqfojUXqvjilwumo2sg2OJegPbJ4t/fpJ4BkEpq3aoDF4FLr1p
Jxw5DmsziYKaoolIhCAiX1f4GHEjZyhsSM4obprX3zApV64HeV6RaznCH2QluYU+
IJ9P0OBWXAh9e+86pgDHNYFanomVVHC3iycbluAxTo7l5knDmyxaUNih6NUyF7Sn
t++RPD+4JKOEeo2Jdb7tFydPdDHwXTuJAxvwTx6DLN3loS6tVYZ63AucgYnHf9nS
BxuSkyP1AW4DUU7m2WbXWsLBsXXwJ6LlQyn8CGlzYWLDkQhxO5LxaYHKyxNE1aAE
6eejM2PTeCsilm6t8D21huIm8uwAkLENVBQs2pkehV7NJMU7IMb8Y5vl4PBN2z1X
jAmtDeXZV1NcyKNpA18IzUlkc4Ao7yZYdrbWkh12OIUMmg+8OWp6KsjdTX/7T2cx
eZ84e23e+nu+omUb+6lImjYdY12tJCWelCnEo+G18L8160x/MsBPqJthWddmvMas
ROWxkuSpcX/vHusxJkIGNxceB+QTZnl6IEZe2F0y/GiazMowiHeXi2P/Cd3f6xUq
MxX7xrvuc0E8NN/aCG0uZDm0Y8TFT5vonntX2ExYeWPPPol8uF+zu+WMO6bVpvd2
5yxX5SyFZiDDiQ2CAPDQ89Z/yf5KA3sPwpTipdpWvj6zRXdr0i6ZXyHCtMyLPShG
dlEzUt8GTT01bEtCdwgHwiNMF3ATUOjg4/EtOvW/d/+/lwbZYaVi8k3I78FxZePJ
iZG7wVtBBMe8O1PflSVN2evKvP/sAvdwE3M4hGCJUuUedv3x9AfChUvZPpCqpCkn
zJHjSZeZijzpaIhFljF5hbxRxIkFig4VBD/aZ2wcZSmuRQlpKHMBnHVRMQ4QbioC
TjwulAfNlf24FjBDfaaSuQ4Y9T6IzIdQQqrWn4+m4Uv4Zro3RGRFArcgdUAxYaJ2
IjpPS6IqXtZUMlYKkxOCP2d/94Vo8tCfXNl3nHjVhjEPS0f1t9fhFi4BuzDtG/Gw
afLI4LqD96TQ0zJkarHKXj+Rmh38B6Uk512zZPiaMGr0tlcTYE8F/Gmz+WEcGY8X
OxYIg1ovYZK81l5mGAcsy9PmV7G09S5u39iCtSkJWItDlJJi6apd0E6UeL10CpvL
xEkwVE+OV1BtV/c9M5fpO4flC0Meinejn4S6pHqXhV8WAuqy4YJQg2KgrmvB+aRh
2l8Usc+Ma5JqWVV0VJzVfz52ws85oCJpFLX2mR3mLSzLBjeBgIJC7um0RIvnHY8q
XpfP+HCihhiWO1zepHEOteQwzTT1V3lQc9JP3AVvVxJGROIXUrRuqJQcN1DyH9DG
jjxc3zLOPHHUZM6IX7a85RNU2OXg/Hv4NaQBvlCXJE1SxdtQ9QsfE+xGM9GQx78U
2bEGfl4bcfwv/IWWpf+abclTTYjZ1vk69McGs6hjLtEGi7btUgpdj+phIfVbHI4w
bc+78kenv6Mlu1BxWKNT8fP7qMYwhixbXjLEUTrWflPboxwk3BsRGl9FZmSm8VjM
VxelDjsJtUvAGVQjJ6FPIe75s7lH4cJ80IectfKMK5Bhe3fxaSMP07z3txhcB8GQ
RDnSHUlKJoQDorvhTrWVxJEg43/iqU58ley2ama20npa9s5gvLaXM7LDWXd09rHL
4HcYAhLklhFFKV/4jFusR3gd5otEqBdjBs6C7m48Oqd9nzOFbBbysd6mx6Tg2tOi
wDIgS4JcYHExtEdJCxYm+SX9PztYdQ7QoojAyifNlBndDQn1Am+vPZ03GAcojzdb
yb25oE7mT6OWZaLFBiS/SaS49HyeURuSAe5sm/CC1sAeVViayyy+fIgcH4VVimgR
s6EChkEqvc4COdYp1NG2tNhrV0HkzdUGgnN/iFlMVAlPYhmGVH3kf6Q0/2ai5Eb1
tEIFZujblCfQiqU0RSrG5cXphpVecHLYTdrOuL1Wl+qcPIzSUZPU1V1R1U/amN0o
DzsIceQ0YPCtdykBpDdLCrvVqKFdW7ajgEyFg9qwJN3aqJDltQ+GJpKxtcjSJPZA
0c4wKXr4+A9XNDOYx5YAHtoxV0Y3vjEgw1sOFXxGoM+2r5fGW+zJgmlO0+fyGZfG
oOEzCkI17A2F4K97xjm5OGTK1KAcB19o+to9CL9RLGIGgcrromW2X1jeUhSpALfR
VsDzdNeF9aeuzLzwfluaZGotjqMQk7H1d9JTYH2setvH60lOdxKMZslle8otFW11
ZWS0lcLyEQH3BHy5mQxNGXV//u5AgKsOYvTSsfCs4UZcYNRgiNBZhmVM25fSX6Ot
tnCgduDh+q99xUnJIp49zK/VM+Uw5osKjTQONmneSCPBIf/76nFeAm2icMMpLWzU
YFC+b5m0fTTVL1Jme7cfKgXlqNCadS+ze8mcqpnJqSDkgdWYIlIjbHYcraS3on40
FvtLtfB/yDUoUywNmzKu3MtU2itPWBtetHeCH7hKGsY3hwpUMRtdDqXPUG6ZN6Tn
5V97fClEiJWeblAuN//Rke6kohNC3BgpCgtiIHFpNTKR/ToHyAX0ZPBoFXltgzC3
1RsuQYzG7b+kEWT4qvyWSZ7GJi3w825MhhYZEami0lmdE8FdDFYYcuTww4r6V62x
/pLIBAQ6X9FCYLTZAKxcBhKjWoTWdFyhyQD3sgCt+ayNmKo2HOB+xx/4Keqr3GYk
WkgusBZKm0yVCXvItKDVJjaeiNeIQfLPnneSNWQ5WX50Y2gimbjksDOsBXYvc+rL
VY9aEnxPtdrMFuljHzJLQqjVH52+J1RuG53AGU1IViCPefr6eGKttRnayqnZIb+v
/na1Qx/BMHZXP/8EHlkfTQVQnDhfoYajl61+lmHhlfivjA8LuqIi8nrBjhlmk+8T
Y2cXl0LiHxZWDmZik0inqjsJ0dxsQmraPJ1Ni2+mbbd2FhDww1izYMSR5VAdqGVL
kZmmND1MjeqOod4TEgVc7W6hPqVTUZgje/5DEFoPuZE9yH7dN/TkuYZPQJP99MP7
mtO0x/Cmp75HQnzeqUScimj0PjIsFU3BMLr/oQR8MHpRd4/wIMBlEkJOzvEe1Q9r
ivz7PThyMyfI+009jJRTHxuk90OIpetVovmeq9cU5MPhhVvSj2MuWB3fIqL7bz4x
e5kJhdEghFvTcvGEtntwXaSlzWaKcU6D1615xjo5BJF99MRLepHfBoQ6dDep5zdM
4S5Wlvffn+Of37Z8l9AqazIrlxne9PWYjygLpazQ35zE9Kfo7AMiaKZDuW7q6U9z
wD5N7f4SB8ogQBfDyxXDtKggYMg8VEnh3lmC5wDVMLzHKnhNlSVXd2T9qVgK1K9E
rSwcvuH/xLP2xFZ0aB04xGPS9j5LCEWLo6TznnvWKan93EEOHcpUpx6zJpHkTp3+
h95ZFWHyDfrjYIjK5jb1zNoGtId0ofax0FQu1cLMOOM5JXdMeRPP/Efsa8/ziPxp
cNpVshwRronXezKBr+xGEQovCV0hIRELWnGg+D/LySFZ/fj39SQfBP19E4C3IplK
YUsxJ6wmM/rHm4ro5edWKuTK5654qJIThPeuipIWsNKHUz6BIEZNuOMARbDkeHDL
nKvOwBY1crt9brWenNF7Kc4kU8/03bc4u/tZVuumyxERULzE5Mmag4iFua1Ov7S8
yelD6j+xVlYTxdgpIPcEi2p3PWUiX+kzTteDkuBVc/KN++YmfzcBAQkch1ErJzjf
6xCb+Rzct5tJaX8LapllLNN7DYJmF120NaYrNA2Jbivw1QwFiNtx2GwFP710vdas
K+5nn7FYlwDsRQEnb+qWjJuwEkedIAveYa8/ECsf/K3jKgMAA7VDC/vq2Xuh2kU6
YUxoo7jJz5W9m39zou1eZQHrLkFBAdBlWyhHIwiIEWibDI+HjP6VCfdOOe0P5RMU
AzXoI/fjFOqyVYafSh5dCWyQGDmN15TpvuVuWlMdvTjsEo2x5Dbn0lu55X6up4uE
xh1lu+VCl1p7n9auat8T0VOLVeW6FZYFYP0+YwswOqocJz7XNtTUf5vhpoIDVhbv
f3IBVpFaks2O9dMFw1d6wX9sYviBlhUr/yj4i+QXCWw1ARm/6LeN9pxolmoEFZDr
3sOVUe/P9LkkUFb0USAGLeLPThdJ5bFn13UDk4CcmMpXjFGC9icuZ+ADugVONae+
zzzxeloCPub75U6SoBZyBrvY191Tbp+LctAlMCyr9KVtsnyTBfqWy2OfiNl0OpEM
P93mBLm1hPRteDnI1sZ4nHysTOwiznO1/LR85d+3vhAVyvyKrrJHAkU4Pe68CCiW
D4nO5HsXcilcDhfq1HJ+iNYX1JJMOrHGE18394MT6J3wygsIyqRYiFuEzpBGUPov
x8znheYWth9CoAkXQUxMfPPzRKC1vuSnmZ+OreUDfjMu7yeHJvC2G2gZwRDPh7Xa
Vr2R+7agmmP/G4wuVDjljjBZ/2J2wo2tJsknd+gjaLMDZ3ierVVI5xc3A+NlpUE1
4aNiBEyfygOmOIKsz4WBVj3A0M3nRVCZ3lbaX5sJv7HO2af2/P+hIkabz4XP+xEW
p7nUgqcX7bmdKT7fgqwAvLKDu6OCSJcYvHkMALJK1glFZUIMG8gPnoxRZaWBd6bU
mW4ZKq7b50HyY4Fhsgbof8kl8xNk02yepajlHuCQLOQcZeBIju8BsGvZfGdw6592
mQ8VaGPV67rl+7MYaFXc1vPXOiDMFYJfbjIFqVpguaABoOl5hxOA4Ww7SZdm3rkk
N34t84P+Sdi1XEYVWnvJMEi5lSP0LUZQmS/robbBYC3qH9oBH3qTZNshsOIl4pX9
FmWeUbb3QWRvFFLEteym2leElU/CM9VVv1gttg+J+6GFF7dJCv2r+1zKV//fo0/A
MF3gYDWakzRX+sS7DA7Ul8d+LQwlXGHsraNEQu7z098HvO9Tscj8bF3VBYQanb8j
nCVRVFa9qvXabiw0EG8FYuYLdxYhFQtkajuKEmzYH2NSmKCCrzWCCk75cZppjd7a
54ykNoct+pCva5GCsltmgRiwvhMxrFMyAzg4ucEsgcDg0FESB7Sv89AWh8U1+LfH
iJuEfo/XURRZqPj8juTLvMK72n+j+R4PhPBwRkEjZdt+/YtS+BIEbn3Dehcc84U7
t5sPRrEM2PpWb2OFIcOsqQFb5bxHbDWIyh2Id0xd03vBj6ZoUXFYKX5zJGpGkogx
JORQXFho3j6Ual2wx++MpyOVu7JZy+dy3UkQmluaibOAEeIl7c72o1cVqs9sp7cU
ISPDEfkFqGSeirm0PyHjWSfDwh/GKTie6UXIYx9ZZfv4+Gq904ClCLmHyRPh8E4B
wRl6O3YNHiiJt/kDjlDipcZk2hgSpDEMWwol57YjtavG+cahz4sf9gWyxVXHhOYl
46u3XxTkIa1nUKyGmGj5peCmkbg4S3IVOOeHCqGVFsYEn0PKBKBilDHdJQiwlCt/
1m0HxvpQLORGmAynNVza8NJWjhUZqvRINDnv1f0NTZJkt2BaKJ6e/z6x36zLYZHO
UYUWWbH3eMihEf0aJhYc1sS50lkbITkvRHFXu4X02Ioy/acIriGV15bVKzD+bePj
wbGRhou25DQMmONT0sstb7agMk8v0Kn4mzPALIfPH4oNoKmZvV4W5Qf84vFiqCmA
fQIXLQr8L9pClLMgCra1rprKntGc/TcYuOnS2N0lPQMlQdw9Rr5RXa1CvcXpNnMs
71DgWuzfuPUNKO05OOdsNk3BfQJKgIWb4FTDUuVFQQMn/BEIFRYtYD5kTTII/+68
B2U2Co/DxmfEWaRcxQN8kFwaB58S3MRw3pfw4K1DY3DjVXR39bX2GHnq+7M1RZaM
lBlD4R8zE7wpI1E5Zwu9EHPs14xZXBQhxc0LtwBR3LQVqGaMf/KfE65wXETOLGeg
HJmBwH4ckmt20+65ZGe/WsMxdtBLr21iid5ErjD71Gdg+TYJSDlTAhkanQKD2GcV
p1wGNXJbLhdYmQV3jby/qp844QzvY+aJCSNh9UACzugUEchBV5wMzK4OMUuvIMDZ
Agtaru2gEImDJA5GY3+Y+6nVLGSAuex6/ONmtBvbYQtLRM4yUxrnccrZbjA440i/
tcWFD6q6jaul9+dnxZ4b+y4QDsKRvN4jn7Ys9Z74RIn2jnGn18NLfOwa3QUfCA92
jWuhkMK5/MVIVo8VfcVf928ZAJv3DrJIMZoMpj5j793xjT6ew+J1WmxhUXa8YwYE
S42IS4I9Fe93Ar9ENmsff7BuJ+t9r31x1QzvBzxNe1wCe+4bt7JIox4uM87LgS6K
12jM2/ZMvuPTvlGyhUZKX2Nokpk6D4ZrhqAmaI0D5uNkRqgCGDt+QD4OSZs2V2jS
amBfidcitNl/3SCr4ikcBR6aHH+A8rhrycOiHFpvj3u7YeFwCP86BeuWEYuaOcAP
HYMigJkBMrGqF5mbGuQzEuJjc36zcGUZtzh5jlwpskTF4PWl2JJ70A8dI6lC7661
X/L+Nlz4e6WBA9z1WNNczf0NcwijC5jSVF95kL712cJJm38hcEYeswNVvfcqLkBP
F2qrnSeYl2bQvjhZ1JO7TrGKhzoTh/oQrfovNbj1H8uVeGReXduRThsaM0GOrD4I
TkRyU0QyYPMzi8USNjmB0UnzZ+QjGnqkOT27o8BmWMzXqfVbLMaj1DpKkF1TsANl
BsWkP8J/98J7UWHOBX+SyZcFx4p71ZgV2XnFgF0KtNWBaqAC+MswRcc05Q4oFhAc
jzmAEaZwIV5qjiXU8a+z9Ycke6waWHz2fLlZKMYYw9OguYEf5HbnMRoe4vDKc4R0
x6tiXwZqHhws7sbwBX+qn12vZI2Wdy8p4bDomUIsilknfFenRnILKp7eW/pX1NAj
n3jt6BeGCp/ruvmeYGZMreftd4hCN2JDUZ8uvuVteugN9snLiAFh7taM2Br2X6bm
XPtCvhJMZV96AS2HQVFfaZoLWvR5aoJ35Jq0AVo8Xk9/8WvpAAMTrpNQBeQBS5lN
U5O3u81rRVsHVe+AjmY7MUOFKGggwPMMlHZj+wxg9WjUqabBTWmkJx+usIwt4oGv
E+zRAVReDc01btS/2+0FuwexlVG/ffaoW2eyZSNyA1tqYCI+BELWAq8J/Agyh4OJ
eJVd5tu3did2UJe7UVDaoIXeen43Gypv4O0MPN8lQ0k7WTya4iM0tzKVqHX0wnIu
eKqTqfU5ncbpfXyfoiHJTHDE6eTJ6vSPnOhp06tqF/ANHQnjEoEffQw7A1kEd3bR
yxn3aJq/ZqiCcGQwNd3Ock8DDmk+ZAiTKInhzdjauUKctbBg9qY5Fmaq/Xuju2x0
sXqHNehS0uIvGiDLNaK09z4Bdap/1KIK3tdfigbgBiITr8lUTaKqhhHjdRjoQ1Ug
fThqNtWfqQpqAYKeUZH0dDfggIje81Ay6F1xLaEzCss3PP49aRlwGOOegD1Old4D
CYqYZQF5KG65GKzlTK86iJyQhujr02OsCttBkFQy8fC1T9A0huoRsQaJ8VPd4Xdc
/fI888SVAC923LQd6ZXDMsr3cL6LU8dZUQStvoK2eWcdG+8vAQjkBmJylWJ3H70A
NFkihsHDSO47YIZz98fVh2xHB4rQet3BLZ8Gi1QA5bhfYIlDF2Qiaw3jpR1o+B8s
wA8AUBwrioS9H2ySCt72FnnV48JGvZq9nPgG+G2wVoMJARyyg157MRloc81x4joH
6Wg5Dq7fioqUi/pxaxASAeQDdTtU255E4F6QBT6OOmKjW3QckvXVxjOKVoO72jTQ
CiNfWItjeoOMOZMHE6PWApchnY9iWwwaEpxgzWyd1vcAJyE7E27j/aXANq7UWOl8
sZREE/fsj7M0PO6/Cz2k0yjIF5UehIlSwc6mLPZMK2YchDCPrHMsINGA4VcKhkB6
rnHEkIxbgLCntFPItBPq8xtDI7yTyNfky1ZWfTnkLKN0FSN+04TwMhAvm1cG9/cx
IL2OdUxoycSzFJOh4q9TmjFy+nwQkv/eVkKeONS7U1EeGgqB9vL5uIZDX0LckBjR
9pMX2jwn6X4ei4i+YlccsCjtbx+3CB1WAahm4on/Ow+mLwMDmh3obz5CiEbAWZyi
/46jG80kMrT9KfDZPJrqpSTcqkM49xNQ9v7w0i+bU4OCTaB5dBelG+2t9uGVEEey
y6jJIIlfxp1FLh8W5l3fsJktcYH8b4HPdPzjJTrSyQ0tgN2yCBXid9OPMnAQyc67
8rPFtD4DT+VqNb9JqnlYlhveVXUg+pJu9S4ctZkUF3+d7mbtDvf6tX4yXPu8H9YW
OK/xSIHLcw0ryOCc4kKTMQV4M+l36YSZZoS7dfONp8eaU3rqoDxalE4MlPz3b/lK
eLGz6EqkqrZpHVv8I81h87cgkgnyJqO+ojx2jElg34z41roD6yn4MD6fgO9VEvGR
lnPJUJIQd/p/myzpKvHoizdc3dtDId2zVUC8QF1jxlQzgYJses+VhKQL6X2hn8GH
XaYCZHhzg9a8QlsDGETHwUhIAfyw3ikVAbPG0iuz/G0GVujxd1SLJppXUCmW8nUZ
J4kjJpL9Xk3Yz27pOdSixamzrJaw+Q+8EA/xJv9cdSuU8wAeGqKQ4g0sbWUuWVtd
km1CK10LH4D6p/277mtGIWw5VRQq0QyIwAOXzFSFhbEVc15vUoQFvPU/01BoGphS
nLnwOtI0qV5VXwLUQ0b241KRbGcHcVRbiCUNmuCnbEundiicfu7nGzPD0sS8fYhe
EQ91YaqqOTGIqgONMeZ6D+AURBXoH/pOlPQcfqukAfdcQbjuJwV3XizCsIWUCdza
r52PH+5rdw4uab2UrzI5qFGTJqqot2P8nKYXyOFKoLdCDUSd+2C4Onf7wJuRMs/C
KlETjDP8aOWo5yKy3EwFWFb7Bm1ejVmMC0Ugy76Zg3bB6yP3fHTq7IxoDnmVRJIf
27+/HXSJL8SS6duJtsa4J4W7hfihhyPfpwK+qhNKBzx4R7FykVZ0EFWr8koa6M8/
2THAMRtPynWUTKHZ4z0oUQLVXKSl66FtZwuBP86ZjeQRW2zjX3hlOq1PEno2a/pA
ptyJq9s2Af/tbdGFcDv/2FDtucmpPnDPq/FDlqigC/NircyY6V2/2G7/bDQ9wola
tx6QmTs/9Bds+u/XVIDI06CTWpKEzi7V2LjfmxwqJ0yWFHdIn88rHMy/jhzdlDJ1
Znqgc11iLTKPK6SYbe2Nk1Fwda6usKguHBtb+MGZYo9dYX5bmJD5lCNzAz+tPOcF
+NemLK5jRHrDPBlSSMXvrHDX2zlx5oBiE7BcUeXXbwgjIiVPucSOPZBjrNK871v+
nkMnYBdohfwAd2shWvbC2hE8chx4E2Xw0H1NYPnzI9vy56p0hXajS+70717hYeW4
ICMVlpT/zi0yj7AooJuG33O41mUcworD9FFIdSwEJwh+WHQPVqrYHqfeNvNDAGNi
mT+LPOyKJ3CB5SKMqQeIORqe+33rY5XrGCya6aMceWyt/TK/q9MPnxE9z4t2B/jh
nXfSKuHwFp6fOm30kLa+M6HiL2lDc/DIqpCX84M4bzFyVjeyurrpp2e5JcBvudzq
GrzLUgg/4cnRUxnYs8JsFUdyVKbjvFC+bF07e/AWiHT7dKbrTVGa7T+sYXd9gBmM
moDht2+BEuya9vFF7LQ6U8+ImBnrheU8Z5aeV3ZFPKAPGjZs7HDwE6on4nyOSo1T
AGOKkxs4XIUZxpMXk64ipfdIbgL+BvHJ/GV7c1K7j2BnOEdXsCTfmgerU2lwq1PQ
PS8dDOqKLv6ONyUIAyX9c4fpSrkc+B17XViOY+Ea2CHXkCo/MX6b5KXXBMr0w9f1
Zq5q/wk8yRH/7XUxsC95TK7Ix85zM4WmuUZ6ztImWrIqyLD3hS85bJFJ3O31ZXzG
k6ieTqF+OpbyyURejV1/v58FW3YUNK7d0kxrert6CJF/kjW8UHeleGaNQsQGjBpc
sG+mevvQ3DVs0cRXV+3XtIq0wzUDtanjivDJi3pWRzIN70KLIEOThPxCo7DOMwtt
Ip0M07EofznU9967zu1qDHul6Zl2Z0iL6kk97R6BHz5+vgfqqZI67jxiteidAnIC
eyQYAA9UqElr0AfVx8Il32M+XkuMG9lLLSCYsKufpk44peW6/LqJl8RJmP3bFNFw
1ws+Eu8OlCAf9r/Khn23UKUxmkIFb2w1kPSC8cyj68eluaQPm13GWSzT0i3dCP6Z
1XcDLixUPVGdBsBNE32efHcUOrMhrheUS0+HXyyTlayhx4EImlKRJv+oAo2oXFpg
rdxUQ5hB7xDEuFX1Y5Y8wplIUyKa3lrvWkjOO+LlyFiZ3YbFlQsthdfXJ5TA8Uzz
rB/rzCvPvBKRa2qL8SWFnqk9Mhb/CZIY5ouIjhB0ZhlPEy2EBeDJyeLmS9Dzsq26
z1phBDbbclw5FQAyYji1UVOM8wheeUAWC/3B0b9Q5/9lDqjB8FjFeeb2YGIJICpw
iZYbURz+maaRAR6IStXgyIjoj92BG0v13EgFRQKZ3XJSoYNY70Q5/Rm6L2oQH2JD
Gv0JziU9MIYTu21Lk5xtZxaT4gOfVZf2A6H/SxlDayK3jy/LUkvSv4Rvea2/hEpV
GbGKcdoUyJ7hyjpqCUR2wthOnzin8TlrY6YiFc8b3kxQBgeysLIMMPKb94in2lgr
Z2ZQcsM3niBtbTZUglLPzGXmWohYDkexpfEyaXVnQWoeeHOjdkkaZt9tCAvE5iWO
FkkUxvPgx32wxtAg4xHuemBh6zqgiLSKuXToELEJMJcfKitmTn8ZJGtp8NAYq9mJ
PuNqmJ28EkeEi1re8Gw+ldERwe8qaUdhUn5BcwhA9J3OfBK3KgW3Kl5+EzDB8hmw
FRpi2zEItd5Z/cEA7uzeQhmBHRPUFsLJfpLwfjmyjd+IiatyWZzsxq1nib6jUyq+
7WGzzGfGPv9CQ4z+7VjBlgoevvnYtjvKULD0dvI+Sgbd0FviKbhY5E+FPQfbNYu1
ranC/+emHzfvv+lCL5FM4ETeKvC7agG4rL7d2d+nOROrlsbIDUOTGYPrlONbs4Yn
tWxnFcQQ4LE6EZoHgE8lraFuJUFSlSAe3xUx2sEKeuz94+DKEwTBk1MC1om2rlLR
N/ev3N8n+HiCE5sMANo7b+f7W2ZCGtr+te1s3VYTO59unZutlduG0P9o1quwTRAW
59JcHfzR2o58wlV9hnJtylkcvNpAQCzrfukQD8/9506y701uR1D71jkCaB37eVnI
hODNmij5zv9QO0svZcYsmOwVoaFzPt2ORYh62MimJICT+QPzfo/jnG8vJyRjNw0H
JS1zf5ZNTKt4EGv3MaHcyZDAzdZS0BWIPq3PJxjlSvmy9h8TpVFInlan5g4uOB8e
u/J4ZBx8ruSZiVPqCogYldpfc1uSIoB5hTlsYImYklwJ+m0PSFSulnQGWNHMcy/J
1v5xweNEsyZhOmjUKSpkDkTEN6DJi4bOBhC3ImiA3k/Qyv/ixccHmk8F+illXqfn
zcq3faHfQEfwSux+BAQspqYe0fWDgD4RhpOa4QGsfsXVlJxA/1q15BhaD+66CtbB
9JrKR5l5ykqNsFZZjUEjHPf/GORbpmNl9dbcNWzNeAnjHbeWieL1qy0RjKRCXByq
ZiNNEjuVxpz5Ale/uidL8FeXE24Vie46KgJ58ZJ0vwvzcItYYOUfxZ+CEV3+mqEo
90N/916koOsN7VyuTHIa459qMvDmapAZ9mtyjGObHwwlP1pcmBRI93pcBlP6nRA0
4yT9Fsf4fmeHA+1+pP+pWJejbCk56TBWIikziNjEK7PtmVSrQNOtydxu3s4Os1sJ
MMAAk81ZH9/D9JqH1f39uHc4hO14Viv5h18ERIbjsujUHlc6Ak8QHPEd2okfF6Cn
eKP0mhDy7maFQxxxdcuY+HIGPTUKA8Rks+mS5o+Ne/LPAtxK+uGaK25n4ps11zUo
1jXTruSJTzKTy/FD0HE1FYodAsueEJyel7l2haQCJ4e35GVjRpm3x6ja1r37kKoU
mvL8zB0N9MRBVOWjMDiR+DBE/PW57N+RKQzq5HCeZqTPmF+evewZ6B4q8wASauZD
tH8lOt1exQ/Tx2Ssxo8vclaCgAb2gz3TukiALlrPRDMKnFXlmBiTKUE6zinsj/rj
tehMBEDQDUkqbgBNhoA2JogUW7i9+U7mw2oC0Y4DtVYDfYRxZc8SFsu4bE/SNwN3
twZjq2JrPvOAumjbQEhOFW5QUfTxASUblffl3ZuKa4nbyywq92/5SrxmJCM8mcM9
3Uw10wKiYUPMDZTggAhRoptMFMIsfz+YmvdDgSBb4CHOTEwmFEHENedy09CO3jk/
i+VRkLtnhKGZ1SDBH8NKJ2MlosXzQRkUmdTHJSnfmLxeD8ttnsn1qEO8iCZKRnaY
GtV7pOjS+nkk5mLfuwLZ/riOHbXLM0YrnTduRDNGU8dZZ4zpHigQ/mzdVXdouiBO
BRNqlv6NAXT9zCvUqdGApjPBazyWEGm1u5R/8ehkOAPe06p1Znl+aH/jEQxqkQxC
ko9rNVjwYz1JNgEGN3LbPhBv+6w7sh/5eurNS/ncN+P1Q7N0xIUI0QOfkzU++2GK
n6i1nH8xt/hQyBvlsJn72n9d962jzxd9BS3SkcrW36O5glXYZgpkT7XniqccEWLv
iyvzhxwvUVsPOFTUeGjZZ3j5PlLoesG84qfY51xzvj2tVTtn6kIxo/RSYss98iLI
9cT2YqX3oGVbngbGyLdAN/zh32wOen8W2ibhfEOdO2HxBSClsqZoS4FIs9NuoFt5
1QFkpNzVDMT7GZBzXe5IdbIS3FTmgoE/y7nm7avi/ETsdH5Wp16hABxrjKORHFN8
4WEeR29lMAgvD7fWUjKJW64akf7VLDeavtHMaEaP4l9j07DY3WzEtggybeLqYWdp
tYO3Od4SeHFTdIRXU6kfmAnufoFuX2vxDWLd5QEu7saEIv5yqjzixSUAyhXMDtdz
eXfuDW03WrKQXl73QxnbQvUjc21yZ/aepMuRXP91MyC6gP2WSu1fzWThI6s1G/bh
C2qB462s+57CIcrUuX+MIOM+JRQ3IxenQx8SE2D0B0E3LJDFrUgZjT6EBh5AV1XU
SwvNpT9bULtvFukgOu4HxFTXcA7DNdbOxkCq7MWbkbcQpVS0BcBNBxWD9CgaK2YE
/9JCQ0bM00lqBd0qiD+jlBRJB9brMF8NYifq+vC/RxANHUV9wxzvLvxa9AGT8J4K
hbAQM0GoQNLEsbtMQE3w2ljNB75ThakS/Kc38tkfKdvknvOG1MkxcBvQeHt9X221
5A7q/g+0EJYjX+HGe4S5FJIIZedZs4K4+jiPvaYcqAej6RC9hzzqbs5++TAF9wi6
zoF0vu0Mi09m0n6C3GtWwq0XR+cAw8f8ceNtXRqLpCM4D6M8flFj9HULqO4/Uk4G
xuoIzOCxmALcgldpmu93p7sUFLnoBn1GtIpKeDWY0hrgq5qLryzobqJiE7laH1sK
e7sPr4b6DBC9LqnHoJitZ3EXK8z9IeWuM6QKh1JYY8+nnLH+7poy7NtFjf2bJ/Rl
tyKgvUPQG2AiXec6ZZgvviLTW6vtNBw3HGBKpG7YWlJgsSvpSJ3nT5f9l6egQR2e
+sSG+5F/lE8iP1rWgkG+FQ2fzCGhJS5b/d9zQ3wt3d5CkqL1NmUIadP2osKl7K/v
EUR3AzdI4v7SiOciWKZ1+WyoyCeLClQ9FELsB7I8372gkpVh2ZmKrGyd0hFygebL
2/9BOCM2DZBBZ3By2IuOaryq8L/E9LuPWbhbGQT/k8Exr6K+H+P59FCyaXEzE6WP
rmpFtTui5hPeDraPbND4ElxuQhpYP9R0BnCav72j+t1zL/DJlwg44XIDcVHNdPiG
vG8sgfH0TnTkKusOIrAUskfCiXU3ee7Asshn+F76V5sWikCF5sW7ktXe+xwY+i87
/R2HC7DiIqZp5MH0bpsdtSmWho6ljK2aNMlbvFkkTpkM5xkGp+HDrMMKX5+mAi55
u9sh90y+Q2hBZH2c/5r2183EQ9XO/5icWg9TGy4Cv4niNbH5MQf5EdABsOfAhjqK
VNODjwJ16zV2ymbKvKE2JWM2pX2s48+LZZEWhtDclwR5WO0K4o2VUoOhbEhIGRKz
zZ+2dZtMI5iRxy3D2eFMQeqVEcHi6mSMF+3/dDxfBNHr1D6JSgKHN34+2bkD+Woi
+c2yFGzS/IrN51cHSHWid3A2E2anEt9qaF+oODKi4roNrCrktuvmo2J9VSzIZ10x
4357CCDorPKH4lOiskiRyAPGQIMr2WpRdCTKxCDQ96sBia6119sbW08dxq1wxZ02
vYPQzo1zxJEGi39N7MojkOwiB+On2XcPKUKgPHSwCNWnbEr1glDla73jW4s0Yih8
NWQCF9W4C75yQnKeU4AiL9CHsO8ZkyA4fPQ1NX8aBxsoJDfjObvLyb5WB6zSOElZ
j4huB/IISbGYo4nKFa+k0QTNE9rKlvkGvaiNa5/7+c3Kg6262QnHqevGiRuUdpx9
V+DlTKWHgtmPpP7ydibFKx8aj59OKqlo8gaKc4L5m0uZ//tfBsJqMRLxz7pLAT9C
KI1qyAmktDqaa6ckjxCesvRGeOvSjKBz/pNBrGMSUjIRQUlvlBrXFi0EmOcCsJVM
rWY+Cm4YVFobRl62tZjiDfJIIXiGq4vnfHjB5Nd1TatItDxOOZNeYhJObcpDQ3e9
9VNdqK+KKSsQjMUTCdD28QFHW6+vvDyJYg0Lld8dfWgpmCNM9chrIe2wzqzXVNFA
+yL78OncViqJ/1axHLoJHXb30nuTT6A3XLnau/ap0hXLf2SEJtcuNfioEIAFrMUX
Y3QhF7O3W4V9f8ILxmcJfLssg5Xc0UtjzseIX7Nlp5cRnbWxVN2kG6t5wVX4Pazl
c62/MACNz0xfcaiEVIGd53F9TQFC+NLIba0aVm3t2YC2KmP2iwgTX7Zd5hFFKo+t
tcRXXaZhdY+hVc6vnj+WArBYAkHkkOw+EGI6QsjiipEtlGB9RMsXm9qKADZ+RMSL
gg5lpvxm/bVR1gZCnatUh27OkiqlafSFIR9Sh9t+PtBkWqQ0xMmSMsbVyUp5WGmt
96c4GX+2Y2zdcrXD0C88nt9rahxanBpxMXuAAvpOmUxWaul//1L8ry5o9dkelKMo
8KNtIb7l/Nxn0YGSKQm5munSSAG+qux6WpnNa3/Hoe/mwx8oki9AvwuH4AUjPPsP
CSkq2idCbtv/6DiHzU6NkKtPGvkx/VNdrGN9Bv9yYx4DKELBUfAl6dVwXRSf5LiH
9apOS6Q/WuaKi8e6gj47mAycA7TwVEYNA+SaYPd7piP5hEqszwsKqHfqXDQbYN0h
Tpnh0QuI1/jwd5zk68pjf+5P4bOgMDJEok6jkm26ES+bBTED7sQn2oYHdmUNBD6z
ZVirmcWKzN8arAii3pkb0AvfdLT41tUE6MUq3S0+hshzSxEafOSYUSZVswDwMoOJ
hJ3p6Ab3pzN8WYNXkXxX0onSDRmItTUNNZy4dfEmjgiyv3shbkLMfNx1uZ4mFfSZ
1gLSCb6wC38/wBRHWOSiQdMxbvkUoeeTuzl0RVeLt8VduPyMlWXVKSXbD7aFhC9n
Ku6TDtaTrTMP/q352pKYLpJicajT7pw9794/bbcaEK8gysMZt0i+micIaj6T7eCl
eWr2WyITAtmoTai+UrRb70Xn/VPOWWnYUvivc5QcyL0n2M1DUFS1WvCsWRQrKBDu
9e+mZGgtn3pMFkpu41nntu+Zw1HUkbDKvVDpNy9vWoq6Tyej/WFUrz4o7piGV7kh
mhfv+KGjaCtdFmncLI6H+5aFN0iFsVOq+wy0Kx+72n0N9exTLMB7uE1cqhTGmrfT
rZ/T4aiCiVEgpKQgO8WloAo+FO4+XUzn+8mRRLGHMYepL9mH1jyuTcxxhEmUQoxQ
agL78bYK+/C8KLDJEjtcnMB13wEmt3nEkEko6cgK5DpQZWXjXCv/gkMuAPsncTOc
OPrFKI6PFOhYqbFHhMuo1iwaS63Ah1u3pBR6I+/ndBrLpqSwjH7dCZ0LLtKAs/LP
Jw3WHh355oh+79Lac4EV+17nEVHUY3SGxytK1nTBR8/SsccyH2EAAwd9rqTlozGP
DxomP0s26jvJ6ObsdHJFPe2Ir64uDM0niFs0PqsQk3XC4te4vusY9PFMQkIvnlSv
wJXkMMD7HNL2ZwtnO1PnIm0fSB0jhdAi1DWswIhjWC/jCXklv5HjaZjKTEpGJVs+
J0qYwIWD0DFCnd08AGQ+KLE0r8E8Ywxj88B742Vqka8ERAYiz5CyVAUR5Fse1VTE
4eV1dDwPZiFzLdAAgyPS7uRzuBgEeRoLZ0vtAWltKeKrC1Ejp0nsshwkd9+LJymf
q/pOCxZ2sJCoSJaEDSfp0lHKUzM58wGAAQKk79NEf3D0kvN4ScA3dVlozN2P01Jd
bqnRTgitf9XxWAAZVFgyUN9uJfJ5p3wSj6EEmQLVBrbQk6i0Z0VDWleZ/jZCIDiM
khVLO1nn5Q972B3+a03MJm4hdas2KsQZJp/Cju7QQLxz7gEqaVsCsZFlKUhv9MNY
TAU0R1RwzZpxebaEZx58d2EXw6Cq+dhiNkSj0gCWRI3NctaZ4szaMQMg4ZjRaMcX
2iUlQQIdaS2ubIya5IeDNC6FFoOKFY6+lSw7YlRxQICNHprb6XHTj4TKAmFeYLba
M0eA2u1+FUEmYLsQBca55UfC7YtldZzp3Pgq0hj/mo1xMRLuuTayBoQiAo1GAtqg
aXPVv165rc/wg18jJR14Nfxm7qnabIXqDX9Lajl6DTTUJ0/8chubtCszr8s/ofdQ
qre7OsnahgPe/nD4+Bv+UGqGUAWHeF+iDx+gC3yKh/UTgXJfJ+WAzlVU3HAoeFJ+
h23OoT3C+KqljUOe7aWVHy0OqiUb9F9WdSvpEIMuwUHV545aiPDo/5HTDg1zfzK5
9UvhEnurr1QApGzurO8AeyluiQpmj8bVoqGlEtuEZU+0Ro9zdmmuQrRBGc3dehfd
hgv0Ty3HZhRtRJ9F+oqaQNG1zmpTiprU0W3sZVHTs94V6yhpLZiTjaAEggF3nUbC
iqS9lpNc58mMGjdd5Nks8NbYfm7AUj798tqi4zrXkx/YOGCbf26mSCmXufKASDUH
JctFcgaZep+F0+w/jr0Nmz2Yvj3nv6nOwpTZngEZyLj2GgffxS1F1nKiE+2++uRV
7W+V7l2GnisRwg9pFhNXXN1lbKnEZb9V2Srp8WrPaFBmyBjpneqhpx9tCJLBGxwP
+V5KRQYHYSncMzPxr6aGS20nbWG1j62wZ/yu82wJp1tZPcsCS1yFgG/FmRfE2iJc
HLg38MEZEBrdseqNazkZjzTHEXJWK4avzDBtdSk0Exq8+iVVaIQl/NTKS5p8bPlk
DVmwindm60hQv5Q1015e+W+LTWT1OkkEO7ZIKoRKfkedEsKKZTldyp+u0Cyl3d7A
BNU/QNHKVWaDgH9c+0Rb6YKoHiFCkCilAh2M0R9xwj18OEW5Cnn3+l8Jqdb0aFqX
nf004sDqlD3vNx5FZ2k+nK5q4NdvhbNrxceXM/wDvi7oUHhZnuaT/Ah5SLjz0KQh
5WoFvPhzmBSnuqACtG1Mriyp9n0arDa2kx1+sHN/6wBMNZ6DFiTR59V+FXFyPhoJ
5t2iisbUt9PdAMPiRODA6POOX94OWQuDIX4PVWM8vd2oi8r9RK37LFA29a28QE5U
Iym/pjYBztm7fYN1MUNWc3cF/CRjiwkRQvRjccl5u/elYS4XbbQB/c7QFoypRUbe
Zsij5xhNO1CnohCUn0SRaI9Dayh/eyE5XFjNijYpdXWSKAwWIF208hS1WKkUQfNo
L071gSER6sOpxiQADWORZ6zweIZF7ad57Fkw/gPhTtLKNpb9KEADBJnRdG9LoVyn
RPXWzWiTwzUYiXvRA2vGxZTC15bLXIQl4VPzVNGTaYkSKnCudJOw8Yx+NM7MV6OI
hcA+VikZFtcn77/qaY/D4nsDzEcr5VsF8s6SS31Uc5bVrHpLtIM2I6DkICCO55uo
d19Gi9AneT5xj3cAL4WBT9SWWir0duPAP9mcAyAjDkozixe7PUPYdMM8CqZpgd38
GV3ZUWwArsr/OpLz3AhCMNO+QY1CZhRZokQ3pzcgfluoxpMV+6G/woksm232PljC
KVxWAdCRohr/+FXhZaoCZ3cVLvfURmt8jyZilsUb5IscKDSX5wJo3cryR8UyHeTi
OrESabKLSYI3eir4NUj/fUAHOmPxYtEyGFWSa05Tsvjyhk8kcdTlCWAi1zun4ukX
Rl8TLIjP6rVJTYeC1Tejbbc3ZCJj0wZP9Xfu2c0+u+rkL5BM4Nap9d8/MRpLvE7e
soe2kPy7v1+IiXPkxMXgTjJi68yPhF3SDdtJnYpHWiubvE3GwlVDw4RfNUcW1S2i
XWS3AAS62T4wt8eDma/ycv9M253yIPQZcaGZUyhGlVV/w0XuwLrDj64/qUCZGl2p
hSc2luWmZzRoEdsHZkOheYk8BlSN0yiO3eXRyFMvJMYhM0uDtc4+JI8Dxw+yYt1X
28sJzAdcfJETzqgrq/4E+6Zl5uYxChOQJNJyNnydTozuWT1YUeA0CeiGauXUFC0N
pzNqjSBFaGb3L2+cBdDOcszMuZdbxDP+62sxSp/9uPLtAUcA2mYvRZgzMFCw9Eoi
OqPKFB6pwK/sxufmsnLtAtXgyYzfAoOVs22czlVYkp0xZj6RWYAuN287j2MaPf84
9bpeISrsS6y7YuZWIJA8AVxO7AMWaw5XG62+QohCib/DrrmUszP6PHbJj/ytJTKM
ZfodrWh8ctS75TYthgb9U3BQmIlxB/FlUU84CqzhilkuBRrC9r2QMzkTrwGriq+j
8K1/q/bbaRhq7FWzEtetI26+O6pLHaN72XXpWAupFlmUQNVp8kFAHGt05x7I+Dr1
9wm++alyDh6tKg8rbW3jC4w5ewA7NVMAxOTRNVCm3dZkfJCZw/ce0TanbRrTidSG
IocEIMbX5vC1wX2lGOgaaHTMAbEw3tfo1/7M7Vcs/Yd71MbS7C7Sdx5YWamsVAHj
S2vDlx3PU6FEw1Xo/WbmxQELl7P9MDFSpKF6Pjt2gXZV8JOdeXPRcL0xpYkbBjNy
blni1HqhEOTIaDmqDeTFNt3scbZhsTAVQNqvjiyc8ILh2QWB/XEsoElBG2nRiBb7
BFAirmPu4A6NlluoapaKXG87koqbn3dUYzUeKE+4E+WKCtOoxN3GeZNX0EqRWHkE
0r9HsbMim+mjdAipDpWtlluZVTMu1c+b6HtNf3Up5ieic4hEE+IYmGoYQVEMgUYo
sTVf1jPFYdmpPYe0ZbZLs8kRlQLeJxkFdwzbiApXvxdQZcUz9poHSmWbqVsqdSce
4JbaaY6rFt9Bq+YZVB2GVTKFLUuWH+7YnVbw46vKYXwkRXvWbY8kb9R/4i0DwnFI
OZDwlNfi4NAT3ZCaKMqCFpbtopmK8xf50BPxEoHpTxjszsQHC9R6xN6eQeNACrSF
qu4/0VchQ9Ax/+VkGrzzoVOgIM9SCExDyWjm0xzpImkxY24u6ysxty4FccbZoBCT
NaqbFS+C2irG/VHwu7VsN70+QV09SxntCcBU9fQpeZCl2RBB3rxBAMXbE5Y21t/h
ICmbLmtZXvLsAVN1fYtq+AeEvd/qdnlR9pIm/ao2MKHwZMVL/rWuqf6P4nh6IC4K
IMOJ1uXEjwscmTooSeykqacGrn8HcnoEpCJqcR/40hDSgnEZPdd/RXPVLHPvYMbx
PwJ7RRMs+PID+eZL+dqR1f4cGQFGM9WIU8rFaLQZX1A35RUOXRt7II+9gVmPJ2w+
w3dW8L7mLBfJM4Qj8A3EnxZXjTN0RtOOXIQ2bOacIIU2tU29pj+hTFJYa8Agzekk
qtTCx+H2JgjeMQw91s3x0UCvWy4SYUPNMEtcTARmdzaqXVkWsfg45CAH6/IOHiqG
qKoH60plkLONJ/Dafmw5aVu972AW8X8LogydmRaf/zTLTSbsK71YzswEh1wvkGuj
vgQGQk5kW/VV/Vc6/NKHKAqNzfm0KOpslvSFUK3rsvSDimgEVVfM6wXCHl5xboQ9
XZVo4/l66loicjL4VLiKn5QBag5yA2khola4HYXaGZnftlNuZr4b3bqtVCff1g+l
EtXGx25ybVJBcsrwSUpAy3AHfKTEn1/CV/ZbGgV4LlJB3Hu3Use7+duEWIayczw3
XVst+vrZ/35YFON0R+T1dm8So+euxvH3w9kZ2Eev1bRVOZwydlKyNhGM5BX8scmf
p4pvc0rT0mcg21JZyZYytcCxDJoecgzDpD6ngl6pVqcK0Tz6ZXxpo2RP57u252v3
XNpCKuPZgniXCKoK8HeHP3xmwRZ4AN/x3UJkMxkch75KNs9jiFGx7G/bX9aXyujm
zRS6Hk9jPSHGIofIw/J65OLBXDQiL9FSXA6daWxwoHZpyIg9Ishj6dX8aJpOHTyb
woONITjjof/Dt58a5ufp+AvVDxnUXQ3j4b7ryQBiLtuBEYFqhAnIQUC3LXBd27/g
6x+QM0mDwMyi05NYFd/A6ubEF1WZb/n82D9tEPUyVdlZO5GlbxKItUmbFYDlE9fy
4D/0Aep9s69B/j0Gm6vq4vW1jGJEOW1Z3fVif4qcFSLaMIcFLCA7NRAaWN02ZyTv
zDSs8kJF7NWizWka4WQXNFaa9APgd8ysaxnr3C+2MUF8Zu01VFxTq35cQxF6nJDP
zHHRwaMHZXGVP7CU8D0ro6uzBlgWmS+sLFlhyosM1aCtRsjC/mDdYD8ej47jdKFV
U6rx6eAXTI2mCa8ecFYGEZzaWT+HEb2wAdbr3jMRIArUr3/EALGVpi9EpLltTG3p
KO3EamC1EjaNWF+cv1d8Faoa1pHbwRR73tuh6Sexskg4eAbZ3umukjr8EsUH11DY
GHDJSwmvGumkGlY+blpG86uwZE5ufMlzhvhCXUEVh1kp/SN93c7V2sobl9FvJvgC
mw84w3KEXtwbe6DtyLAWh5YcboCMkNao/fiUXBK3Lctrv5YEooBnO2Y0K+Q1Ijt2
KdhBB/2OHbVK/01hP70tGI2jlivFQswRUVjwhUhCYIIy9hDtgqT1bRdY2yD9fcvQ
j7xyUOuEBB9TjaeNxNBrratjOKmuOfb67Q0Ni7wI+pablfkTX4Qj64DqeLknAWhK
Qhi80UAa6vldJg0uh0WT8gAiqmiLOl6f+lGj5qhgtXLLCUanN1zjoMx6pQp4FxIC
RFo5C0VmlRZpwo+Cg29nL9kQzu/cAyxt69AOsd3vJn8+FRMhg0l3lGHpk/tCHkuc
Sg1SLCuRJoU/bCVAkULsKnULYL4JhfuyCmz6Mdui7oKgHN3vm6KJUNMQeuA2ZqR5
7pdtdLkgiExCdB4GTGBL1ujBA5qK9QJtx3AlaBJDUPMv3EGoBan31d5Pw0lqSAqu
t5Af2MNw6Jzp9Zyn8LwXSdzD6gor0vTlPtkRGdWR2y1Gt6ZpKK6Ol0EXie32bkzy
Bnzz1qAmQ9vH79QASm4NyKQ2IlDCdaX39AYQEK5OUK8Lpmaru82/RrJCfeOGZu8g
PaxZX5CxMJkV5VkkHVWBnrSeEGNLeCeSUEwo230aoPXJ6QFYNAsBmWyYE5idDhn1
Ph7Nrw+abDuWWjrv25XPe4jiGkNHROcwdb2c7ikonU4O0r696YyP13CGD3eZLjsk
IUR8bJincRMi7A4nF46Qks3uFKv4eYLYE0hQo0K/dQbtPycr9ksUjFLkkAZ16QrW
/Nn5X0foFagMaYEeLUxuwuTG+RhE90LOEuYWpCfmOJLC9kJSZXH8N/cPDCXlKLra
7D9quj7/jHEHTJ9I8rg94jRzte4uAqf4eSLPI+mgRtxaaqHhFbuKKPDbImliYhW9
DcTW/te+ldUtv1S+ecoGd8ohG6ECPxEruIBiMmQbQ3oR+4kITsEdxAQck8X3lNS4
o6yR5aG6gzQCa7rF4/7zMDdWQ8cMcz/a0JlWt1az/cV/a/3TLgqXKHPVV4YbZjaG
ZKludO3nQKlZnRFyrQFbEHsoRHT5r6THrJwLm6CNQWV0ZgR/e2ukrJdo17vwmvpt
/EXjqIdM9VIcDuOfO4oDv4EFvNkA2WRq1vaiBwRWjx/3wT1ltCgR0cywIUEfMFFO
JT5TUAqlmVB2h/PZpJY9T4GlRiaN4kuIcMYlY0wpzOcbxCbIwTcX1R98+Rz0OjQi
MZ8Ms8cyqlTMqLFKPep4AbZkvQtWYZWDZSadfdgpjs1+ZKGcdq024wgO+hH22Hhi
mwpnsKqO9T29Qbq9JmsSLtkcrmvl4YOerEx+PeCNwkw84wJcAvlR74mKadxXyN+F
RSrqfrjmoE+fXLVO83x0tyVhl/GV63QDHD9GKr/37sHH1RPbg6UPmInvaU/umiF4
DocaIUuwHuWCWN8pnFGeEX1QvdosMBKVrwbrbOVxHUHgZtiRPYCOFAjcNIbEPz4c
JZHg2wX8jyK0h6EqEWhw+JlRJDqmDd6zTxy19T9aLvuNpVYyBah9rxmrrgdL3Kf1
xi2VZrKk0fWIpz5mNLaRSrNrtJ+JkrgTskZsQocNqgtNmpow6Oq83AP4xPh5ZAxR
e7nPq3M++hVnO1Cpt/EWrHB1cBLPs2HXgjE3ZrUHKT6KJ84win1IpoYKEiY4iKj7
lc8t1/YcSy6gVUEAt7vKB6p18zNTXyhzZH4ihdkcwRXuFqs+fztXH4+NODGH6fYj
gLhu3DQpOztuU7h7n1tTKaXJ3FCgpCBbnSqD+5SescD6x9rv5ljREec7qfgfRbfD
2Sg2iR7HbFU62POUTHhDhdN2kqWNDJkKNgK2j2JfwtFoSpGe5lxRbcy1ErC4Aqv3
viI9jUtY1WMSKMnNkb7E1aRWbnyqx6xJABbOnR1am4ANTIDMfoCDQBdiv8poXDyA
fd25sUX9vwQGeBPM+kocFSRonGJ/JfvzmeGWUaWFcA4J3sGl0dMfYoQZY7VWXsnX
iU72o57Lup7N3S0yBj60pTCF7KncqolMQokLH35fEiK7N+XsZSh8XgkRNXZ4Rfi3
AsrRHmnec2vq6tSZmkViIUeOgJC8TAltXnZEIovv1NQnCDF1Djey06xmf98GOuJ/
jMNrYPlI7U75efEXrKVVAFESYI6Op6/QvhW5xuFFy/MuafBUVdYpyMf+QLiRFAVQ
3vIBCg7u/YCM6rCsODe4ZBSqCiHH2iiznmM4zjIlItT73nrPQioXdIv0PvfC5JJB
qDWzNDV+D4SectHkzF98knXbr0f2JhmCgc3YC4Q3/jMVeP+j2s211mhkO08zVMhm
XHgVpQeSIFqSBi9gjPDspiUqWkAR0DmA5a19yxgyQpxMPzElfOuTedL2ZPBkcP+y
N3TYCj6JYnRqkSROaejSM65T2wySgGF9QZqeII5Yo7tmFI5PF9KSfkSC/tViIk4E
CxCpaJEyXlsWJEyLiSGDAXjSPb3oE8XxFTAUv9CZj6MH/Nt/UIpY35nEzzzhyXQD
Q3tZncjtrF0ggYTAQj3JWDiq3IgA+EzOXTJwz1hgp4mJjjimNln/W28DiBEibUK3
0iAh4utHgXWu5sfYDKFD+7ovFKeqQ18iFxrGsPr67yLiMaomfg3nIuSDCN1VfTLr
JzWsLAjOSndKD84Q/GLWFYqfSx3gyEeUzz6K0zbSt0VIMWR7vJjRhOYTwtdm98Bj
3AwLZSpoQ1k9r8Y8aSd3vvHDd/yHVaP5mfp2jZtRvMdc77FYqR48BM0e9VDBGBgI
DQ2lLjnPdRMYqgL8Lf9Ff7qBq/CG2MubTCMZzJV/exaSOeN9/CFEQza7FVvm211a
leGY0eDbd3dBLjFm3qua6y4Ixb3Zu+AeY8igHJAKKSFIhTAh2PJCiaTwWZDD+BO/
Ej2ej8ro2y9ty5/n+qE+lE6GZTgwZIzesGzbkBjdTeYlHeKVpIXcbWEZwuB0jCLE
vfP/hBdTx8P/Hy0Umq/Sv00j1RAnjyX/FJkd8yTL3obuVf0vov2lxtfH9E2wg/l3
duCsQ2BoN8qdqK5Ri0GNNl3+BycELXNENE9zBxwS3D72VLnpDeGNlwxXYMwrdY1p
eZZ7mxKvOIa+3YF7bO14olOenRaieZ/xnOF/5DK+MWeRLNfBk1wQZkMRbJ80ABs+
kuGJ0c9jS3+s2fvk+uyvOBk7UHIF/QPqn6YPwyETQmZlDemQTbrtL+7A+xzgWZTB
8DJj45A1TAHmS8ne0XDTsQwxWjqTVQ3SLrKDwn09VfswI3dsyYC91uXYvupLhX4x
PTNGSNguGpbpip4ehJPrsxuiU6CbsUJUEFbVM8BsLShAJDIC4NRZcZqhE0gRLLh2
lDWKDXI5ov+PIPKBh5IAmqVnThbCbM3RNIYOO4k/LWYm8WDWnYviruSQjE3qSP4F
7IeWjFjYUTLV8BDy+HW2Z6Qv6eAkswKsQpkGlQlwBaSOktG6BU1lejff7MdR6NMd
DyGx3EE6fJBU2A1HmiTl36CUURrFkWMFCbOjU/7by6R3ltGq+CXOT/wEltaqNsyg
hxWw8CEKPNwU+pTEtn2cUO25QPlaLciY1u7uKuC5cHNiZ2f81pyLWtm+SopOumjJ
hjGVipXMFhUrizLB9a2i/fNnanXIOc8+UzryF3YRRnAoQOA1SK5ZtgfiLcMtkxp3
HyAlbJie1jPyNwFAGAB+4/RJ6xuV3UTD/+jYMWgs6LQj8+oJNfCk5FqhUv3Fs2OE
oKE3dSh9TM+lzVf/VXeDOVFDkaR2UkUpg11C05hixjiA8nqV8XraPimJegbAeF7+
Hjj9EWkjxO7CbNvof1mm8gsmMPIYA5eUZ7YywzuDJdvmLBAwsHjk7vmdg9gaqcbz
lzfHyIUoTRH94A9Xx62CAhw9nfDCz5kiNWmnlZnetbXfIQVFvf5xGkJCLMGFvgLv
BzdgTDelmmTCaXyUjyKngG9tRUqCN5b+fQ//uIlyssexj04s9L15W2yA2u0VUSVH
wIR0FeuEmTh+tK9C8ak6f0KxJGk1UhIG91qS/ms+27gRMnPRv9oNBDzgIFzZtw7p
9PqiU5wC7i7FkejzdScdpvt9CXGFv96DErC1hamo0jSPzOUnb5rxLbsEdEdzv3H6
bWWp+125qFoXHszXldi6dn26vqtbZNzV0+VHlQ6pK4bO29ES8TIiGtw4VK0muhRx
7rXjbnw+yz8nRRceJBoW+mD4a8L6FiOpkjgspnVE61WOzsUpWgnokDo21u6jqX6m
+Gvyt1CjoP/bfHrixI6KnGDs77SGrj0QfM4hcqTY9Ilz4vJyoUqbuZSyeadvRZEh
FrSO+HClNvXELQy2+tLrJDl88RzFN0fGv0RnCpdrssQ5HXdhddCZ7E2f9M+9JJ38
hp6QuzihPzBWvITHpCdbJ4KJZLZr3DqQ370yLSplI6IE72n+gnOVDzOUylu0y2Ib
PGua2AcH5HOLZP9nWi2n3oIYmmAccQLL2Iv0oqjwGUWqrJs/LMJoYP61cWm637/S
UiV2tsdMhPQ9CT4OWeaz1bh0lPvGhDvWfKp+Ipkm1kATJCVwICSPXamfLRcUEOTc
DDjlo721hd2uWppDvVXQtCfumavNKQxI29c4Z9uliOjMiMl1WSg2tWBugLXj4eop
1e0w5k4A1WET+DOzVlnBev9f4vPS5bKGUJzYBdFPn8uIAVsNrt9BXWqPIjkUCts6
cVjPqW/Kd/A5wsgRjDkiOYpekIuiiiF7z9rQlPZG9p5/W504Lrohaxso/ntV8Y8E
NgJ4x8134lgOj5I1XNtKtCTZIEu+7uovzByu8AVg8ax1NFnxM6csoESrqsIMfZzj
m448ZMlAZIr3yrpfBTYNDdO1ekt2w1rW7gNIhRgFB0YNuCF3Yh7YVN7Fbdo1UdPz
PlsxJFBHQp/XWz99gjjKj3dMZmr9EYjBgqhdZ17NwrmD10UFrQYfw4kET+eoVbhi
7x6Wb/0SPwjnuL3ymEZi7un1ybKYXGO+ngu0VU1mRoY2uUjz5peuzXOGsl57mEUt
+o2k1cAIIPRG2VwKPxIlhlmNS+vGTL7Ek1eyBoJZHmqs2Z8FsvZvN410xCcvk3ck
wnHP7wlVqyqPCUPRfdRuBGAfN2SkI4GFVAS9V17VI2d1WyFfCxoJ8Jv8kQx0ub/F
e37fpPxVW/lCrKqxznT97Wiec6hkRRCKViipHHmEkjR+vuVyzJVnFFh6r6ML+OlD
lEgQV421q9Uq67olj2z4kXVBLNW0smUrSlEZ3g5uau41rk3PX1HQBccg+ifCqV2L
LcdqPE4FNHW3VT5J4K3XT98qzbqGuz4l9Nk2MQO4qtjPeBK5HYrwGShKKMzueGk4
Tzp4RSO40pKrKkbty63eyRAbT5OE9Nzib7hUPKK//ncFV2Qw3jFkVg8rmi6iSjfY
ptNixmM4oMd1g3fjbiw3MeJVcOhPxKOGHiEm7VOf2aJXbh954DvVz22yhVgNsER4
US77rgiKxip+qbQaLvcv5TWD0uX5LSfFGMWj/UPiCyTBx1HWR/vp2KD+veYFqQvu
R8mI28zNQtE7LAf4McMRoLAwXKCRv5pMvYQXHDQ+lKzskqN+pjKhcfcf8IMC3XPc
g9WkJhckg1oc2nO/3j+jqeXLd6/lfAczFtAjrxsW+EWTcLieyi7+RWtup82ZykTw
LViYArW/4IavaSg6r9qr5+sJXCYlOdv4HMrsMtmYljG0CpB0d7ziNV3mFlo0J/K3
0/F8ai8yEo+Q0j+w1YKjVdGzeaozKVna7Xn3vTwHWcbhddhCJeTl4hlakV/PxMFy
9U8nV3NdQVoQz2ogjgPkxRvPdTBVBiEFYgUwKetUdCeMV4vq7CAGhn8db0nLn96Y
zID9af4gpL9AJklhG241q20WSvJOLKeGWaeMsfvgT2KfwbpE6JsSwbhH0XIdSXYS
c2VEncZPaRqhfgiKDLG0cThpD5cG34wuJVOqUjESN2mOyY1vOhdYzwxHxUwZwlk2
EiZEhMFYcIviIjv5zssc+ldBsRiqN48Vd13sIUHIW9cC9c+SWwC/TGswbfbR0zsK
YH1mQ/sAouyxhQprdxX4S0eJ/euTROjDq9rHfaJRaF8Yk6uahPyE0k+5RnNiE5ww
pKuhCLqGHtXsJTFDEQjuyWyaU5G5Hev7HqNZw0s/txMMwfj86PtPwjIqn3Qj8zBj
fjKIq2X+ISvye0n9dYSzi7kku1ymrGzce6kzVYJ3DR3Xs2jjd/9x/nUS+raJb0Pt
kRe7Stwz7QKy4s00ztmre7yFWXHAwM9blVR8VxdLmY5sTH5qxXUQDmalIoLdk6HK
azqUEqs4nLBZopCn9Vg2klMM76qYltRylJQUUU0U3ir9z13oHC7Lc5hQPm62JQwC
N64Bw97c9wDaVfkojQ6jBJE1JqBkuQ2Wk9A9jfWRlKJa7gc85PMm206sN9gwSfkn
pEPXbmhTzyGAmVOBxkzv9+4Vzul3jgKZtSbnfteHip/V+Xfh8KlJ5lQWzbGhPs66
marFvc4B/kXliekqTNCSyduc47F/w/vmv6cbx1BAKLsaXhFMekWdslg4dFy2PbPm
Oj9dFby31VW5E1yHFfcMHexh50B1tXpCPFuNHj6AJpLjBxSQA5dqQnNzu2uSd/Fr
BG3HGEMH5dt9d5BVrIcj3SbH46x3TYL+oG/SbKIk5bWArBYFzSQFmvCwqjQHnZdA
Db4SM7SrK/67iEDMqrvVdbFwYc/NmuGLZPaa5FrwpCysBQPRR1fGx9cNOsNjUnNB
iYPZIzc+PId7GXKwZAXvWMUw2L5bQO0Ulh9mm0J7hfzzTSeWidsQKgU52PmGezlv
IOXRAEL8F4UeHg5plhNQTe3yCBZaGzOpXHaHhMtjM/HOAn7ntqPdBAa1XHGgWT5g
QAidu7pY3LfsyooLFo0JlZAvMS84rm/6CW5MWRs2gz9VugVr5Q2Ly0mI85ger/rY
5HtYi1MS3QxSmT+M7LydV+AQ1vT9a+sOHQKxrIjzcbEk1vZNcCgIDF+tDgneqC+5
cM7Z2PA1jz62G61pG/Zay/q47MCQLYKY0lfD2hLgI+zyNJ4lUgJTli2FigLaSUsg
nt59Yy6pE/bhc+q3r5gvRKO2WzGa4G3uI5PUDoOCQ56Zs5jRKqZhrmgGjZcTHmo8
MMKYRpvaJ9EBBd+Vk4+FSS4Mm8jleicZ8jpnha+B5MBVi7a+ws3fblPf9UTTYvuA
OCMu0IM7hkilBksv7k4yEgqGRxi/3b/0fRdF/1UijkK2/TieQD0Yh00farMT8tMn
P8CbYPnaFgWOfChvtfnyik0nEGZrO1v+omBZNvsPvaIopvm1ptCgfhjl82DAVGY5
DyMHDte+uHxkO1JCNkxiOHu0igRteDM6HXBj+CEAeNQmi7qctJG/EDEzEaPh/D/C
qPesGqkZ12ItSD3t4ygYFa22nOGvi/b1BIU0qSbWzR7eU01e7+lv5g8QC0c9gUYP
/McnenQ/YpC0L+2Nv6zvF+zeyv3ux7IZQySNc2o7Wcu8IkFgwqO+4yHvT2lD823P
Uo4YctXhaJbE7i+kEV/L2yxfVyvavRIaBLREFxiQK5X/ZMlbmks6eY90XIsRJSvh
vHFFNvjgZ6DpwHNikF5IsnlWBQ6SP/U6yiVi9FFSZzzujdjl0OmQdnjFSjYEq1qD
U0gWSRoJ9B/oIAVVY4GOtt+95EaTvM3ZEkQrNlQzO5A6hPG2EAyhUsPOKgEPxrZJ
VCABreVbjVyCWURxXCRpDfXjyAm35d7JyAEX5XnCqXb9jVFLqOzMZt9SsOuQ9D38
iDFncfQax7PIqbz3dFsG8mNBOFWuvtQ14e80BYD8MFoWzX+EHZr3YStZO+fuWtV/
ds0JS5HcOsdNIvggxlMHYQNkRP8YVFrNi2FKEiM0nHnHs39L7PO5aPYkO6y8ALVq
XbWtKxIgC7w0OleXvf12AVBQGlZtI8VaIqYV1jdSeZdKnDD3FYtTH85xTKtpkkcI
p0f4I9hjy+dHP+CN0Pl4cNwyAhMDPGEqYRs9IAgf55Br0PxuItPM3EulV95QF6c8
RM6iWmegOm6b8mwFiX14g4WjmUH0fEdY1h3hvj8wQ8NLFMN358dXZahPENnQHd+0
Ab2+3o3M/0UkQ0lr5cpK8qbeNL6Q6xVOP5Q0wjKogyBjzi2m3jFqdG50clmNW/zU
15QsC8KGa2MHgh08SufFvfAAaoKGfPud/dBuT7KmjP2Ngn1Q/ltspLiImQvAIZqY
k994Do3+mGEJVE1Si3JHu+D8L7UeTB8KC3L5runHHslgTw2w9t0N9+H0W1aCrwC9
l1jBsx6egUUbx6NXQdMvVxESD1WA6v6Vgy307n4jlkJMmX3bjAwAFnDei0IJQiia
j9bYHk1M+CIa8199CQ75d5Cm387dOD4JiHtpL31icM7c/6uMSllofHVyDtlwZ5hO
5xLdUQ5s0+LCcTXe4VbrW314DqknMqzR6SawIP0+HLZ6Q54DKhceJ5MWcvO/gunr
YIvAG1PLmdVfKIyJksLEN1ED0a60QEALBNI9y0Z4Nz9KpvcXM2l31nPleuhvDaDJ
biqUPuvTmVpPS24lKfWSQtOPBeZMw6NiMNVqnLLm0qG7m8HcvEePgmY1kfofkdhK
2BO624BkycjmUbV1fF3LqIYn0B8iOv54xYdQXm7Li+pT1S0ki65etq2NqgxMz6Uf
ijZFiM/LwD2uDlyxPtQozb7tZlerixRIoaq97uwkoCtt+JUnCGqx6IGGOI6JZTNX
HDajKKvt5uu4QMXs1Z4kvDLFNaycdlcqArIVGVwiT0sjKbLymucRqTEryoJZJqCf
aohmUAslr+L/iCLaI85sKm4cB7OeojLkSheXKiz4ZK1HPV4rJ7Tst/aHupAa7cnX
t+RJJATlttT8ZWSueYF/afYc/EBf6TPJA7Eo48w27M3WsYDneaFw85B/Sn1GZawS
xkGBrwFm/HpB5zoDLIqNHXhafP721QI4uijq4/shtBB+B7/nCeFsfoWyyWgO1HHp
eC6AzE08Wr2bUkWLa7of4DDdmv4EogFvE/4wEx0MPdweqDczKamYkElHPfHuAgzn
a5x7Lo35zDqW4v2ijabZD1TdCdMDsy3NGkQyAUZyrGoRXlERQUXmntNKmZLegagx
rQuhcEkV791WjKeFsTwG5+PbwQvfoq/VbmTh/ngW6bJm7mBsmAbXlAlaaYvWS2gY
OZGtAXiHSpqo/nr0JehRnWhVU9H+VnMf+pJ3pjRXp4CbTDxBy0JElOv1fna7qW1c
nppzsxyUvP6C6eQh0egYKiENkMz+ABc1njTJJoCnfULWMN+TiqVi5LhntWCY1Jzh
Y3aFrl7xP7JB9yna4hl843sQpU7He4Z6Uu+b14GvmiXqt7Qa+L8woKObhWnuXeWo
UV/q1HVuBcKMdhHLTq/M72bV1p7enEZAQbPTA2oKNhSOwyiOZzp6WLQvjrBCb2J5
SS2yMawaJ1JMsbMnh3YeEF3AvwTwDE9ShMNDXWadXlpz/Cvl5XNz5vXqPu9V9hCY
deya995sL8ysDNINTV1O6rOoq/WmeeI5C6XvI5hBvRtdkRTdDcENfQ/Sb5LuCcLz
kwMKmkcgCcIAeEWRaPUQdVN+jKEDBA7iHr6m31qD9SzdOki7jTDSraz0kp6ePM1Z
s1+niYveoyz6ENlB7wymWIPAwh8p5R1lbVHPkCzps6PFuA3RdVrpj0Ufy8j/wwX0
gKfEZ8dld0dRaqFH4VH4Q6REzW5szL6dpmXeixoqj16cuz6ySsvYMLVH23+lYTQh
HKVQyK2s4Hidkvm78ehBOntxMlvALIW+wBTPQbvKL5nzkuGR+praGlwwDf93M/Vv
6vZz7O8d5xb37jmB4eWA13c3CgX2O8pT2bhhWxWQUPTCM9vE+k8zbhqOx/AHcltu
gFqOC1SvR9WxbTb4/qreZteI70dkhqAK6YGQg6oNYP07K23NGms+WvONnXmBsU9l
2VuPvSe12JP9QMmUutYM9OzAr4xZTgR9yjwkdzLvKIDUTZwyMhqKyXPLVPj6QGW+
dJ3O1u/zWm/2/hTIrcn5VvxtKxJrX/Ils+EAbF8mFVrzjoWoPkJDJGeUp6MPjfI3
F8fPLpv/9FwJcTfxKAHlOEX/LJKT+3Q/vNk824K+VzFKwJNSm9lTNjTz+qVkZ6xu
fj6cNoIC+iAO/nC97PfOXtGBuBjAHWHrbHpIMRHCnnSuBGnm4kR+rodX1wj76vrx
+fzoZtPtaDzLPnY7bDeQsAOIsrg5T35GM2yv5U84LU9T6v80rsxSi/i7Bl+Or6+Y
2RYJOb1zzpc6R6lqBhG8xYzCxZzb95yuL6HQT/g9SrNaIA4XjOdCS6U3x00k322U
qZwTM8hPttcFw1h2AXiXgl4PkXAWEysE7D2WlTxWF0bCYUVmeiTPT7SFhf2xFRfD
hD/Z2FAyixz6ZdERZZZUp7QkvM4yfzW2bU9OB1S+XzgU1PA5IiwTuwyqkq0hrCn3
4+CDft0KlAV1fezylRQaD5MU0uWV1gUwn5qcegpJpki+qJRcMFUUoEqnuFcAs0NK
Nbu5OEM8pZoVZb+tx1kR7QLs3eUloFuipokJOSekbourwCZvqvy/DOJ7HVn/QoEW
ydGQ6mcBeu8raRKPX4K3cARhiBnfOCoOLmpUw0ZczoCelNcZp8XFyZewybNYBCsZ
uny7Aih/87MafDfAlEqAtu0AgpSff5cZVK3D6rcraWDlwpaKrACe2WuC/Wg+DxkI
AOGp8MQFq1+70aR+K0f61KkZ/MlB8J4KNXqGhfjw0b3F58Ch4EAfYmuuIdwlXQlJ
lL96o2aGMptjbsfW4SqpB1Et/Un0+qFMm3FY/J2TSLnHEbSSoETxV/AmhRSjcccZ
M0N8SwBZs3GuMYBTaO7Xr9pwGOmollRhSE/CNWNq/LLKhVOESBIwVjvV60PM/8R0
sQSe4RyDEh0OEnpuBvupcAexpotaOkTDq/RFJrYnrC0XgJbt3VQ/3xLO4l4CbsO+
hU6e6qR8A7Q9+gILHu66LhSMd9QxFGa/xTFNr0wqu+NzVs19d4IOQmSGxBcYRED0
Siz/vqpWq56SFcMIDnz1R53An5vMCqCGmyjXmcj+iZ0x9JkTfkWMApfYShqjxR23
IVV4+G7V6hEvB8DNlA9vNY5I84Ucwjug/kc2wDy2K0FP7H8G7BnjjZ6uHfwcFye8
N6XxBTCKV1GxoeVYwpojflVCVIi3BR03vKkQAxmK+A/VJ+6ASomHkamDxcMUA8DS
zQG2du5L1U2/0GFuLgPE4Pmmg7CmbAL75fxTgtg9hiNk/tuT86rsfQW3OHpGPh7F
v12g75lCwlPSyHDbgylKxhI+/cuqABob3lJSFHhCXdoaFtyDM8x6KzXMjLZf0UAi
A0PGgDH7XOgLunXP223+y6kn2yj9ONhYNZ5wBhSuk75/KD8IZjuOupADO+CNr/Oh
cqC/v7jV0eito8fF2iOs4CtjW4gR+IdfGr6Y/VUv7XTOQ2M5aJF5WRm+K4K4aFhq
534ORFNRkKrbkiAm9bQhziWte8JsiVhEa/4+wnY4DIMWGs8diJ0+NKpwLZ53VzRl
PwDCXH5Hh5E1OnC2zVZlO5b/7DUYVYXcvJGJ/sLrkdNQseKyNXnbMJHN5WMlmSPh
KhIt2L56yJCip36H8SrH76SJ+eEy1ZH4UuHEc+HJ8xdaf0G31AfJ/EhClBSJ6LMK
DlmtDG5xGVPNOE35I2bAbixkS+o0GA4PQos6Uw4L3UqyUtmQdKbUUYUJ9mLssZCg
SN85QPDTpi2vavi7qnrUhPDzVO9B6ufkp4/lhEbwKaNK53hXUym24EjW9oF+JvE5
3s0k10EnF9hw9hOiae0IFYSAQtCjjY2VDsUrIScuvB8QWwuXVSB+wjwbxtfwe9kZ
hjIOwZ2ig+lan1zIrRSWQm8oIUJY0paVX1rfNIkTPoMHD2zqHY5POBP0J8/S0be8
7g288Ir+plysRPd2xNzYJPGe73WhADzuOq8dATJ9BE4x+v/l0hylJrr85RcSOL7e
W+AHUYCELeYrKRF1BCe0oEPYAlid+e15H9Ws13/nzkUqF85cxKD2KW5VMBzk7n/s
YvFqdz68tqxjs5pmJ+swLTdtk3LNGLqfQ0ZcD09vY8Ep6riqJ+Fp+zp70FMeLv2V
6g+aF0juxD6hcHl38oSMPiWI7VDiKc/vwnAaO2X+RewpZT3yw21ON6ozJY8J4A3Z
zu8ioxOd3p26pjQjcoQ7UGj/ZewGLl2rk5DLQbS1mscHAut6VPtorrVhLdeavWtU
Bh0DQ2XxxWZilWK+0aOxwCAlSxS5dJpV24M5scgqCDZsh2Tol/bUFzd2z+DneePl
m9P/VcHNSZRlyYC67033SOfU2Z2sP7P6xGv/SMTeXA4nLm3wUXBTSwv1kFTloXJw
UuAtH2YH1qv4kvNO5+DyWkaJuDssDIgU9Q3futlXSCZ/P1BM8R90hInAjMxrJ71D
zQku4/9I50vpmh+Doik+XtZzetsZiScch04oAEnC7uA5MZBG3oa1S4ipv4ZV3alZ
xaAaWxNbdREEuj9amXQBQAIwREC/a4j2qxdVWsAGJQzOOagapjfyWXall4jHGOXl
eFZYyJFVp5dY41pFMMZnvgTbZC4ZW+fSu6k2/C1ZjlqVh5Lmem4Pa1gs2z0aTRAA
KyYBTchrBuiOPatAf7GgRqdruZ2z5rW0Y8xIA9QKz8P30xapztroJv1wydnqjmux
YbL5vDgVz/eBN5ww6PpoGp19Wu4QP3nPKfaFSAcA42C4a0lkRjx6ScLutNrxd8kk
/DI60HWjgYXgijWtnPXHybojD+kpJNmO/bTzCv3MIF+uYLkYfabrTKhYBk2hGVFa
4qq3NdIGs+WyMuZmHOiuKqOnv0Ua1Sdj1qAV9Owxjjn9aJnlc5dWqMxC/Csh79Ee
lAsSDQMvLjXLVKnbS4KhjHoO1QbhV2R9Fa3k66tkxrxmbSR8kGWu/YCEOH1FU4n1
k1NlcrfBrmJhxGx++WLjt2ty85SWAl9kmX3R86MAQdQPKJyrQ5/XrrNP/sc0wvaM
avTJnWuNXkEPSaJTnIUpllKYhsKF6puv6Xwwnvb7pPzUYL2jzZo8+XaEMxM4hFQB
0UrMS+1txCapxUDSl3FIDtpEui5Wg9NoTbaBdcLyuNU8IuIRT67O9vFokqTfGdEx
xiotAi7+moG0nAVejsLFQiEOY4HbmASuv/QieRGmk3Qwx8LW13CmyckH574TFIQd
S8rPUWeQBVJJZC4nTdM2gFT9SY2liKX3ewfV6OAPS0W+9WCF9SiHSqxXHYafa6Y5
6SIRkxsuh1RXD7joBOREM2rce1i18FuBaxLK5spEoAEQciTKc8HV7np0Y9Guq+1B
76KdMZbiXvMviDGusQaf39zroOHxfi9vjHyl6GIwlFY2LTDLy26SFf9szGFGjJrI
uDEtAObKB8spvQPff5c5JTEYEYDTq9thTS1D6UP/XwYER5pNPmsYBzJG2qWchTVg
ZZMh2qUenu01KtgxXm53a5SCd+a59sWgBRUChk5xQGn1n4/LR4qqta8DQs6fautq
7Qa2Kosorw456y85RXW7637TXmV3uU+Q+nAMRonoE6/9lpRjlt85uKbxTr24YjWp
Pki9LOaXqVUeOtAoOXIbuYZBUFSylNAAlIWrQ2f5xUHVF9DcoR/HyWTb4e90Uxrc
GR3FaJpoXn9Qyfe/6ctNQN1rG44Avvg9kHXIxYIIdF+wbOeEUNV995MmRtPyBNbI
ZbfqO9a3tPaZ7hfuFEpVUB8z4OoTTnPgwCkH1t87F788FjVRBTrWcsqgNFNOFxww
cQZ5zhiCL2UB9xQcKjnMpxovp7fKHFU8B4aHdKqD0PJQ+q41J6NoUVsi+AWM22eJ
ERlI1oPmNuj0woLnCkDV6HNBibYj2jPcICstO5U1hrHJbHZgMMwi3kPz9AgVF1CG
/4lHexEYQEgAc1vWGn6TjWwqfPUG1gwiolAcoOXZzJuKEPdpI7ejE0gl2sROCOvm
PqAli+sqcOsnl0a0xVUITiiKE3SAAlqckslfxG1JB8IRylL2VYbELBt6wSt7M7yY
V8ZXu+7uR78UgQVsJEG/9JksyZx6rgAoHxqJcgGOC+OViLPx/i0EwEDAEz+MxCio
D590B/7gAd9S7YKLkbqUrvcHq8AQYaC+KHRB257oSNokUspIPhQ4rhm+AoA+nXDm
J0U7yT6b7AN/3j5sl4p1X7nsCW7BHc5DTCDfq4xyavacwOdzOgrO+DvM2aGKhNEl
ZDwmZV1XbRTj8YVL3Cjc1IWZteod+m20UKHY6npvkbvNKBGEPuYo8l0Q510qiKBr
0lESmZu7Rps603EJdMivT51qznmmiRJOtgSN+4fMTb/4GFplXY4byS/Pfu3PdC57
pTAX3+r+WQA6wAEQEqYzuiUUVONUFIv0J84SOIA8zgdO7RsEBf8p9KlrDldZxlcG
XwsGMWZhtGQEy8kBLOMUHm/PSe/N2f2M2ZcvDq0lIIMUx1QA0t7XOCOxIPXQAm91
uxZXE1GfkclwPldDtuHTA2VThlKuOHlHPHfGQHWaT1UwNQLw0Nta99GWLOrbdIS/
xWA8KoD3L+iaOf8Vv8IE6TyA6fQQNkHWdaHH5/1NAlfOqsrrpEGLasI/MIUtL13T
J48u5YNBLA0xQNkjrRcNc7xxYc+O9uE2SF9+ZzrnUN4r2svr8Sv9FllYXB+epjoD
/IkINfIZCerfJP71z3JNPfMfj6C5FJVda3C8qoKc1g9O/MroD6TfoMhlUqlcBd8M
s7tBXAjNuEUBhKWoZAb4wT7qF+NOjQWjog+mVgoB8bTdxsi3X+Ng7WtOt4EX2AUi
L8VNlXjycwqKuaNBCSZlo+09QUv3FHeO1nzeIzCvvC6eoEWGadrvkMeqG7ca5GlG
N7PtiGpcTLdpyumz89+NTwk+PVqvEDgr2bVBWPrueR1lkzsBUx9fP/W/O4k5Lp1A
QX5GgthfF1585y0uhL24MzmuOeo0q72XJ821jSsimOB1HnzltfF1gLKwapNaOHIs
wU3V3YKWTtbLrhuLcsNy2fLJjuYQXVIdLajQfY9GKkkRTJbt0ktD/cNfl4y49SVI
/cGI49U9ADYeU/462kk6zK5RmGrdo2ylwySciU5vcnhSyrH+P7AZ3Pz1XBBu6bfs
hHwdglAdg1noYRHCDY2XKCc9Pb4mZvOUo2nMQaLYXMtRHGNRE+0pm46LohtVIHzN
SxxXBDUTB3PjUw9Sct8BFEk+VCxNYQmBMCQGcqrd1rayufTgcICg2yNAud+XP8Co
Ut59edpm3fwnWQPPvn2IpyhaBGoyRcAvq5ig/jRfMg7VGG2/zqY6GX+e4L93j/w0
esmven56PPrIWvAJGOez30tD7/dLLye6LmtvbAHK9kQ5DKXbd+rFro2Pj6br9xjY
//thJMIfV9+aXSU88WhT1xvGDURqllEC1IaRCeJdmdRJ4ZwFNRSBzg+cefq81Hh/
9isQgWfgXc1M9P96OzogotUzVRxy/Tb63QYWUit2imjM7rJzqGq+JC/MLWsypPmU
yMwoPYx59JvEJXDk3jSsNz3XySX9LQnraTDo/WU8mgImoJj0E/WmGLg++7+hn39K
Izd526u6XAUaNOlNvbkPRZMdVvTxiW3eYB4s4hpkdTIi5yvGy/w3W1t1uX5ZB+uu
dgYtntOH1Q+BgUwJKAbWElimDR2C9dCzH+iY7XAjKvrqOj0wRD814o/xZIdPiPQa
Rghvzt6yCh/R/W/aL/CC6NoVPEe6YYmDmA67EdO5m/GITATHOjNkGMBpRs+N/VLs
ZWxqVVQg/Y5tjauVDgFJBI55R+/V4sSnaBY+sQZZQujqHFN3BD1Iai6d2UOV3tMx
1mm8LGFI3z0tRHlazf9Nehif7k17lPN624eeexlNVM4fihk3bI45SYKuvxpJr2ID
N/poL8h7lOtbu0Y6ODEGlsdajKzYH85qJnGWm8Ugk34e5uRkn/lKsUBIr4Z3jx2+
RgA6ek63tST3XgdgG+4HmS0pdNCS5n1H1X7LC2y+btk9NMMJNPqg2tTzwYe+o0rA
6vOlzdhDz+4E9o2Zw4EjD1dBDyqFrrJ3YoXpQLjXjecj3wiX2FMg2/h39AnsQ+vd
q3uKAzip2MhGAMFfkU7JupRpXukXMxW7ZUnwICJfH3EwLei0yiZW4uDkKBwCw3fR
swdoSt+ce8lwoolR1Vd69aR12+FpcatWVT365VOPNzQLg7qz80cqBJdcGtNT61kv
Rqi7M0aWe+41UglanasjRsM/wn2RuwSWH2DmyVRvUNuHoFi9Nv0eNFrJLpeC8tJj
tLuZ9WJRZYercf/Vag21ej6mm4nzXdNL8Hos7loMraJ1wwKRoCybEBWCXKAN9Lu5
WZddGauw9ywoq7vMx3Y55C/nrU9fHt/3oRZ7qhc8HVEPRYuQZ5dfLWMHt7hOiTwV
cHz1ip8TioA5edi4eG1ao2IRN6wIKki/mPyaUE67Tx+hqELwIa52I7Cn0crhJPl6
C2MU8luOoJc63qaOYON/rBv7hTYzCtG72FgmEFhWg5TKm00wF5FHP/1TyvZfvj52
bimRKjQzgSr+OXse6iePNSrm0Ib1vxIuDfpY1QeClHuAM+EVVCGhtTM8arpNnl+w
/5C9MLnr12BNgUZT7E8DlN076gMDXipt5Ozn4wjGotnnxl0Gv0TiEJgFY5DAqlFh
iJ0HalxOp4Mf0jJWZzeCDgkHyZbT4qG83Lx7IH+O7drpMhRi+xoVwJDNWCh5+uDA
r8IrBWUwp2g6+miSRC3K+uCLjtwhy2Z/xzPNlFlFkDb4Ph5TGnoHe6DhRR/LHLZD
B3W+fnW0qP2ZdZUcjCf7w2W1X/kW94acXgw37NyGmewwyzsYEA1uZqsEYXSHqRGA
nI/Q5a0G2AuJHM5vcXVDZveXupUYdMEWNWZUQG6/qp4yHLLlm2G//qGRMizTp+/v
bdhlcfF/wSZlc2m5GippPETTyZSP2bM3nQNcD3rkYTbCv+Gad84gXu+yZJBcS3Ro
Bx8SeXwS1nruNEwoqbAjiD+S9MAA3m7sURUk4ZZJqnTTXeTihMA/EQlL28kBrwkB
nMNzC2OAzh/Es96SYf/0IrcO5A0CRBeFUf9ONnta/Cyr9E3g/4NfH21f0SxpJ6In
BhLVxKPfCbG+wR60P2kF2/y06fdFIs/jJIM3MftqyeLxXiDGMOqrVi/TMvgLQuDw
NVXlTtzcpihEEDGjjDARZyjgz8Z6as9H5ozQljd/M00yrAIO1AEmAzU5KOHJa9OB
u+cDnxhOFKRrpus3+NGhnSawQoeS3wvhJG7kRcLHyqI20oo/smhQZWJ2zUbi9Vsz
BpfCYy7C/QfG1zeKUGwa35LK1Ih5EF/jSfZ7EhrB+PkXcEBfcDySMp35gYrJfzXX
JYFjlPGBLPSQW4yn8GKh6EJpaIpCkhLyzr1D74nT2tE/AGrOB8VoJLF/yH76pbIF
W2XhhKTfGBmjxQSXOK98ZFKDn58AMb44wkkrGkzDdZaPtBGkGubVn/exS18ge7BQ
3coOC27MLHRVnkBcHj/vJK7opNEnuIy/xuYF8P4iivW/CKOC2DIPf0Xoff8c9wne
IXnuwCw9H8GabcgPrZQ2f8bsOFcK3yj4HnxOPePFUpuNliO+ZkyqGNzttDhBnDkQ
VmiwAm23JUK33eD19cHS1xlMpN22YHsnWKtk18qarN5VeDY3pUCo+uRzw9VJMKpU
FgCuJ+BamozTDIMzgVQkttbS7kj8MVsOHcErHiOCv45Gw33rxafjLPL+e2XGiizg
IQPFjlo/PntzVWw7w9BVY6QyG+IGtNxzRowcH2cUGUQUYiHCW1AfkPkwueyIrOSo
07Lsxa6128sdtNjk0y5FmYVTqZshYOPBnBYCgoLc94qQmZoUsmOsFwzNeZ/FD0Xu
tBrVvqKPefnkrmudVYA7CTpzXKyTFx7kuzP3DXBGUuAj2a9WZI8k9qt6rvSNu0DC
epqaTfacokshCuPF6GMmuVPV3yKEVR6/a86Wo29DC6Dm/1ENTxhhTs6RhcKSzOOH
uf+7jKBCnuNFZVbAV8p7QRmoF6hvSuGvMWaysO3xlUuOvkyvWD8aA1XFCUD8Uir5
xlswBzHIadXaEKS9GZe1jB2r41TS59bExM6bNp7rR+eLaJhPkB1dyc+n0EnYdWan
qaAe+dr9qo/o8297w+zeYmq2IIH23+Bzy2GpY8slIvM8uYM9PrYWUUxZNcJ/9xAo
BOGa6Ux4pnJwbKVv40/Fc3J4ouiX0DAHi7ayFsF6zmKf4DhyufR7YcO1RitGeyfx
xqwpJLDzpcs/zNdU3t8fM8+mDLWMrm+pttzaTj3d4pcP5QqJIHFE2InT3I2ChjrB
MxpdejjQty92ilJvkF6+dBoohw6eaSj9s2z0v6exlgBCDJGAtjSHN2eL8btk+Hkf
eBazPwuddK79lQZ9XuCR/xY3b4f939+yvxqPGaRnJuY6nJHny0FFwSgi9AV9Goo7
YbFO/PpQ1vSVoLJGBm1qWcJSeFKUJeYytuN4aa1Vkz6G7Dla6hJxS3TN+X3ctZrc
zTUov5KkvGZXl9E13CR723z/VQRQyzUkvXXJhVv9yYVynMEtHAnFEb7ukNht0umv
Gftg0SKsmwNQmoped3Xn9EkRUyjAWfijEPwiV7x2MjY1ZIbUj8GE8fiDLt9OJQoZ
zUc1wjGq+UTBhyVpA9bsfNBmmSYUrxG97LHG99Ncz5U88HNUO70qpgtEhAAuChVL
wINeYUjOykaPzv9FCmshtNWUxX30md+1ZcWC2YnmJF5ghnyR4vP1IURvsMCSSVFx
9RaFPnOKnNhNddMAlOWuq+1WBI7pJ3MPCP9wgNE88T3gtitK3y6YYs8VgtM9dBWX
Fp1kI6RwdE7ooMDGRepH56+L894YEIZ2AmxDsIB9bqEucNAjMy1yPUrpPGZdx5R5
4U1rpqsrqf1ZnA8PJ88IyNeeF464t3wEOIuwdORAqiLlmM8WPjGBLot0Wz1pyM6q
7TzpdHyNL7wmHCzUtydt5Ttqn3BeLH/+dBBh/9IfT7CFfZp0DnULRCsyNqo3CdTH
eR4EK01PE1Ki04NBzx81F3MOeJkGCQW5miTFfSs/I931kVg26ff/11D6E6wTegLq
5FElRBLSOXJSjsBa728AWB/lnrgXCYRZ+5ZC7tjeMcb+XJx2ANxCj8J2HD4EuHLU
3r6elg97FNUO8TkSNOqYumYxlwrJ5i5PU/YS9MeJZhq1bjUbsi3wvpocFr165SwU
r4cFwWTzvPIDWT7Mk5ZtjogSNcE/XmXsFoXODcSV9Pz+jPEwArxXPSBooXNzpA8w
4spjCaXeX2AO7NKLs6JOWSdgalBh0ujdbMkIPQBIjVhC++MzyvZFm+39P9n3sQb9
Pntf0F03dzEHILu3lROJ9cg1EgoQx+2WMToljhc9cHImbECzM0L6KS6cOw3z9KSE
wnae9fEpLagjKRWciLysrwpp8lI3hMNsx3hkKyDLIjowjMxMIFDFJFnn9LqJjedH
i/pPecT+12oVGZtGPVwkHsxGIKi3gb9cerOkr6J3YP+VtUnSq/jrl/KBRFx+EvU4
rRtM3MAd6dmaGU0gV7aOm81BzvJcgc6E+XTNxSVKrFWzXRM6acawUk5Uo7klWpTS
4qvofZ4Srqnsn6FCwr2AkDE8izOWiUCOhS/XEACjc1ByIp27uGtkEkseuUoIvZpZ
SUosc3u3AzzrYR9dt6ja+seg4fmZ07ocFpdSvLYcOO9JumMC61F12+gaMkXwWJR0
RV0ZYfRAJiMz9dPBuumOdGD6qTP92/jOeA0wambCqAgyHkBkvqR2yEVf3WlANuVg
jLsGbwG/tRbh1u+Qhh89plML2+pGtX43NNGv2Qp23NWkHGk4Mx2+EFNM8mMswHpa
7QhYlT5kt73YCJwO0kOORaSz4MPIyTdKU0V6nFUDBEUqi86DaHUqisrg/EC+nxuP
v/6GNg0urOSQW6SVchMnsoNYecVo66iTNl/Q3VMqF0LEMSjaZNCIWjVtaAiRsXch
DoGtvdfgenUmeLqOc/njphrL/nyNV0DwEq9KmE+XskAjmg0YCHEebYPUvSd9xmlp
tnqB7qi6P+M9wLA+9xu96gIFdLzEtPdeEDy5vjbFVmEVd08FWBVI56z6EtC0bNQk
RfOjrWTeTZp156XlwU4ICuvSEuJf0sIqvXitYkOn0TO1MGsgJY6QjHQd6dkdbXDP
pL0gzV1tWBHDe8sXWir9rtQ6VZRMrrfpSnPu1bPM09LIwfozHKxtQbgXc4X4dIcT
69uqln6cz3cS3pMp04LTHcZMg5Q/vYqgyIJUylas36obhbUGWLTjp37F/s5liJXf
HMzbXvE6R7k3GOQIPamdOu6idFqVf+RkBD/IqwHP/8JgN5pijdJdM4iGArDMB+db
fjjhjUnMSqf/zuHp0swGxnR4W/rCUYY1QCu5TqJKCNvQTrz6QdlJ3f40k1i21oxq
HjVJTi+za+nI9aF3i8uBW6+Bzao15qi47cqHLBHKUvYVx3dAkqzuDA73jo8H1CDf
poFqeSZ9jZaosS+/KFBbYE75QOraIqCG17R92VotazLXX1j/e6Rp/vefckgdhqVz
M9f2jb5ggCUS5ZSDFHJTKANJ+tlL54VzBQRITLB2R/EMS8tXZBBtP+D/nNZRdnX9
7YGbV24H/Pz38N+6HxCJF9XOjOFhtBDJK3y27qKJFqE0V/lSGB0pXc1/dNYfS3RV
6qVd5IEyZkjfDqGNljcuG+IhNYzLIdC40TwzZSM+RS2yVaUExZCjqHHO86m0jqhG
3X6l7nAPCwuYLqs1EFG593iBdRTwXQGpzT+j86mK+u/5ZfZgas3MRFdrU4Ybjoj4
K9U+fmkLP+NkTkfoT9ryDe7KIexGKnTDFVrie/l7DhczXr6JDXXvnXbrOVspDxMq
DSl8LOLaI2h3PAOU+yxv1mEq9d0OYSXzHG5/cMR3eK0fzeMRBzFCY/uvVoeZ1TSl
vhaFXhc94dIcRVK58XP+REn1Fbb7qRVcqgDLoX7+By4Og83QNyO6y2paK/wYdKEy
bSl+l+qAUo6WaEY5SuwHfqupd9OIOEz3WU6kKmxWJu3nK5IFhoB/sZfZiQCvXtEN
i8+aSSqnlSJKLhe2E1CgErdswWYAI4ZGlp6ei7MGQehVexGfXsDGtg7r+J4vrHOJ
iRerUpq6/rGcakHzHVKh9SClazkD5F/sX3Qd2OgLofhFe6+wCThwboP8Tj+YaIO0
hm1FS0OBR4PPHlfv0d33g2joXK4OqDGUY2J9r95zFleewCNg32x+FR6kZ66cJ5UQ
hEUXfuIQE5ED0lrrJJ63U+9Ff/PAe5CV8JeHD6gZQ0bCtA3ZhIaGPFR4l+p2Fnj/
O7wKpumlaMk7cSRcVd81kkSFRRbcMZmf/uU2nKQYct+dRph82s5aJjVmr29IaKp+
9Aa8wSK0WIMWjVlHaWcPOJ5mMkWrs6YY4n5xGDQzjHDc3qMxMsYHw33GzsGZWwtK
c9eLmB+IJRcWB9Ggzgwpz5sSjG5jd6SrsEh0qkmJ0unzCFqDx/s8vXYlIDeCTfNw
zQkoVpoTgOgQOKPUXQGeXmLjMhNsTw7+TCmd619r/KAD317fKiMA739aLnibPfgi
fZmVQF8hiMcY8CBLBdchoSLJX4rvuH8gRaE6Nqfp93J1jnnuGgcXeaB6KBbxU3Z6
MYgsmNrcMoK0vgbUAMBt8WVGEvusGXS25jql64fkbf4UNgggPMCljphj33zzfVMu
H+P7v6SXd5hftYGK5deBy47VXxkgkeSDLsvA0WWpcBXQAvZOfRsiN0Nv1VYtbSKk
LvJDXh9gQhGAP1FgnCN56b8XrqhDtqkR55zenID8sAMK96kDDGqm8gVrENDMXZZO
P4i6fQKUSkhTa/AXKcEDHym402mTTVhWsda+0lqmxkM8jp21hVtvi8+ywH6QFivQ
Zwc3OIqL4zVANP7qS2XqvbpK1ZnDrFc/GAbjZRP1RYocAkBdw1sMWqD4zsUawqGg
en+rF+EQo9nlDRpfmF9wd4Ukv7jZbTJtwDm4s66wnAlXlOhtCLNEz8UtDof/9zw8
1ak8yZqVpKiXtCol+sR9/ItNaa1eEoVRqQ5GV7wvI+yCokA/E0otAasrR+3o+wxr
Ph+ycqGrDCa6JiOrv+nQodNRgdP180lhXkzoBD3/0WbAjLkQUhfn3GmhEdvr0sn5
ke3MHeBa7wC4velofrqW0ZrWiiMYknYE29HjxLgq3j6IsM3xcYEfZBeCogl3qC1Q
cCZhjzr3oxPMHzpxG1WSdkp3auRGqYEyrOB87o8m+GC4IN059gSGJhZjLAg3IJDq
Jnn3YIKiq4TZ2iRlI6HEya08xhqEmeBv8qDjvNU4kezMBZ28RKG1b0ukKjHW7JHJ
iK1SMKBJFk8HP0qtaeW1PPoZ8HPaHgh1Pae6W/T/UfNK4jLE9JDn6q4A3HXSMGBq
4SMp6lhW+92XK8rsbQdaxdd5fRERBj9g+AEQh37y/rXfYf82BZErUxe70/XIjKX+
CFDNarPvgPOkNEBbd0+PobjqbqsBNshH0EiM8bKAKwLnGHdAAF0Es2HBLBzQXjSY
ItzaQioD7deM9DMPdgNNk3a0WRYbu9tn+S8cPWc6u6krH0RdLxekyvGEO8oSKVfA
dpFD/Q9jG3xUbuL6cHAdUakqxi408E0qpWbOaz6pwS0jI4h2TNsgD7hB63hNasiQ
2e+naZ6Dm1U8Ij+FVC3/+j3+Dk/y+7BmfkafCF6ux1529tyjV5k1Kh1tsz6QTJbf
8wKGGnCAHXyase3OO2D/sN+ykREKPyXhtpU9GYY5HgVa1eoIpXNY1LCPy0TCE0a4
g6+yNkFXTbsh46V4vin21k23T9f2SUGpQGeMbBZUx5WGEuykO/fu98wGuqZ88rs2
Lr8KjKfqrrgiuQnaS28uoAqDX/nRqLkMIZXmbkw7H4jKoJcBfybRmToF1mbspO15
QDd45CvAckHbf9/CifEVVfOZZ19IiJPLkF25cojCevqcSSBl7mmJmc5NuYAGFM8E
RPBp3xN+3btAvCrfLzG0ehxD8y3ru3itKqb0HjUgiVhr6K+0OXMuJ5nS95q63MsD
LeQaybb8jC7oNhvsGiVinqvR1Ai3HUMIEEmtezhUQifpGU1TE2pI3ADyMlROTFGN
27EQog1jO0GtP66xQMQIpfPd0ac5hr3g7Klko52hA3MJ4UtBOYiuL9VEx7tKIuhb
6VH90hg2YHw4L4OqHcKIVnELgfW5/jo74Z/k7wFKz2GIurHUlJAduqCXIQ9gbJGx
ryoJQt1OsiJ9ba/2j1LepKcTWXk3Oc4FdzY0rYv4CReQVfCni57wfJRDGNPzIaYA
8FeYJwrR+BqGXJWXX3xW2wKOmG6fXE86QXgWDCmoCnl7iLKfM/WeuyaAoWpeCm8a
ZlqPWmOefJ5Uo0MLf2gR7GWm3WK7xwZjyB0QlWkekcYCmPzDtxNWpcRMnM8KKVAg
f3jI/uetaMrj020XhaQp1b333Jy04qu+SDxSekvmM/rsppWCEapV+AFL7Ql/8dJo
+S8JWKQTLrVNOs+imqjpiOpvhXmSMlU2yD1X5ZTngSos7HhMzrkRfY2K3F7ET44d
lrCkoK/Py1MqiJXtHXH4Vuiuc3HokcOuKfEgPQ7rQMoWs/aY3EUmm4zIiKn7b7Hg
Gk9erdzmYuP+rsdAPGpfUX4XJR4DPLS9pKDWDXf6bz4g/Nhazfz9L5v2MIRcH7Sq
7+6Hgvy1dQmuYegXa5k+vtMRj1ALeUkSKPK5f86rfj2of7fGtYVpTiHK10txe/OW
kAGfku8WjPhV0d9A4zF62d0CMdigPrCcsBNKbc58n6ewVOAi38tMo3o5w5n/9vQD
B8OrLhc2s7e0rCYc8e/wi2ucX95VW4m9pI+9hWhop4fr/ZVl7DmxJ88QVmOc0CUF
/uCpxM8Scy44vEXQY++oTv/chhjaxyKykIrb9alLSV9ln4Lq6mOeBC9S8So/kRmo
OG1BJAcLfm3nvyDf4/tZ1AebF3ZPtqP0P0PQX/7d3oaqZvR0ifj//HFMJahYqbrF
lc/XyfQjnKmsaBvjT6BnE8h3mLsS0s4/DxCQkK6DLaLTeIKj8eOv65VSE0muqaRp
0ASuZM5hXB4OiOU0ZA8GaZlh2bQUgx8yoJ1P7/+nvWV7PZb8diuOPPl5dJLsyU1R
EfytBM3s5EBUSgoO3Dj/dqydrGJ9lDgAS/NIh+OdWPHTLKnsZhD305S/dSkD2Wai
RZDcrbbCVIL3TeIgDeKgTV4laDdju8FlapHbN9cdPFRvKqv/NpTQkIdPCgljQRVQ
VRA3LFR8YXA5wOIPTaiQgY+tUzNv5PShre65G4FyBSY1t4DlFxd7BYI96T6UlZ4k
vZjoXlazy/iOIGR/1ZQ8dGyFYaNP1TklntksdXkrzRc2nN6kq+sjAt2dI5rcfrSt
2fpsXQE2UabmKb6Yp/pWePYrXJ3uPkGBS50GzdRQhVpDKOLqOP9Y7cXGLgi1WqSz
7ZZcQxba3uldKMIq8NJXdkDPfSNW15TvI0H7uYEB/sE6pwd/MaybZY/c2hp/KJjv
9a8eWX6JgFIjOvU9lSzc1Tc2QbUCYLgXt0Do8FmxpNq0lk/3YzknoG1Z4OH708Y9
5f+ALEbDh7K+eBz8E/DgQxYG4c1IFhM8Hh71Uf/Q8yz6TwWEsWJcZJBTXi4yxQ+h
gGEfZfQ7har+ynOu0YqXYKiOx8aTQANSHLVObAcpnYuyPLUhOzbZEp/UfaE/etmr
S1bklD6O597apkodTVxDPCdppnEsWzj+qaOdG6ZsqBY3eB1YXvLRG/jtnsckN4+5
LRiTb/OJM0T3K3NJ+v2r34G7MeJZMGqboaaxop9eOy/1GKYW9gFbVg5nuIaE5KlZ
+UAXAEjaobc0sCo1cS3/65NIv65Fw3ODSxOn6LvUHrVlMj8SwnVSRMgNvfpNKqu0
Tvjgk7qdV2EyYUtM8opCKfdatGpNQKq/EN+KimT1eDn8GNP7p7TAjPsv5jQlPyIL
4mgLYjLvQUw47Q9fuKGEacYasHuaDAPpCW7QV9RxyIaqt9PhZ73ey1tPMfspVlE8
YXPe9xlljuLyAS27XWR8yWh797OGcI/lwEXPRMJtDEZN4vNu2n4BSTPFd4oQ/7XR
hI4AkSPny9+Vl1JR+4o9+CtZDGnIKwhu7F0SRi8TcAN+frnot7H5t8aqLnP/Yln0
cFUKZeXLHPJoxitdDvVr4Mm+HogrRpF4tH+0zccCJ+RzO+3r3S6hih37PXeTtuYL
zaX+MLg9QrNvOrj2hPt+8BNGUYXUnm2p36hIhPlDxqIUz1BI6zqzhB6rgwqWNhIs
JAY6lwAKqzMOA84h8FpS8mfgsnpjCDtxq0PYJ4C+qNtOqPFT5fIQVFLyX86EbKs9
EWucaUBpbJfldDGwiel8HeQs0liXrUmiIGgHL9r1BAC6zCJDldjK0zJRMfE4Neld
kwbbGd2i3i9lZke5PQ2BcQaZzjWqpfQXkD3/3iiaW1aZ1gZuRnqNAxKQX2rF+RTP
fKQlsDq0g7KWWxDFM0Lun8fEYgX8PFEA4hv305fqQiYVQ9E/ptENQPLtMH98eqip
22fkGsh9SpGIotXTJynIIYZFYRuPhQkjKmZosSOEljt3/Y3NGqqJ6Y+gQL3LfmMw
xlvP89P1BTs53W1zgURPGskY7WJ0mLeEbfy1Y7gq5LFaoibOLbrVsl/IBFMxsipv
MZdkNVvJm/SN/EH4a3QqPbRV3cFOhdKC9EX5xDBtVb4Ql85CZzeHHLxBYHLpRphB
uOR8mP4CuPH7dHf7OGfr4pOHObINOgRTITUaMAy9ZESbS6S/4BFXBkdv7qd3jCe6
PNNZ2HdDbVTRwilRE7xzblTi6Wbk7wpNyka/TlZG8RM+EIe/KsQiykgz+X2jIn5s
YRuHaQQr9JWy8XTRo1GZCatdcg/9ae9N1X1CMCwzB3mN4758ywxcozIzM+B7LGKq
81MUZixCmkz2/NldC3jIqvMeD9IqaHvwWfbP1bzYzW64fSJayQ62IPLUpYu3Y7hq
doLqFCotOCIaX/H+A5HNpW1HesAh1TH05bMWNEgr/nS0ew1gxxhwjW9lbIg25Nse
aC11ffuhYHMzQrI11zuWhLwm4Hn0JlDcse5ZrFKqILzEEIvjZc/YcvDLTIUU9xmx
KWlmHHomg4Ew0CLfVXzGTUBteL5EBH5e0rC5WhcKAwlgEahsf5lT5zTobwgOe5PW
rheW/3O82MiMkNc0njqTCPOHEFgdYbHOL25/UMsYJcAcwSmgM65sZkP+/uoESPls
9w9K1DpDbByqmru7b1gjtBMxvNN8znk7Y0Iq6aE66tSLzfLqZourpvOi2UCyXFWP
jNYy0vOv/8l9xyvl3XOIFZmDPD9seqbVe0yBrdKXRRrbvVSxJ37w8uOmkwngRsfE
NM2XwDhALe+0vQNITpzV1d2NF7js3fMp+N9mcXwpxVloSZpvhgGPv4R0fevXSdol
aR1K8E2qDN9P1Onq2+7FE8XboHLad0PB5vQ5CA/7yKnWA9Swg4a9LTBEiHHDJJ30
ByQeyGVj52auYxxjHzJ3OVpZm0qC8S9QH33sBRTpAjwYYZmWqm8MQwaH0nD0+ksq
No/FxARW1aIEA0ArXKsvg3Puab2M1v6rwbz4U8lQuGiriX7y40bqXpAfg5uYX19w
pCYTTjKc+x9D+khQOm8bTMx5jUB2Q6/ehYa4+MUEJHv9Uf3S4rnwH9OSqFv+oByT
oMsXNNGfN+S8Qe4Wtpu8f8DgOxg9nlj0s6NqaEcKElvE5cXt07RZADh/X+dIl+RX
i4mp0jJX1bzjnGmXLI7WXkza1AZu02ofkUBJrASvIsUNE8mExFwFlnrXMSCI1Q8E
R07VT18PmktB9VE4D9S/dKM1oh9O5EVWmaE4ZVS3NXWsgCbgZdVzHX2qjKbrpjcm
4YZBHk3Oo0/y5U7lzUN1zEw5NLaI/hIQtit4P29FlHuMh7HldhTWki+G0bKdx6mw
Zb0F4YtofPtk+hLptbSQCp2XuQeFNR3002fy5AKkYOPPwGsfKBCTTdW46kda+KgZ
Xz9KJqp/0xU8DfEAldqz4VoZ5ZLZLpduQ/jkwkyuRcF+/CUsH3+4VGtJuUdVKpbP
ueTWcE1QAnfRZ2MBiRCi4pXCC3OD/vgeet6ctPp/6GlVRIBL4djF7K4M+cA1SDFz
sBElq9SPpYBe2MIYEw1vt+zZIr9AJAUTGDx3QIBgJV3KhBG0zGe5D9AIfZHhcEon
Yds7+1pUeKH2zBSSb0OiegANxMUzffyqWncf4lQOYNU1/mnEvyE9ksgmpDhnE49v
snV67Sg8BhUxC0x4Gk8ZZYFtizKTVTXziNgYsMTYHKeDu+PVPD6USm3MqBtpLCOg
aFPluygP5GTdcgnXjHhCOTzCabY4Bs33x3YGv8V+FcOdkwQkr2LnkeGctoNqFH4N
Iu3vlnqkrjkX/71i7qtdm2ouwwOQyNMgD00hT4WeH6eEMnJyY6Yw5SaBA14wY7yy
5Bla+iJ9/L+R+3UW0qdGaAUi+2lgXSciuvDw6/hgKknvrVgf8o7JjFFHMlgF5eBE
yAc30+L1Rsn3XVxZ72W6XyNOmKB67WTq8+QX27U+VPW27H6Lfel5jfhLOsKnmqn4
hPIFVyU20AzpausGh+pXPLFCHIpSuoRShRCjuNSpO3qcCGorewbny/ceE81YWza3
b213gccefiJH9DnoFq0xTlsMiDjF7+tl8tzVEDuiIwBz2B9qdhAL/mjS8UqF6fbw
3PBpVdjOeC3xYTbdKC06GsESIGcwKgD4mxCc8FpPY9EUhQKClo2Sp1Ogq+YcIspz
pn4XNdBO6wiPjlG5DibzJ+qBuWWPZt/1Oc51/ALXJYEMI0yEuiOEvbuUHhcpOPzx
fXa9rCTpmCKZs1fr6P7yAG7VYQTFkASVGzXz8mho+nogqTVpVYS18TED0tnGamdO
OKb2X9wMlBiS1kBtd2cVDJHjyhYjf7I8lo3rRYmApvqeDJPKv8IUo9oHa+S/7kPF
Ct4JfLNajOSFjIGiqCFbT86tGVNqin7oOpVPZMk0FN7LDsPUiedpXKUdHZjvcQvA
O5/jrPyu5LJfWt3bMPW2MFiE1KRnpgasRoWRRbF2uyjBK+hJAZJyy8HTDSUulLoC
ZY1obIByD2TE3YShuKgI/cMobrzYQf9+ql3xoW6Fh9fIGyVcUbrO77yu5fK2jXzX
dnBPTpJEiUPIwnKnBFgBYFvSYX0tYNoU7+fiyrFsDOosV9bsY+gBCBFXxqE6OCH9
RJ8TDfjGf9hYC46Ce/hwBLrKvwEvPtO9GzO2HOzYY1rG8uX6eEHu/f8f0VK/TTAn
t/bXAW813HwuLkU/hDK4JPsHMC5A6r3aR2Iohj0eRt/e2Ucujc8KM4/dwfzyym+q
PsoZNezlgGZ/eIosL8OopqwdQKvG2xGafMsMxGAC7rmaGZLci3QGQKjO1MNFeWFv
J1ALMJEGqUVlKIq0rEuFsiEYfIXha+9y4zLIaBQwPNEv4bAGxfHDtLDJM2dknEgl
FkxVij9v28nlCVapX5/Q7m03i18Rz2mqGmYEPrcUEKTr33BR/ANNd6vj8Zc+mCON
T27FVnHuQtSgT7oz4bHIwZIVXRmBBnqg/Gy+G5prNYLwgFR7rV7kWodTlesAqN3O
O2gqnvxR6L2VFHoVSY/FZsBm51vmmIrLtiJN1lB82GPaFo+mdY2JWvBs84k4+j4m
ujo5CRLNi6kbqSvE0ptNhrblOKcpiaB6kJvlybTVn28PK7JXow4QvYq5YK0Up/zo
fHYnimzuLj3jplU8F0orMTQwUnZa+t0VL+kr6N3Hgx0KGU81pNGk922K9M+irsR3
3d5tTyS7rxa8xlj1OMIR1MtwXOf5Cro+GyxtIRj06lgOXaHwOsAwha4UMSeo944Y
tAMDRvqFkO80ezMymFZXNrVI9GgwAMTWkhXBrwFAFyLeGVf7QVz9P6CTd//TDYVa
cMhbNeC+EgYj+z01mKm+MFldmckuP03xlScUUk5ubVjS/U4pWwkUftfAmEFqeoFF
TKYlH+ORzYdWoItxVnjcEhyg21YE5sKh8U6y6UTuuwPCXINBCoYVfyer77CnFs1h
2o8zOMSCgUphiT+4RfINtih/ugvJBZmS/AYsSrNsdnqL6qNfphQcOAQO1qN0arzq
/tNoSwgMGdIUMmwn5kGbsSDBKU5hAKISTrn+s9O238TlOekBWaiiSF0hgG9Vzgjp
GOLs4Xt0WAnBbMVWGlYaDwsfxeCzhquW94626jILt56QejZqvN9K6K7pV+vOAfSD
qEzrwY/+QAaneRuzE867KP5EM18lyfzo4mDt03NJrShtT73/izkq1TmrNXsB+jS4
2HGH7dg3PLcDE/8FL2yDmupZ0ycHdcbWD+prRBdpAY5bpYXvJCnLEa6aoHQSas1s
+kfmxHACVPByG1/F8D5FEwadPf8C07rHInnAbPskcX6iewYXp6XbW03jwiSmlpDP
s1WIEPtFvyMvtYdzKJ8KVKs+erDbj6Qdwl6WMmrfyzJ6gzPRGkcvqeJrw7hn0hzn
Nqe2gZ00f1hOYNwE3en7QZCnBYkuVl8EW9lcSrOJs+kme5JztTdPyeScg8B3y3iR
freYQ709QvN7QEhvjx0EqcSa1GlvGodyd8oe/+WiiXjNEwjc/+8dbo0z+DoBIUgW
yJHjw49WtSFIe94RGnGZojftN+VZH0XNCeMRrafnb7/yvdWc6rtb2uuEX2Y2FpDk
lc75dkKIKd10iIGWMIu2zTFGkislkTztZBIe1pE1BpK0Gzy8VLo6MPJgo2VBDUuG
+E6OzKsCg9To8CtK4yMhZ0uWT6IBLA0nNhhcZIbwVsoQUHzyACAH9tEzSB46RX6t
dLv59YGo/WH0EqxKCjB6OjnZifOX/f9b/wq4SM3AYumvuZhZgw0EA2tykwHW0srO
JLETlz75/cVfU1U6zZ3y9iD7U2CbKNGl0uMVAa+wlCDLZvYaIPczvEfe94PvCbim
0rYM9cQun20r2hs0NPi/jlCaEyX6jrMos+VFsz2lgik4T/BR45w+7XXft5Z2sQ9c
iUoIJaNOl35+tTYBFjk5wdX7FcSe0qcVG1tCee7kADicZhocAuyEe6CmqdkcknDL
ZkL6j0+UpY+LHDiQw+L7SZH+Wa0U2MtbYYroomep3pdJU7uKx9OiYY3fdVzetMHS
kDqRSw789IUj+R67Y/2881B8Mt7neyzmdCr3o2PBDm7113CreTwZdaMSBYzH1wUl
9jmjycmpUiW8o5Bv0WFR0LILHrKTnisunPzKby/DChy36eHtHOseDNojjm5wtCVh
yka4oGpKLG4dA43EZOep6HWHgh1v3uZx4Ju4YzIYWrL9YTd+FX67gj9CB70kBkk7
VF7Qw08dgPr8eVDu1Fl16y7Pc6cf47bjv956MjK1p2gO12uPdW5zLI4WnFJm1/nC
WjHYuAjhFCSPzV9ccmnpHPf5JYV1cWJJpA8N8yHUWZWHsu15WMHdUjznkA3QUT8Y
NtlRFsX+g17Z5bpAJ3u73z1sdaeosDKh27J5XPJ9vqwFLtSszDCKvjV0RyJTjR0H
ce4EO/y9TDPrGcPwXkAjoOSaseJlhinfRQFo2FBdpRwXCRj3aU3TLEoXkC+YFGXm
dhhuxTVxrr5UVoOE20lpQViA5r1Jb//q6mCAePoEi6Qz3ZBc5HPMbqj6pvBHIYpJ
IDGnsmhv0WIQTqVkD15I6w7MzKpsIIMptWXa9Nn3I6JEeL2Gg/HTC8wwvnyHHxw2
aStRLkJKSqgJuekUsYhG9WME+0qkCNonQo5RRe77eNpj4uC02NWDWriqthlDeS6Y
MYPUiOzD1SB70OFHt3m0A3/0h2juuJDzuh9jTFjIG4yjFXfn51giZBeP82zFZnxG
q3rtyctXmukRg5hrB+5UBjqbgvqKcuRzA8iXWK9dZDBIhnmAVYOKYKoEgGWExyPw
ws5Cffdxnp4yZPZ1oArVOm3QfLUDg/DqgyZrhtlS2L/wnj8sa8h0X6/2xczkjW1g
Toz73IXhJ3vrFYxvSAyn/ZE3f74meycFfk+YP9BEyyZNMlpfLQHFKPVNSXfns683
aPTnBu6HEdXbnryZ1qCTAUrQ6IswDAIRst5r5luV+fiKxOlpAhlG1ANRx9wBOYCd
7dA+NvdlLOjOUIi2fIBqRXxRJ32Xr3JVhWrvQD4AiEA6/jKBqQVcEAL68FASUVJ9
QkdheQp4ti6ojV6AIlpbFEvz87RgvLWxKL1d5DtUfGd7L+pUxhAwTp5Jbq73dMq0
RUfNwXrhwFDhklcpXxdj44D/ydYlCf9pe0wpXVgWeNeuLnYc8ivZXfz6CziSiqtW
DtrBPTgOh2gAfdn5ryHKFkALzEgwj+/Gx/rHR2A/u1t2tvvm/H+4jEwpCD/tfgyX
UTJSTc9lRL5DdM3gZ4jNN203E1ygk91ZGPneUHdg6zi1UgpEoteBWUBfkVqnm9Av
q3Vp8FGryUoyWLQ5WgjeZ7q9MFp8fiLK3OTmCPKsj/xyo1Cbg9eUhApLovGDolK/
Or8JFD3WHtSoMVUM+YtT4fRYPwwLKRxQ7J64CDF2AgdvcRJN3hbGsYqCv6v+eRzr
yD8i2I1g99csvgQvISjD7IC1f7wGi3xzOqgSrZpfVbgmZ7480A3cdGsS3ilKkWlo
M3lQyGXns5BjyegFmCa5IPN5khxxkXulNYOvTW07WM3SJMtukI9LOELIgbqKecDS
kFl4QtP1NrjRdw6KPTP5+sICE+DdkKQ5zMdxSJTQrCwZKEgKAoWAONCVYXjD6bVM
kr031yrYAD6+S2tMzOE8yhCwE87iKIr4cSwmvy9vRaM+LaxVgmzMQnSmbjExXHEP
lWtLH9MoDfL/lg+kOAWA0j1Z77pkS88oK14ebYL0fy+UPgyX/IXvmc5r9QLa7wql
cQUiMja/UatTr5NItXEsT2n6YcP8ZGyOjNup89ogyOYWLxaQsmJSGD0ClnCij9Rc
n/VOLnicVfltKIUgfFf+90sx3YE1A0U7DGJlxwSO05m0RuRmCmOTzL1wirIDd8hj
8mt3hRDqAs/8+24DBqY6niXIDp5i4d9rsl1mRp8+m4Vg2HhN20s97tuXlmL8u6bm
5TWEmRF/80mn0l2qO7tCLgDVGGxDpL8EEKB4DHuB6YZyywZ+zXJxbmD3OM+wTuK8
K6wWr+bA/aHJ//E6M0L5EUIjCkHWHdXGQ2wjJfFl8j4D/s6Ky6xzojqPwcaHr56v
1T1y9qyjMoYQ8isYOFS8iCGdQAidmQNDyfLrmZNupATTclFP0H4kW5TzFb5EqKlJ
OyPqBJ3NhilQKFQRkUn/abKzX7ulnQ84KNbVCrWMzijh3MHotUQrXxz3Sni/hyav
2VajKHoCsaYavU47TNEDeSRD2XD6mi73sZ/2JvRX8Ujq294rKyhSnxSufde4UQlO
rJgVfIq6f0qlIrykAjK+H7yZCtuGsWHYJI8k8p/mae1z6bDKzf67kyS36HBqoFN1
Pg3SZuCQrMDhM7TTxxmv1Qg+CAkf/BzDPHL8vkqg1YaxxoUg50Z9Xox9ud7PUsyY
zQdMAt5ZL8Y42wagWA6vaaW0jv412MG7KT9JUriOx6hw+se824cmfWA1M752xzBi
3cTRSDH67ZD98RjWP4B4P57ZpB6pby995j5w0094R2hL+7KodcUMXa2kBRO5xnuq
T5LvDLdLRw6W3f85LMsZ/3swCSSb4DwxHrr0idhoQJtyAq3lrvXCi7dLOCG+wrSC
Y7fnzDI+hzdhOCCTMwn/1Iel325ESze30lBo0I1OzbKuS2s5dikpbb8B3qaYagfP
BMzwg6Yo5lVW/87Na8k0udLmbS3NJSMtFtEvXSViexTLhvwA3mPtFa/txeQfG/lf
LLLqALRFfyHIDRth5wnyojGzy7cJSGnT1YWiddRt+EYal2s8IV/JeDLLZpLq/UoB
/STrCtO4HM2yku3K5WrKL2calbxsDgChS7p3lt3dyYcWmQmMOTq0hwBZnEqIhPRn
OHGZl6tC+0v88LK6Htke+gCR3SBYDSYsYEig97SXsavSNlyOxpo8Yx8TwfOROUN1
o5NH7LoWC8sCjBY0yWrKt2nQpJWa0ZcMS1Y7qwmc2fzneSrOkNw1VJWnuNktwqL5
br9XvFmc+7AUFOTCrHlKr4igieqLZT1wAOZa090BkgerAgsNZKpYgbIrBWj1DIvn
NzpDoD5NB/IzcBhRDf5Vgun+6V+qRhfqp5AZT/SBa1AuCox+HXwv7G7Wter0kYV0
r7ek8u3keuuoOuzBG6U8rBh2onk+nFKj+B30T1GuYHpHxdW4EhJh6cr6Igb/RFID
om87og8BwTtiTetQ8ZMecGQRE1zppXlUOKe3nx6ihKo3mMk+yS7tYrLYJ7BTtnLA
2w2NJM1qGXHfAisc0QoJYppROQ0qC2EDwi87DWFgI3MhOd2g6/WprY3TpePtC0Ie
/5IN5DBkOWOlcSsUKOC6F2T8vzalsWHshXSM7v8XBfHyAI+j2v84239SJKlypQiV
QkeHtvQ3HKF+zyTW6TWwWoT9zqY4tQm+0GgERL2qmahx9QK2fI0HEOrV3Me9TPi2
x0LWbdTtEoMh50nkA5GI32iE0Q9kD4y2TPmZpZ+x/KJrMQv3xc2ZNQ/MrwRSvzFW
9FTGXu3sDK1e1wo2bytumnuNPSVtRVibvRiypaf5FuBB6CnW+TfGb+bSMtNg6g8e
449ex1HkJ2S5ydG3PO4O95vH0zlUu7zeM3vYf7benmHJr5lXRpdIYkf7e9fhGiQm
A9Xd03VoFYEuxXq86NRghbAi2lc2ZlFNYYtQFnuFsedu+EqEtxa98vDeekDLUUcn
xqU0q5nbVt1T21ieR8gBEjV5j8CrQL03MxXN4ne3l8MkeguV/5WcsWolq9u4J1Kv
wOeYB0sEqtZf+mCUBx/qPYx2q7wYC1E001jhnn83+7hd56evdYL/6bgbXiQzT6tj
7FRiCgjDHgzvI4ujcmzdvSyxAQdZUFWaAvfcm0aZPFCMtZc91vNJUnbBFYQ0epbg
N2lNIGvz+DC8/P25TQ88bXQgnZ4q0tMdz0PRAM0TsMPLXMlsUQucTH3TLg/5ENIT
UEooEredXS+SkS1AnYtZCR58UfwhcfKicX3SEDlNvvItucnn6m5eMJT8sXDCrAbF
X0sbMrPow2g6OmgWqGJuFWUSDCulxIF3eNhqeOqi6aivCi6n14leMC3fTlQZ5Mk8
bM82P+TO6kVsALHBhYJ77OENezcngM4tGq6VVa4si6Z4W6r3kr13sdX9gfupQFeO
rPx+krPvTMSi48T/PPerwewfXqvPUdg65C2/6n47awrMOUjvcP2G8SpaSAUn8aDk
FMtBWMukgC892DMKdnloaPLD6NxcY9ZT5XykjVUKV9iBXZSdPkFDZFvouDdNyds8
WSb5pvIktHiSdPxmfubgsBqZ/X1QEGaIYHeYwoCorOQDXDes3YJndWjBOuItAc/e
4GyH5EenxYJ+afFLMcnTKJh+UPytAz/bNu1REpqFMO6rfKL/rTDDx6o32xn21bQN
qUoGXBT7KBy8FvFvaVjEKP5AfOfSJ6Mq9Rh07LRxLDT2AI5fnEa3jLPJQXjC70uA
kyvTkiUhe5qk8cTRLjX8kv2WwM1WhiFCjeQXOcIYO0K53BvHFhQPo2dUU11w7DNT
EylVgZY+kIOecC6pOMWgRWS9dK8O+52Gs9dhAHmS5449L+Q09lEyeJqAZNos5ULV
EQ/9r71ngeZrf3amlJze/PdIislQej83d46sYQZ/SdCzQut0trEcEjJLH7JIUG2W
FcKvTU2Tz2+0Cw74KRLJFZYFSlZ03MQRPe930cF6Cs/jC4q28ccklrtDAWXi3MA9
qlE1avi2HgRTGjXeCqk7Pu+s6FacZu24Z4iFtCAgb954igq0gttfVVBpDZ0NjmTB
Hjs4pAZtPhFVdC7afd4ehcWoNIKCLC/PrcUjC0ODrIYy/9IdZ5EW6eKaMWHQ/bij
rEt4qAXtuc6Go2PFJT2v3tKvKhaSfXLUwL8fsnNlGzObTCSfirCDCc2YFMiAyO9b
rW96sAxOvWPaCzqSzix9x5oCGBwBViFwWzkz1aKdgmr1eB5wNbO8xDb0bHbKd+eQ
eE8VJJLKU0aeYtnbjPM5kLUoY00xpENQmXvmSLGWKBDtuqAiiQve/965UuqVHVs9
s/nKDGtLFzL3UqgnhOmHTKPtETMbD2XTR0YdPFTQzroUg8sKGnX5nxH3xxDgVXIz
Gx4iBASESyTyJLZssMQKIfFRbe2F+7BfSxp3CC7ZRk4cgK58Mb+qy+utelXGE6Vi
FDl1mIxwV+IumIRAfH7QedlIqMPnGV8toX8YuQhEMUh/RE3oFOgV1zGdnPZsGyX4
76mBDcOkIrS93QiGTcjkv0XnQukDBBhkfGeCOx5GTrwe+3h14QhZ2gESmjRdiLGC
ePo7T81FhN64uajReMZjbA46pAqGnukTIGCCLaMbfZ+Mfw1ZMm/DCAWdQc5edsQp
K/2D0x/pkyH9FQ4SotvrsFizLFA7R7IHxKtBRTO5YgajHeumpDUbv1IBkZQa4g4h
r8cTsRHFYSQQwZ/Lsq/dsuHoLKK3VsSP9jQwx7N7Tso6undvBbbGTC696ezxwWlM
C/R02wfIjpzAAETKtV+9hKhNdN+Xj/iigaMEkAs3sUr8POkTSD/gQ1zBUoKbeEyS
+9US8IrMdIcqOA7N5OgW4QTSWMyrp/lCT6h1oPRtNvOMYGsAdX/QqGVoVQeNuaHS
+kSRV8YCXtzsNSorrNMrVcb+zzHJaA8IyERnudvcb9N8kJo9J0ZOQ0NL4Y4t5Evq
9JbHCO+nYgDlFC6T5/eE7e02eN9wAou7zLpwiGvULRMwVR9C5dyO8hTNIci6hat9
dh3cP/u1or8SXanU003Z+lAV0EecK81vApPXOHm4lXz7DbsJRNTWwFTkmNYQ3HN+
RLWNkiUQn084FxRsGxmbgfYRimk24ckwYAGpLMsOYeSsVyOBi4nrsjxOnilDzNle
o1+4XWRL3wzfQYs+o2suamBXcwNDeLAiFuf6FpggEHthhfQVhI6xMH8I9cbQTu1v
eaNMIxuJFA0HOt+xMHTxPyaOwuEMJqD32SvUU+fIDdAr0CN+Iuhf/mYpzVWApV97
G7J+i15DJNgXiAX+9eY5+llW4ChWWYl0xyqUOcQBh5n1hSPa5o4TGuhwPibtoUxR
ONr6c2FTevALyPm/q3Kl8rL4Mp5Yob4Suwu3ZcnF9dK9X/zfMHjpabQFyouBxT+p
dxIE2xOkWLr8NVNOmMx3bT0Ctp95iUeBqbP3EXeI9BmSIENbBXsd144/HOGV2y+g
s0o/OntWM3ZKrD2qSJYEDNf/ug9RXCd+JRYtwy5kZvhRqbcoHDd+6EMh7oHGOkax
ekKkusyGTYTaU2mQa/PRaSBVVMH4XsjQkEolE6jF7AGfRBiJD4AzyB6IHR32sGmB
f/7ri9qpPDQKxJUC+0HyPDRt5CAO0fRMUSQdqEVHUC4rLm1x4+6RKEkDUszMhvkn
+BvKItoGooKQJwWn1QeXyln99mJkSok/UAamIZm7DiZyTvuVbVi6jRgykW9KV6BD
H834ZsvrOSxPbDJZxtbkHqeMiViqMa1TgfGszih5O30lT1GBwD3H21z28PmDqvt+
My7uVwaRWfyC2x75jbYxYjOpjVz6/O+A/u4vXDarorwufWq7dMJ37vLkfPTtLAyw
VeGJBDGXLgtPgiTsNf5VzaYSI5ksYmCx7UVmuCZOWAa6H2RYCvZEx6BgJc9AQiW7
lsdKvG96g2wh9xHMwZ7UsJc/Sg5xCRSQUgQwqsbrTFr9W/HbjsSK6qsZ/l7CPxJM
IUpfqVGZk3c8cutzMsZeATjj3d5XbOlM/3MHqZ8+nc73IEERnoGy6RUioU+Z9Ru3
8D0ZeKTarMd80f5+VBBsaemv015xYvHWXC6+E/eZHirrA0noSrcu3LsXg5SwbgxK
p8Xgd06EYOKzIejDl0xFeKjeM3FJrXkTWiZFhkkmt7guttkKN+QrXvd8szESirok
1EiGJFZ3mXPf+4FDVPI7RSQUB/eQV0LCZewCTiAN7N5+XFU9yE1hm4mKy8uLRodn
pSaf+Rvf9C3ZCOY7K+u8aUO8ODvkzMQ3WeGuDMcsou3SeFQBEo9hxbBwHlvlIxrP
J5KATnNVL0Og4kWseN9tCL/wmUbGI7wUoiTW6UiT386dh8bMJGLLIwbcJKItywbG
N3r34HvGZXGZLBJlfYeH3xD76wGmZSChaGsVlVBCxPSymiysNJkcDf8K9Ebn+qE8
eKNo46nWIwdjk0LnPtkL0dxZFZIg4yR/YdFkAsZbffu6Tand8CDjN0UgkF4kTJ2j
ysm4s96MOeuH9TFQRYG2rkvDu/N2VmkAIsTqj++OprrvdP7Z6Pm1giBf5qtLTwT6
CmTYFyJl2ak3Ge7kjfMW7WWojTSKEyx9UMsM24HlYlZ0lYrBVOOD93lA0t8O4AkU
fbbRf4UaylFNKT5MEOKD9WvTCbSAhXpLKIZN4oL3kj9wFFzATnlD7EFuUMnsZYo7
euhsPKfTOSX9FctkW5Dkte9Iu1KFjDqXY7bdL/UndjEnyAbskzlMsq9+NCS3AWpE
9PoKS6me4ZzsafBdYDLMSdjE8L45AauuAC6ePsQJemmlTOVFdl0GR1JEjH0tSAiS
iebIkq1E2r2RSm2DRUmKunp0KD6JMvlwakMJow/Vfe/7bpy7qRaKML2JvjzbZCZg
EKVkPCLclSvTFVu20UN4l0Cyzc7fA6BaFklYpMbQP04EdjmuAyfMOukSQQOPUsJI
25ml+p6YeUz9l3LQQTmJbjnIEDBkuwVT8VvFSkvoxuFYVUnnnIsGIpPnPDuj/EpQ
I4ElSCrR6d7TKGYz1P6ol6MkPIcQEkCtn/YP+NLWzAUmEd3Tm6KLPw5gq9rj7kNg
FPfDXUZOYvckcioroNPdhNZeWlvEGHcZepX8VVoMMQ+id4bUsqnNeaEwLoKBOtnK
0QXWJPJcyJKj2CGUGZU1wFFYCniC8xz+Dh1Rdio2b+7QEBOhXv0cOPFpNYaf5NT2
dwf6S22b+T4CqOO+ssVayVr1fex0XNkH2ru+BL6wIAuIeKVtfvCGypySzWryRdGd
gR8vMwItqOq3hmsCBViBTBZgvKQIDSflOz0zwZtS3hHk/JQrkMzSfJQhDHbJwbO3
1mU6CyqgGGCXRuLGkVXJKcnjUmUhWfSlrRat8ohkQ8ECIjj25Z09CRgXZALMv0Hx
odwK/8u2NuV+z+exY2iZpEqxzUBx4r+2W3Q1xGkR7ci3fhrkH65h6W/xVCVX5iOB
g9u49jlencZ2EaKXEN8ZD3+j/441elDsHRCCB9CeJnngBdQ3u02K/tCNQxKUw1q5
oSJy2pdVI/hijj3Ye7ZfeKdyTs7xnXo5UcPj1MgVK2LaoJgI1K25BE0tJVG0eJri
lkXabuzkeDHEqbxt75e+UgJ/2fGf+ISQaa0C8WWnawL0r2q9P3rlG9TiQyUuYG3l
6r6QbwvrxbyQDngeC7KtDfeaLkEtgol9GcD31hsgKsYvCQv8s1tCErTifX8Bsqj9
k70TS8kDgf1LMaSPxpSOXMhVYFC39NkzeU6z6uXPwASk9A/sRvKMJu23ivh1hRhf
ZEbYF2tk8e4PM8YbuALH8k0jAJzU0NGOWFC/RnmMxqPKnrb5QRCP7VHxthh/RFpi
g4wJx/Q005oIBUbgUhvmApkGi8n08/5aoKn2ZOxt5XGmYn7cV5lJ1Lo2i0314my/
utzSybf95hq3mg12r8rsQKolY7l2qemILZ56RaZXH7JQe/Z3ZlbqTIhfx1Ph+DLL
ZZGLc4qkA55xtFVCG7iHBZbeCKnv0B99ZKJp+Lt0KLXkAFrx9cQ0MsZ14ka730bH
XG845KxDf4umELSTaP7ygZURqWgC+dQstXvCEZcC1Vwg+gipwPrnsTuDJPH7dodY
JDqElF/fTz3uQjR1yYLLsuvDJsvBJLJuk+3ZAy8iKMaQHdJlsN7V+26TKG4+mpIf
Hx8fPJV6bXj6YeP+wsLhOhp6c71DrZMRUNCjSiDsJF5XKfVAFnoIpaBV/nz6gQUr
FYftxmH/w73TZcGVfrf1GoTt3tb16FkMStVbRXicMVBAYL/gRFEdqEUh9fwMMihO
Gc94srvKm5lC1aLNf1vusB0gDmZg8uYHcxaEG5551y5YkYfW/p9l5h4+JsW8Ds6P
hH7pbESiaQSSaOg71H1IxGHaBp4QPQlyzq1wVHrBmFvAgZq1EaUN6EdG9Pz0FVC5
g7twbGXp6mId7/kczrRs7ftcbG/3fJ9zlfSdcTUFv48i5prrRkXlKEvUzCMKJtSS
nkiDPsBFTmALGvWfEai9nGTCiQ+3uWmP7q1RkO7sHezrjcT8zHmNQu60Y5yp9ljT
U4NSGMKI5atGMEXShImmB+jTcLB75tjihd8Bi1y/9D1xNHNC2QpM7qsWDU5pQyk/
zOJ2HFoSYhaQ8toaXMhqvEDreD4L21TRIG/wmsPXgkEhS37JqcgcJc4o3akMl3hw
wgm2qgnmfO4wPc8jQuD/o1DNZynWCiaRtnnphLPeHWryM0RdpFYlfkdadnYWzeQc
iWbwDTvG6ykQFH+I2ymvxHcR7kNFXqR1vt+h73cKTaGWELgdPW27EBa0hDaiSXTT
qIQzJcyd6Kga5xKp+MqVcxR3g4DWagT2Is0WkcPvpj20NdbjXg8kuu8cXKTHeFi0
lGPpCJ8bhC2COhK8v5ummnwBs2aPupj2eLDbwqYZ4YesPC8S95q1PRir+OI+HVvr
WGvvwKjjV6shG8Bu058HmfiBJlazvkfnRP2MhXCBoGL5wOg1eUiTGULdEOpbPPE2
WSE+vgp5t35Gtlf6ptLYEksRwj/oE/6hIZkk/uAR8xWICGj43y7ULKg6KHlHRTcd
L/+W2IrC4uYtAg4nlmnbr5BT8tXH24Xgm/rdd4xbvedsQa0L4Y6AbP2Px09wUMbZ
FBIj36nIAMnBIGtF80jqQjpo7cphMeuaInEgMUNezqwyvoBCHR1FjQJjwC2ER1V+
R52yviUPNcf2v6uV9JRaj2Bh3MUsh3kCczwyRKHlT1rMJYaOQkmaDey1QfwM6llZ
UswuxXGM6I4eqXPJpogLBGkoW7ceHNamclHSndOo3P+015jpJcfgKWEEGgy868Lg
uzT2FBsQ9NwgE6eXJew40Be+v4LNiqWehVPHrldcIEoJqtXRpqgo6I90Ye6ALIQ+
3EKdAYnWHVhfcZwn4QqJmngwNk/T1yVfpvgvaIBf8JyWWSD55k8C+uZjtzKfJM9r
5dr7R5j1ByWZhlrLeOVZKXw5eI/tV0c4e0eqxa0LXKS3TUW3UpLFyaWI7Mk2XgR2
5ip870IUxXKYBHAA+akLf3n7QQzXCCNpXS+2W9N6o53aYTx1S27aNbeqP0LLU4Go
dafeOmhs8HTdEeS41PCSBFJH8ZJ5lz95CG1b+rjdANK2KHjB3vBsRcqXikH6H6kP
EukdsFFJEaPRLHdE+23BgdBUi7bZNJirkxRqazgH1xMTa2/mtNapL7riyd1d7jQ+
Bf1Fglj2rbEsqk20kaNCgQbsF0g8sqO397IvkjDfZhZYqdKRQ7LBV3BWjr6Xlss8
sr/qWtRCnvZk0NeuUU8egqeJ3GvA8BT3a8HgYKo5LFtKl+6nlaljqkp6XpPfHtZA
co+6qfJPYlK/ctyb0VuLGFCHlAs0aYwPZnAo0tPsNf1I92QkT9b8paczJTgqfI2N
JSembBySFNgJ7uFqv1GZ22oAMX/jquZ+HHnhT7oMIIQfO9RomM2rRIGANWq6jVBk
d3767of+NTtaL0FOGdI64Gk3Tx/4NJJLTQbwPP30+ImnioMTK73bXy//dZiLo75d
ePHr9knU21eOxVqKVGAyVksqicPVxzdLRcP0ZY0kmfEtKg18zv3To+QH9DFvohpf
wW6p0m4KH5nGXd1IkCKfuH6utxRXnCW+tACJNknE0wgTfNvlLtTBcEt/e4P0/epK
owabe0Bafc5G5+f+Uhgqt2unP4EyR70ZD3TvTPqzdMSlP9As02V/sC8Z6Er2EaaG
DreJAv6CqzrB5TvKuEAHaC7cC1Pw/pfab6tpKeE5N5UhWqgMlS9G6O9JQIclq+vn
wA/Zbn2HOKlNEWlTzXY+C0Icy6EJhZgNAx92Cd6vy3zTMAzLj1E4cReKaeieMbJN
EQP9fY0DtvYbCBvl84Afe/6dB4dM6Ls1kzDUItUBRT3JtSo+8bkB5dzNpM7PemRF
fGuz9Xf1aLloSoaWz+gx8RfI5nIEr+gVdZnhRNXN0V8e1kbFefu4WOqn3GuOVp1C
b3pTIYdfsfNeMKUAfTKErs3uNE/y1QF1zNxHx6GJ0FW/iTW8Ge/vaDdrOBrnf+Vi
HcOjE/rP/De0fw/CkjnaHgesDIc2fdX6FJDIsQG/VFxtB5OFAOjcfD04XNDX9TDl
QKEeQ1RXC/Mdyn3M4wqzUrJBVk98BXR0Mc4Q6HH4nqfjE5w+TZSbMrsGcagUkmzG
UyVEgeF1DtJPKiFEfJB2DPS+0naXh3GU+B3mTeuW6oKkesA9Jr1H0QcA+fNQn/rp
365WiS3PNuZkfrsQZpuudN42MF+8v26TZTknNU1N/64q2u+AHnJhE8RVpMad1P0P
Z2qlLXSfLayeBgekVxl02C6AxfeEp+yguISBhPeAw8zIhgPEhOcj6GGjxP95bjXJ
pkHii8WRcwwG3TBNac9Cc0LeZTDpLxvJYQzdRNNe8Y2SLmJpKxSWuf/S98KePN6V
IoaOFj5B/Ixklehr3mhZ/36BakO90L3lUxQIhnoWhwqfx+HzUpvaiByOtrQ+MkWQ
Dl7IuITPVLHs33J4SO0sMUaHOwxnlK/WFuYMVHzmVLVie0L1de5gkhql6rkhqFPq
IPfXIk2bV3nhU+0vwkJoAOCpx7Ue2xGx4aqbxiMoPXUq0onW0tJ9x2iVIkpcvY9r
cVtIv1R3c4Nzl4qQJRmGvVoB1twMz+DeWrQB5xFjJD3Xsp/fQnOQZsIT2VVWgsiu
34ka670RpqiSoICPGthz6ez7hx2nLhsBCz5w4y+22LMho/uGy/jh354p1s7BJ8Qu
rGOINDfx+fQ3RFP1NDhocs/zh8H2T7lvfXNje1WZ3Q8jrOx3/qFjULKxt07qeBYE
UbvcerpDaVCrG+yN6uE1lhnqe5olIdSEXCuHVzpimEYpuR5roK01eRR/SJCypZqZ
iiDqA/wjVGAskBanUzjG4Fi1VG0xJk5Fc84zPqOKC+JoK1GLiQ1jhft39UOGDmM5
blcObBXIFypCV39TS+HhAGfpuI+1E6him22wJYgwqFPKabesMZohBHEsNLpfYWQ4
FScJd0RWrj+hGeIIdjEYkbJCUNsvoDg0H5EX/z5D6yp2ydt/O/zPpqK2kyaa8uOp
ApqznVHnSOTpXan3GPMaalpp20cKcgoFMv/nWbvqYRzcrY/M/MM07XWaQeVRWejg
dZUSbA87/obB+cOQy2/MZUJlD2BXu4y6Xv+wp3NeSqu1MYJKYjLi6PR4t4DSovR6
UPm+gYNgli/q3nouUKiJ46rMmXKE097SEKqQKc4MC+/qJ7gHBp3B52Sh9ypMY0Se
+kFYIqDtsgHqxTM/dhKAujChWuvkJC7RsXHx1z3EEOMVkt1TwMcjTqBc38vzj9Sb
Kdh5YHs2oeGgXeOwUulu1XknZymBPBTki6n64smcb8Sp8oQn5yZ+gBFCb4IZzEUc
1LddZtPq2F1eEd6LX/w+4WQsb3Jpg6ifVJLAXFFEZx5+lvvZWyZoaHlbEuhgBlk+
j4ao02nKbgHHCy+jCUKyYy+37OfXSU9KsCes3fx0rHtzduqz+dqcumzp8p/4ftiR
oRlhZNh0i8jfTkLUOGOkkxbAWALUDMnHPNixB7p9GmGh2ZFEZQMKyXnsllU19mfB
YXUtvbo+ZKKxTlLaEiMr6qSGxF1FhPD5Sec1SqJGrny0R0s6NvyXULK5SPtftSOK
casRh1Tu/fo/LLaaUlYL7E56TuPDy59NgLxdeM8md9W8OHKUCzWdgV4p3TanVn5q
MD6an3Dq6hoFyW3eJkjlvz15g3gaRgKQDXD/B0QioHLwXRjxJTSGG7b3sb5q5xkJ
6e7zSe1Fv/arZD3CzdWiwd9Yi0nw6xIn0KeE/lfsf8wa0iBD+XitnoHbBONhtmyg
gzl8lerx0Nb4qiX/JNGFnOtdNfPzQoVTi46MU1piMRqcj+KX8JbK7AiVE7o6IZOI
zOBzPtOfl1OQ4TXoh5AhVuZrTU9pVVl1DYrLQthiZG9s8xXqs8z89OoFJWUf2Xz2
piSLKnoj4TPVImuwgip+WLWUC/tCuyswIuQkqXCgAJpv701V0lN982l4GxtaImnJ
RCvlooIkvpwBcI59nzniClPx6OlptEaZJHhfBTet2skOZpKH5qjCcB8r9JJ/4rmj
5aGTRgj5y62tnkfCExe8UQ3fHuQoZQMT2yZlr/ki4YRdLGjbS7prov6tglSr+r+j
NU52jyWNgqBwpaDpiyfEBYtadAts1Y7kKlyMqzPIaUrdPsrYiIIWbKpREnNOCnY7
a5DXh72w5vCClL8kZkGxFbd1vc4oUdC5fee4lwUYqZ+QcZwKD2Tgx0BCtbHIexnj
QikGXa6ui0gYbFDIZFVdvlTpa3/PurBCen/heNe6Zbi5Vx+Lf3uYRJvghFT2yC5U
HAPXTAqm55RELa1Wl0XjFGb+VqvhSfjF+Wz9970VWsGUldJ/r/CyFf7vqswM1AbO
ySoxgEFax/pTHD0TnMMmX1STqYd2j3kgRA+RPHAPnoJiNi/GvKyepNx6X7rUUejQ
GaARPbSyYkvJ8c8zJBaidKZK+OOXzwkmBx7rz0BjEqDK1xDhxpeSvBnqBkEcVlXt
bK8nW1AJ2sNL+/86rpf82IhHbe7B0QL7+MgD9u8YTB5HxPOnhSJskPJ1I6Ca1sqr
85qORxm0hdEqjVgDw5R8T5O+VCac4LWoVaT+DPKxoaQ9H7eihidoMam7ujpTKLso
KjKXn8sITh+UBeb9/9lD+xyW324/qXltStarcz9toj1RfpHKXkfvyetWr++IU0hO
YTbEi4ZvstDF/LwQQ3vIwMVv4RTukdgXB77LKmXCDP3l3xDqo8UWNimAbSNTS7XP
Eupla/tFfSLJyhfc32THLoM4EKZzI56pregKopp56COPvDnQQ2NMU5xyUWoGT9rU
6HNR7uVHRzM4xhJ8wHzoLVMN8p+gtnWKENHaHsDJ9EdHmoYTdUeeL5qmAhFB7ejh
cIazTJMYTJIk0VSkgb0RnznGDTPS1fKIQMN5WxT9OrXTzKfaru5cx4cRHgtS6nMd
sVJOKf2qCgtHCzSsAU+77j8uv/qelFHL+WTseSB73Y7RPd4kboLkjt0pqOBsZuf1
DwsVHw1kQiNeFbiGli/aZvGhv9aAOSmxIZfPr2w4nbKvz5PX2hok+fhrLcrBq5aX
nws+CUvmm9pVjL7OxPXtiKgLILklEMES9isnqz1zLUQcpdpcknnxix7O9IrQQMLQ
Ywdfj33ggWi23lcjlfFVHuoeQRTHwVOJVEVCsEhTEa8XGdYue/2zcnpeGxRqbfKB
hgP8YVWSJGhSvOJxKohVE+S4egbWiysaFmJEvR9PWseG+Px1bsYguIJNUBMySNko
D3/F26P/WTf1zqNN5G0RgEWaBpEx0YSABHuO+Vv54g9nGegpWiy9lukolyTafjsP
1O1wcav4l/cEHKM5bMad+q3CXiM5mmB7B3zpZDssA2eGjHaf1YK6Pa1dXDT/rUfV
OvUBoI72CI46LPyktbHip6PM8eat6PgyvQiVkRaAVEcDIYdag1IZDaxA2watRdAx
tPQ9dul/keMJvWj8UnQ1oCZxtkVptMSw+goHNAJ5It0Y/45gtZSfbpVdoh1kBntn
UA1F88zYfX4JoxclhrQ3fpO7gqwUGNKHYq4bCTiY79CJtTlwC8r2J6hovAi1digF
EHJDytfiwDVu9MgSAJ9dP0bBoNnnY0NHMBSPNWAdbmhti31Llp7m49UdUefdwsld
HM3FjdNyrPfT5JustHK2e6qldYsagl60GjW9aG3Ft/koA9XmKgj6snk1IU71CujQ
Y1yk3neEok603p997vCwENZp08iW9zVcWYaqjuxN9EnAlQOHuql/KmAzbANkfUqp
93KPRj/bWxqhOxe9+AJ3WK1qWDdaC7P91jSvrZDNrrgdhT+ZPLhVj05xV4yLHTKB
vxZy2ezyS9LFMmpd29kIdA16TH0B/3k0NAealmfrGfxRheHfaGrfkPgRRNqUZ/Fo
lwbIak8QDLSJR9iRJsxYTrlI7Fvg0q4jN2b0EbBQBFlnTo6nT1cNx5tclS0uRD6z
7jRxC3ws0KoD3pQBKKBEp8P7Lww/etMgJdrI6iobuwJ/rgL+HZP5cPSrftUTJ6Da
GMBZSP7pAShe1ZwkeEYFOsH2mljw+8opJm4NLCOrL7nYcIh5sDhlAXZiOX/7vI0N
OBufePWYL7ls5mXF8t54WJ5fgPHk7pXaU0QK1ZwhbLzJJIgYjdsVBFawCOdRNsui
jOfrFVJbVb2p7zkCrrZDAjMSVAFI0/PwQdPS7eoQEXBoruyROIU+iC47BzRsw2M9
RCuLeQEyqjR3eHOJeUH0LrWVi7viic2zPIC1b2mEDYpKfQ4AvZv4AErldmu2CT/q
uR4CVv4sbbYatdXJKq8gAvfS45TBznB2CHnABKadA1G9mVKiSEENNCb4bPszfvBi
2H90o8jH3Chr3EMfrG2de2D/5c1DzZPJuRzAi387qLS92n+O3W0YFsPW32AX1iyo
pYNDwNFkYd8XFitK97O3HtdFcb5eWb4BH7+uGWeof0E+/uTVf/ldo5UFqJr21LAQ
vwveyaky9kpXOoPt5gPylaZ8WxWl1wcT1649OHkX25DJUVDWsRcp15kcOucWTZr/
RHemlx3kMMDQ7lexxWteMtkxBAUsTkd0CFLSkR5NHvIFQ9JhfIJIc0U0L6AFBxDT
ZMYQYFYuvRmz2IieiQWWZxfdroRScv1G3RMWajRrHewvQGiJyRWU/xchvzMYGWSR
+qSu1PbADfUKt43ZIXxA1x0hWoWSHXT4xE3BmKt2Zf7u9LogN1ad8ia6Tjtbc7yc
LhL58A62MTUJ3ovi6Hm6ou/g9HZKNlo/GfVhWSKCY8LKNfCPgbGXSMLexbivUUt1
6fWD5SymLj772AAmPLKPv5xcgpTNQiXzWjGn1B8KNDZy2xusPl9xI4kb0AxZLsOM
VXXVOBRlFUVODUqWA/+qw8diLJQS1ys/sSMAu57XksdrTImKu9/5cXcrQ3ZL/PVk
6yDTx8tnnN8y1n+KIaf5z22t/dgWjQpj5H0KorkV6wWCJY3WcfyzVL4dzzyXKhMr
utH0PcEMyEqi4u0XFfi6MdQDhVvar8M3WYnfYFlhNpbFH9LdjdNv6jQzDn2rBSNm
OTXyFo8WDcxq+o22VKc3lBCt2QjiZrtVFQ+mttZeN5vFUwfn2WU50BKKObsCpbld
cfMl6fY7frZo/W5rWY7law7OIg80+JZjmWpq8pQreh7AWqJN3yufQGTCUOlxrqbe
QQr4DpAttMNYFvRDcTdmkLVypNyvu5BEvo5WfwQA8PCMVpyIp4OXMEtLdbTCNzgB
8nydc9ihSS/Yl8I1oXsKRoSAmpdkwDmndflSNwAHApWeKksxnGj9mvymw7mK5Fie
wMIG/vpc4vrsOxiEonA7r4MEYXCkKMIoxtYhQ3kcVq/PUDaWtYCXGV1CGvER1h9k
DPOc1tVm8MTIcx/tRKHADcZ5LUSB5sFJKrTW9dNTFqLAcSX+f9t0vX3wAx+bW5rZ
pNi9N9627GammLqqX/QGfal7uMOk8JeWl4yowop/MKk7jGpw/ISwbu0Tsxr2P/bJ
67Wy3qo1JidjAq0k2KRvor6vE9q8TfnWCa7MeC2TT+SyPbnVar1op6OhiIv6hCbE
WbsrM6z0SwHB7tKi2425Q/HsDLnUViXYhWQF6IxdA5p8dTKdHiYzq7WNmI/Y+Nr0
ehF9JXeru6TdyhM/m0nNUOu+iS56jRU72sbyHG7JxoJHICwHx4W7nnULUG2wKYwI
NTJq98Ee2H40X8sfTLAyY62vbM4IOXrfrGfb+u5bw4qDizL7n8nZOqdMsAwPnvGh
i/4bA2JjojAeWYHCXJ2pWmera5pmUnSQkXice3Gw9ROB4IS5EMObiCTV/zYZVirQ
5CcpRuLBBwiIOefxn91poWV9GOs5pTX8Wb/4LDJn5j4hr7xvsACatHJOWwXpuxkP
iXI3tYDZ1xh7IueTzy0nrzJ3MstkgJqzTwmdhXA5J8KHkq/RQnQfNVy3MVHj/sly
Oy1cdUme7hpAvdkPQL+KjCKpvFnQ9sgMJMdLqIyJiqXjd4QbxtZAovKz9lvOp5yB
VKqCSVs+78Dw+EpihxJBdQvxsxwskypNaVjwD84EH3ZgXD2CJ86NY/x1zjGem4jz
3PGBS4UVd9bUzpyxGxPp9ZO2xPziH1ydc2qDSorSgr1H8+PFskZeYwLOey+a3aXZ
tRaM8uAuGj6pXrRkKVVW77AfMKtF5W7e00ECNPuyETVzNucDrSN4iYllVhmNs0a4
d9phIr3UhDbazPyD81B4fyL+LOt0OnKFTWkQvzExhEiheaMXePMGbDW/QSuoIvaG
bxjAD8SVuck+IUweDb9dO0BUabdtICVP345iqiNn6Pf1IEjvPguFy8ZYEKMUtG2o
WqOHWViOGNaECLHncLVX8j12cWn58IyGgDJYKXH7O5HW6Sepnt3SsUve2gSeNJEA
SvKJg0JnI3smlPdh/sCrm+Ww0lniGukCySWo1168IJB6R/OrZVmSXWHVLNgtYxkK
LrHkOpYpXyQuvoMstddPh8852L+49wySvCV9l1sziCRv1lwO6oLfqhVQyk9LCF9D
dcHzbnU1GiCNHQHzlMW/IoEsxlIf7hTGC3s07xu+IGUSyl6+gPddQgFCdwzq/1Ro
ACUFHVDWt8zjsnXT7b0zi1QYmsm+zcs+UdEjq94yAPeTSHqlNiCfoidXJcdO7zPt
GTII1s9tOB2KmW0Ls7jvAxX3ELRQJU+10OyqMBmEDcjrJWR05LTi0pRUWS0zUuFx
9lCCWJiE46/f+ibjZuwVvhE+UpuzOZDRmp559EbAT5nPm5b+JVvo+LRqZFDP5vBS
FYJNIKNGqXXkuGALHY48Az4y9BSyBNcESFCG4tE/D56V9Xaaj3OPHFr21kY9hbUf
WY7tbQjEBFM58Wrfvd05+ZOZqQJtdO+HJ0zkYM0TS01j4a5jMt4JTArfM12a6bg1
6jF/DsTwjVeTUtZTJPk/BGfDDcvbTbpSDKDvvaEw+CRmlxvtn3mwYwRBl9OXWuZP
eFzID51Q2U6UsAURYaUFIaxl03YtdVC9KM/5z/u2GXDOMH3io+wmIL6pnRVzibcI
ongCKC+KYGEWk8X5K6146r+J8DhDfb7babt7jB72p3OWDAq8/0MQSa/ZwL0N/86H
15XFkZMCwMD12DKSxbvJR9MIdDrwFeiiMx/myG8g78TtS5a8BiQ4ZSpiXeT83kLd
/xl2smARBBEy8oMWEV6wUE+iQxBzGF0cU6ZsOUoRKvkQTUWPnPIaDkt81qXk8WIQ
NaELOYHKdSBXTw9EST97cB/36Ycj1ZVVGbNLjCePNnrUU5HFISH01ZYdEDJqDICb
eQkCCOeX15lHhhrvQm5DCG1x9XmYrkxDkPu/O76SOpf3lyIhxpSIjtQ0DmZXQEw6
NflUQ0L/PU9WjkYnv63VeeGefpndvYJJSuiB+Mb5T0vcb19RJK4cicXT9o6nzrfl
rkya8/jEgC+GfEZypvnCYZdEMXX7l+eO0qR/2Xkv6MZDnkTpNd56SNObiY05bVlK
9cZ3EcTnH1ujSjeFRSI6MV0u1r7rXNOCGYFOpont4JQMNIrSY2pf/EKJyco8iKka
/OFbEDyiyqe6+94SZiU8rxoZqwyhnEGwkclArvnLf4a++Z+XW46IfSiAJEXn8hna
bKDQVqbpRhWoMmxMQ8QeSELfUDmdrvrZEOxmRrF42QCLcsjqEl9CGU/h79rmZO4M
0AL/x+qyrH65fClZ6T0LhpSmcLlfHWfwLeMhyJuf0//QXvo/MjvjXxhSeN5CyMZw
cZ08dMbB0wX3y6PGf0YOdb7bUWJ9+V9NlCNvGO54tcmHN3g6CSvgRtudPjFShy8O
wEgWchea+9VC64XGI+eruRMBLcXgyRTDCdv4Efw6tv1bRs/HW86NifwLAJr6OX/f
CMJZFcoYutgAojU4AviFGq8K7QbbPcr2NPwmhaK7tCTnhRK1hvee2xe2aQ5ISLR0
jAni9HOFgmtTx/QEOPR+/71hDurU1ds6L5/AveRhpY6PgMc62TO8nLgu1XWvJAfB
ARw2RLkZjxfVX4dyjnqQnMYzTCtzzV7YONu9xWRiHK8HpD56clWL0eUzjQuqfpgH
PkdilVnd25mycvGNioR+c4C88Q4rLV03855aIv9msFo01VC1wj2+19Z7FOCGLsy7
WOrQVFFkDBxG2Sp/6S2Jr9TooFOycIHdWshLRSqL/y/GGEgbDDu15abrZlxpGvIW
7FiYQrkUH4oIcOzkpGlQ0rkjbYBzFhx/DCPW45QhQngDlHnC6ffSEat1AcM3Fcf4
liZFXjJNjP+WnHj0gTYgErPuP/wGlG3k3zYToiGIv3z7gG38dfRbplAktfnpU23N
sFrA7+EUqRBoRvjR52pMWjmtYOYkqfu1aeO/e+1QVnA989lS8SnoSgNvX9KZQnaI
WJWzWUZd+08f1S4sOgWYYwPHEvlkjdHiTu7Xt0vSTH2LntWRGi//nAzmwxyOjjPm
UZ8oCcQV05w+nLE4UeTfU/XU/Tp4YzGh3LuoV3u3epLqZSc6TCUeFQE1/mSbcwmJ
opDg63pjRvWGqcK4mJsGUFMbQAxZN4EzhErMDL/wx+W9T2pEJ7tw7Do17XqYBkhj
SXxp7kTi58xBg3mrkjLknr4DZ9hVply0L4bQRCovLa81zi9gWk8tamikTloyRbge
lB+PwccNAwAVO+Xo8QJTV7ifJ39RHhl8JfQaMRzETLqRcP/GKREOHiAatSeGNY34
4A2nyK2nIDZbN7NAZb0mPQ+mbxUJaIlUuy8qQBtnIK+PbsZ/I9qaa2UMvsTnuJz7
jPbv3OxdruTRSOlXElJHsBkcIDQfKR5uWMAWRlYrIlgi6sUo9Er0bXqjdXkpr3kO
izVIPqm7EshX8+/76BrzHVaKzegUcBmk7DcwEiNVq2fLYkXNJlCu6Rd1s9OlLKLp
079yCjn0JI1WStiOgGlMByU5d+fCYgq3oK6eVd1JaTaVv3jrPlA9CxizT5kM3jcK
GbIo4D/lSUtDomxuoT5kDhMjrv+La0b/A2PKY52vdSGesH2gAgfPOvFng8HUyuAz
1gmlRJhDGC/NxxBpG3zergaZLOxxoeqsb1QCFkBvmNs++LEASHXy5lgNFrbUZyc+
PQ73AmdZN7K5N7WBwfq1JMr6revuldO/QUc7Z72uRWstIxQrRlaOVzfiBS+j/7vv
zlRntUpOM3EdtucsDPWa0+JjIjHgiacubnbeRMM0/z3SPLxNMf62zsGrM7Ytm9hO
Xd5QsigiJ1r6Xaxz8YiIM7JMuBNuGcZD0cM3kLlDA+aNoaaIBcxSLQ7N9Y5355DO
+byqBx2c6N5hm0OofopeVgFhSZ72DegBfJv6FwcvghnIQCqhrqT1Rj7OknNUhyHT
4jYAZmnXasxXasCg2tHuQv2mwkdV3xOcPuHyvJfOG8wqMVfr0iW6LHdGnT7W5ztH
N+AT54nsyKKgAfQ5vDg7lPCm4qM4EjCHj9oV0ItEdhRfD91IjQB74//JTzuF3r49
4kHWzFp0Pgryti0NVmLQI4E1YevVXTR9xV1JPY5YMQ5IhqyNQtGWifiuyHK6z2gs
l8eTeme+pDxxhOKx1B8olc/8g6+/hCL7haZnVR18J4GUhLILjlCAVGrHzOW8o6NR
TCVaHUE+Ro2/EqKpFvIP9KcaLLr6JQq/yQ9QlKChmZ56l4O2zHAb1ccksc7ss7C+
7rahNV1c/kmeW2XNDP2VifXyjFcqd8dAk0NzYeVQCUzgMXvaEaKfcAKS3j5WUHlo
mOuZVZMUfGJKTusL8YSPWAYQmGgwZgj2nVpX18430rFRQKC1RN2b1PRLYfuPXk2/
5OTHO3xEdOOzDwXAsGGo/8Kba2Tajq3kVH0PJUZKB7eMECa7RO5K4XPqKvhbOtWb
LK2mT3p6CB+eHeyvsenyZCAUNWgi/0RcrYuSPWN0u3WCI/jpmF0yKnwpHA2uNQo2
3mc4zaORQTLrpCWGFXQKgV22FtSdR7oKWCdUvECwld5RHO9lXYf2BLCV1QiOOVA5
d/5oe6KbmmED2fg/l8CZjXqeuX/foNzXyJ28tY6b145TSYGa+egdgmXcUm9iow3F
v+enU5mmDyquVke3iPqRgkWiL05hvhNy1zYnhA3W3c42SygifBrfS7DWb0t6s46b
M1TxXmk3DG4y5zUrM1HyuJN78nc7+SdihFw7HHMjnC4sR7V8TTcuLEMneNFtbCwJ
X+obloymEWpCYx5QkNmf0esTbCKhqIz0/+eATtnxMjkiYtF+8DFv4vjOIEXxGHF/
hsuomyAcUQEyXtOfSDKp3tkWckWjvRzlJkoe0WuUQXjLfYt02nKfmtU2mW0J9lbT
Zu4bHQLq6uiaoXHkls8NNRpXK0GDW/o8SQTY8PYzG6b2QqehJLBY6od7K1255K44
/SOTxbU62b0oNDql0A8sl+hVd1+rU6dc7pws1ch0866/ImRpBRUhtTJN4BStblSU
heBQlUnKLKsFufjX6jdpmFU2oiRbmfyTf9olW53OiOxJgdoAwhd9uiY46r/ultvV
ywfqgFxFIBIr6Ht5LGLtiRPZAJd2l1ruLEvh0ok5BNaAlk94lhdYq7EPRcE97ZCQ
M+fCTi8g+a/WtFbWkK9MriDsQV7Vc/RA00aGL9r0LrSosL81Q22cUo/+g4JPmO/1
P7JmMOEsHBPi1iRicWlwikt7DHbIiXPcps0O3+BmopiNFWavp+csbuIQh2hDG8LX
GvXHfuzs3tdQ91lwxtb0n9+GdpEdhyO13F9buiCljSnWjpYEc9e2uH6R27V50791
vM8UWfGM+EbVwXwFHZlA3e+yaMH1IK2l5e7N49h1xYfZIITbZ8AoEyIGxvepwN5w
EWTofw6XmvsWGPdIpzFK/Wb23Q8uATuuXzBAnAR8i8FV0VUHUF7crpd9WgIHIpz2
1FZ0aVmqs1tQZfOJPoSGC6eYCQq+4zL91MD525y2+7EOjIL/aFlpBNY2MBWQGxiy
wtzYNaIfovpd2lhOiYV7xASWA9WtVCiKPnUY6ur6gemR9zm//8RJuHtWAfT16apg
o14ONcWbdXQ4RhJGWnFQc3OzuV3+/0ntl5q+QGCZ8PiWbSIxoGZfLtff5FNNqs7Z
ZlHBeP6iKhJlAaKWJNJ3krbHp9i94t3aBHT72PVhtN3IwydwpvesmYUn43wMKywP
a1zbsykhPrNeyVUS5/ELwZ7StLu66A/O53xfJpbPy9aesAT4EG0a5Pf/YsOxQJnf
+BhrJ9VhJ8frV3WZWNEk9+InJtdTdulTGvyJ70pRKB/9mOw4rUrqwaZZg4TZFwEA
942AxjjdhUN3jWt8KDvqtlTz8TQ5kSLEH78+1++hwZK9INYL6F8P2FWtmLNlT/6d
L53bNU0gthwYD2MX57vjeVzwN7kLkswLKlbPvdGndjteRRRJAomxppDkMks0IqX2
WFINzzvpl3KHdaI1n6J26vIpTqB9spd/IfqUNFP5gHkfJk/E34UyEMdVBsAi+72U
HQcU3TBeYwNyWSSvXoVW7NWC/EOff3GSaz8GI6LXC61qFvpbty2DnMslhpPerSUo
v0qvlYHQLfdDDdnQkyuB2xsENNsnDpyYJwUi0OVtonn90XlmMP297awbqCsE8qgw
fE0HTVlAgXWXUUKQNE4QaJJYVSkxk4/l5ZlDpYFUfSkWuYgAkyGJZRoMHS16qyDz
/yx4+qo5DaN5q73cvFhehWgt4IdMm4OlRIOCC8CAHIBEbpVWeb/SV9lNVTwi7iPG
DOY0aEKLEyS24/pmhSfqxivegghwP8C3r15ArOigUdMAVOSjJiE5Gn7PmgEERXA5
aXtZfXoFq8emGa3WE0WUxg8c78ovPGZmZ/5O36qVMaxh/tsgpz2GSXb2uuvd9la7
70719UY7VEtCud6VnygUpozCxlteWw+ChoEWOxmhKNmFSe1LiFAmVybK8lIQf3ke
HKywuQ8Qa7JrjYNNR+KIcKJWgjPF5055uAUUyu5IslrkBHBcvALj+5SUv0b/dTZC
n62WKgHCdCbF+eLGAqrQ6PbzH9NvgH2ZXKVKjxrs5oVC9zln1AWPfWYsXB8Zrpo1
BkqOwK/1EjgQe1jseeqEdRLqHaTGaxOQptFNjPWdDW23DYXNOpamrNQOkEthx48x
g+cvDqPjGVNpsB06m9IJaMBFdDEZotP8p8bwY1Zz1qR85O9fu/uT12CqB1/Xnyjj
aIj5RxxkmpqWDZhdjHJpdauvqgCz3p8G0whL7rLZburk2xSgdowDZ9b1TVf4Pywb
uXkAu09Ntcd5opt0AG6XdZSw+xZ1Efr9fyF82K9FTzd9ZaDD8/OooCdpqWhHZ69+
te6GqoylQ+ZJhZamLT9hgZ01Qa8pCP5KkIYCkUnddZej6V1XqE2pnqqNjxQNYSO9
DrrjwKi+QIywv8p6Zgm1iKCFN0u9yRyNGAMKl576QeBOTprx9trBvdwHCi4U5CKc
L10iaNm4LEFh/9Lha6112+TuGwHQRa/tHtYWb8WhDkPiesG4X/vi62Bco6cKWle4
g5GeVevBhxg4kzq3dDVD+4Tj7lM+rVZACi3YIn9vl63F42fEn2YOgpyifHRUwoAV
4Hjh1q+YLLJ+abG3GOP4s9gmLlOuAj1XLdoznYficaiiqEkelCftD3cyqNgrXUeC
ntiTS1Yp56waD7nsYa0FwLX0GE2nGbx8eNC3yZsrPuceo2EW0r20UJLHfjmVVqOu
HRRCwBK7HVdtmH5dqDqRQtXwpbJNf2AmWxWPrjxCkyquec2G3v+MHEEpxRey/5az
NWyJy49/w9UhECSYwxeSPnB2+p5ZpLyj3zloST/AaEUY5RWamVyg9FV+IAhVjHVE
aQq7/kRnnvbH2JaUizlGjKpDueEQdMFMHk3hkQnwkueczqQXEbLe0KztayteyT4A
AJOq/mRJ120qrTqfBRW9T0gEDLgKTequOXp44cLh3xg7e/68T68ujLU8DTVQQm3E
a/4dZvCAxn9XVRm/hjb7nt822ReqH85cX9KA9a7nviBttRNO7T6gK+PXw/U/RVXx
WqqqG+AgexD+sZzWX4LVryST0B+3HZbWlI6TDqyvvJ85Yb9ZjIMnOp/EqM9IS2dL
9vFFBC0cNqXixVhmONV1Xe9+1crgD2a/C1Np8LwPFQjI9P1YHptEYwJuFqSAwBDI
iIc2HVYN8kENmAblrhfrQeOnJfqA3KpeuBArTLCcl4VpJrXNCCtXYqx4uO0fH6ST
s2dYLT0xG+BB6unahiy1b5hBMwR9SLDreXpDKmf6ocoMnFkSXt0KkWP5MHFK9Fub
FE7asq7Oc6fMGZlQBi7skoBah83uE3CqilIRGOZngc+cY4lEEUKV36c6CHRZzIl0
pJWukpvJ02TbxA2VE9+zeIjJg4RgXEQmY17Jz+FRuVZUitNgtATTf8BexHCxBmFc
en4ODzBYHi838f6bCHIwjwU0WXwUm4mMyam0WhHODS/fs1DetAxY0WgOeDx3Vtks
j/kIFUEht2Z5PAuHqT8RFyDZtC/srPBPPvGi4LwAfim9VFi/mLMBcEYYrD9aXOzK
4ZR/XQ+dTXwfuzaUzK5SK0CwWdW/O7CZJbRkMt2bAvAXNATpgH/AYbF8L8rvx1nS
iRlO++vww0j+chvuwteFZ0CvN4A5APbSVXHjtSLF6Ncdg3IeqnJxBVsShbegsyz0
jJW7M1IjNWJvSY4CS00T8poEiy5GUB6n7nTxpFjbZxnw1RgxeF9+P7oUZ+90ZJx5
smRpqqpmzIExefNWKXzXdl0Yb0W2u3bNUPEPG2sF29i8mJ4baDZbqf7uIa19JRz5
deonOuR7cl1b6vpS1OUq583JXb9bTHvKTi8XAOilSuZw+fJ050UW20VazcitvjfF
gTEL4z1GKZPyTNixGIAM7T+qSIinG2wbfLbn3zjRE7lmzkBcPg5ZqiXeT+7nyu0r
vl/W6/uZ14PIGKVQks9R8zZ5rx+Kg1qYmJ8IQVRwlZ4x22volATmfwmf9KXbxcAK
ylirpCHFAav1rQR8hq4yXQ3eqZ8hOSXAxnCJOQAYXCilgJDhiGWBK9HC01PqbZzo
0ExAanleON3VD8qebvkKdGFxBJVrURRQdLoAyyygNwqXo8tMjb+WP+/4QxdhvzkP
5kBl+L0ABtoiuKsDxYoVyaAO1pyjqO33tfYiDQW5i0BHoV+xnkKCHWSBoI3sqpn5
3AWbAWn8MCMunTbGF67M/M/2TC1dj8Osi4PsEQME5/uKd9raUiG+zQRNbSKn9glB
qp2cwU0QP03p1ldjq5Bxz3AoYfUyOXkH+i9qLpJKbxCEffAv3SLV4XzL74mIHBhj
nzvjLireZGOM96ybq5n0IBlyS53zYcrjZ7mxRBw3pZZhUysiZXe63nc/VB0HK1cZ
5eqkq/1UrIWz5vG8+eA9pGU91MTm5d+MzIx8UZ9HkakmC7PQJxxYTomc9JStrSV9
egfwzZyN+QfxBjkumtKmkxc8PUv0lkbsDqOy+8qWw4hwZv0utqPjTMXGdB1q3wMu
pCZati7K6xt6O6IzbfVktmuwlxfoiS+wcoH+xiG0CkhP882jnOy61F4QQ14QpuOF
IQeq25aAPAI8I3vfZxD3BnxAsLBMDMHr+IrcpoEGN+hnWZPRywNiz7VAaPO0k3NP
CK6zNOYWZ4B5AVCYf9sMHRIrSYuyg7wdvLzCphN6vXtEuFodspsATxcEZhGchTGZ
Si/+XfzEbVt6rGeMQwVG3yBpU1kawq52S6npNaOkWvKIfnTlyhs4oIpqRZ6ogQrI
3vQNu3m4JR+E4aWg7MuNVEmm1Rl8mHYO8/hzTAAkJDQJoRXeO5ECnrN6vO/HMYqN
6JsfwHLfB3dJrUk3g9ibOD3OEeBq1Zdkw+qgNoxrNnhAsmgFzyMh5Go0XGvrot7K
phqbZx8dgUa4wBwjj1+Won94Mmx2e1XeixJRO1EHRBFz0xJmPjcmDuc7Y+XJyqkB
L1Nu9FqBSJw6mVTnQm7WTn7V2pM3AvmgWj4d7OhY4XfFjIvvc9NfpPApEOxyiyyl
5bkZoY2E1x6CytmGRvwklEk0G9wJx58WdAhlpa47Y+SFNdm7T4lPEC2HNZBMQoh/
LA3eVPqKA9BAYoJ+TWJuh1uzmu7OeanhsItd2fz2bMUqiHLOzVUk6CC9tzaMq1f+
CtS/n8zlq0nTo9rfXKRiHHN3lwfQfPjr8qDH0FPieaCAa1A7xXsvakOe9sEjz5ZG
O7V00aM/5I/0A6zhk25HitTDXBAzybPbPy+TYtwuU1L42spn2u31Fkw67MfWNm9B
cQflaFyECYmCFGAeNGjDC4yW+/GCp7ijQNl3kQF06CU54ijWAZlWpKfPc68Hby3G
xjSeyMMe1wSXLmNvVvdgFVREOM9QzlRqoqAzFE24AFiQX5rwDOv/CF1Dg97BTGBB
1QfzBe3jM6Xx9LWYUrrZwcEnEnQ2ZMHIFUfBN+Z+E2Rf0tRuMORVf9ZcrnkOAlrc
BnM2bb4g6Tr3cCcHdcU1e7HYSw3lGiMbV+5QO1awyq880WUvK6N9LloHtCydWARS
ufJeY8fv8viIuBDhCV0W5P988ClmNyoAkyuC0pHv5mavQ0SHxd74dsparcE20M6e
CtntWcmfd99sKj3cP/0j8iOIdgrvt2K66u1G+OLS7voZdbMP1QujriMXTDvrEF3m
KPSoFJZnXbrV89DhlhCu6k3kISU7hr5yHhfh6XhN2t8VBcjx3PXiYJSa538Egw9U
l9Fe9QIUZ0QhB3rCSDL/lRCbQP9e9RzXt9pIjZeBvR3ZwpjHA5L8rYcfh05HsamL
fpIo05nrF6GUEntBKrdC/SuOkbw2msbXyvirl/k7rFIyBbMPUl6T8mxWaA6dgnHJ
RzmQP23M5gdvHvdZ0Z8gLr5PAix/AmJHFYhki7WspPHuqlaQGtFbAMJDAyHBZofl
eW8VFukrggId4eRJSr64ar9hBonV+3JMP33IM7OZFBWjTfryys4ti1MNbfoeHHrw
mQKgnHyuTiwXwgHet7tAI9a7q6dZtIEiiqwr/cf7SOlkHcYvl5MI1f/NsgL/F+Py
hSSFD9Zj7xzuOYVMiSVePFNMFIyi+yUGPEY+whEwOO2TSyzlJcJsYaftQX0c2mZ9
1gaSS8VoEvloPYezMJzPPF9Dsw2f4+j7CLipi9cG8Z6KVdxLV9gST20AQ+iwJHcv
go+1FHUiBnELjAVTVfU4edIdNrM2hJQqk1Ou+7FUdlQQioX4S5yH0Vi+mCCqzu3T
BZLkW56IoZbqBBCp8cDyg7AMAgvFHcmLRhyADshrbPGzghcTWjvtYuawE7PwDVMQ
FQoPnx4zAhp+WZg+XMPEooC3X3Uxs6RGGQQVwscl3a3rWJXGO6RkLdbrMBnriWwT
uIWZjd9e3V1xtSvpFMd85NW0miphvtXZ1DaaQwd3gs2UoXYoe25SfvbbBUZ3Prbg
HU9nBZ3kPTSiCHHMk0pzHe2MqGNJ+HMGEwhyVbhWLuTK3tsS2pUx/FpjVlpbn87b
PnUa3eJTKO9x0heLfyklxcQaLeRFPEVZI9by+51S1GErFEqm4pgmwrE+m5wimu/N
JAZ7MmnO36kxs1K/Oec+bpWIoNYpz3LRBGDAqciJ82kx1uNJn5CL6DCTlrq/+f0F
koTuTmawwiIwKS48TOxtHMH0uBaTNfIzksBRaffpMRG5AiKqFmlISYs/gvHLRDbI
rWHqsZa1U7/ooTHmUimQ2O2SNPlZxdR8/bN/iEJW3CS/HsscJEcOL6mfaq7mYmkp
IUDSFK7+C3ZljBPg+4BYiH8oHvrAmo+OgUo+u7VIu0ZXGPPgUO1rt7XeAlWIZZtx
V6dPYtljTa5fCfJ8O5bZkc0oNyws5YtgY4Gs08YYD9WT4q5Wp4Ak1fiRtX6fhWbl
xW4mzcgReL7B4nXxD9yCqkQ7nzl520jz4+xXhpzvTuvU0UW1A5LYYudYETVRzYQa
LnfCv48X9U+bZ2DkobGNpw44mXGJ86IOeFJQQVPQbzTbNNtq/CSPEvhy2CdVpY+g
YXEtTD+HL0i58yMG43P3Cne1YoqJYB06OsfP/xXhA+bt/UnQSgwHPDqhmnmKV71A
aCRPw1gwUalNuU8tFaSKsOa+QPOxD5Kwn5efzhPg97qVzBlo4R0dLzI6po3+d3uV
fO9UG3GCkhosTz23bKtgosX/O7O2PDYpzUu0SWARYHwyjZCJINqXUbZbGocpHOXW
gMMfXCeeOfcClnbk50uuK8DOB3hxnadteLrfgO2Pw1mY/lH4avhmZJIGy4crqKLj
nu+4ac0y5dgKEJ51X/T7ceim7HASSuWpXpgyyRgPDmIIn7TA5SSn/66EbpIsu8Q3
+amlc1MX70auFlMD9aL4O+n1evj2AvWIuR7woLlVQEUbgZE7ZUJp3IOYyO6g7Ah4
LKLBxpOwBnw1S3/9b4FOL0FE29QRbubabp5RUL5slp7sJizplZHdYTR7FPT8tAwL
xRaY0SdmMkZ0oARxh5I+RYQvSmCWEZnPsnxJ1TtdTzoQOWGTzbTcZcuBudBd8mx6
bCR5c/OW+d6VlZqS9I4hBAYhzJeTVtXIm1xF4fV+V12CBvK+qbd/dSH6Z+HNLGDV
f6xQxXyR0fgZflL+zdHrV7jDvjCoKkPqfAoBXtzeiIwkZeYP8Zw+862L1RYiIiFC
RT5ib0CeotBK05OwQo5TPV1EFUZ+b5sIqbZgmhOSeBIP869vU2TbqwBt1T6wfgNq
4x4hT0j8NXJktKVJm6W61ezFJNsqhMwatAM+NneWLfn9HFYUm6mP/6+jikEq9SIu
2AcivsyYrpn4UWRmcrqDnlksgGVi/CYQbNUtJUI+GlOIAaSkZSSQqMaZ4gRdtWFm
RvNrVWeu0qCzrzFK8IntGOzcIbphgPIgSaiZASW6XA4K1EAW/9/GALSomXBWYgqY
qO/brD/Y4xawZWrdxk2eU3DvwVBI0ZhsWMIfuII8v6LSyZX0ziywwejEncJ1X28/
VZlew4eK7aM/Lx0K2vVOdcCeI5EGSt3ForHygCgmfctBZjBChUUpsd9mzyZkljt7
N/wyNBSNnTO9CvFZp42QwUqdQkCAOY77hFdFNjIxzMVGzV43Rjzfp3P+/cGTHvbm
0AXJfduKL/ZGZkNJ0AvzSPwX4uAOTzqbyebap1KqHXwzPTRfrh8Sq5tenIFLDjpc
8pNmILayDqTIJomcNRmigBBVaannG44GL+lfVF1ABjVM1/10KMIXPQGy/J5qxK5B
JH+XtNBTin8UL7iikjOVLsIP0p5UVWkKZyEGuRYsCou74/dMkNFV9q0HW+aZJ5gq
MFiLVNh2PWf66KoM74ypoj459ZFb0OKv8yxSY7Dg8AI4Kc4VfXsL9dQs7a3VIq84
flShnGKaozZ8ld6PziICJNLCHgi/IY9tqpcUxoZbs/fVgD2q/ojeyjIm694cLsSk
5NJiJGS6HsLR0/tepq2+5JabmOtTxDd5KilgSLq+qzXdqYpfQ+x+fsooMi7y4sfQ
wwE/0ybzw5MFTe1dPwEX+kxFMyZweeawIrE5XKfoz5rdZ6h71BciujAzPP1uqRuh
E9R6ncdBvWKQBMuEKtQyt28jC/OTMfHECO29AIrWgmDoi1RDsc5HAimwixHrNiUg
hXYQCt3aOylvXhEOtL7HiPq0vPo9EIjyncLNxWyniB1jb3cHXdlzbu87YVw/WXlV
gqRBaWUstw7sSkzBf0529wHE3lv7NomwiD88k2iWtGDEkDVL3bbLXs1E6nIASKfR
uJl8VleHabOK7ziwirH4hsavntkLJGffIOBZWPoLGfTwJ5von+g7TRpgDOfoBQ8E
xFpSRC8Rc0+Su6nSBXmgRIQZTX/zVFeSxU4cEesVEFLdNlsDJLmOb/A+ufG6P8d4
vtIuYtvGG7AnfCUl7hs5bHkxOVLl1PCW79uEdqxnUT6t1Bs0sYfmGF9VASdfSYQ3
x1vT/a3FGzXU0hGkHSJTODaniYwxZnRid7GDpj5Zw6utt9iKVYaaB3HF5c9sfzQo
NUjGFjuz+aLaw/HKBLB4/WEgCU8kzzqWyCz++x50wVOukv28mLmNNSw0Bs/5/nYD
3oVleM/tIBrjW3Pd7JNNwKScQbUWv78Tx5p04Y6PAMbcbmCmiA+wAha0GnuCALOK
8G2k2AObVsFl1dQfZRM6AtddhSSs/3YkSfHfqTZDIA06N0KyCIcUxMUVtDdW8vkz
mpxaUR6OtigUOCcUUXXot1SAn/exqegdMEt3GpI+67yaEoy3mruQbJ9Iggoe0JWT
88wk9mlMtxJUgFuZPMSp+3lL1pT6bBQWQnGIXfP/XN5xj7cJDbA7C8Biu3M+jwir
74hYP6K31JuP/yb9xYxeB4kBwpIh5yuPBdYEotMrZwMsBpFcohasAOqnQMzIQHQi
eXniFKoxeRSIEaRQ29eprVhpnc/ejcB2Gm++fP+860yIYXb+3pA49tuN+mgnCLPf
DQpHtMeKvmkV6BMi3GsNaGtZ2tM6AiR2WbWZ3B4Htaw9ahwkuq/tYq/UvE9eKvKu
w9unjJs880wqoSWpVBt8WGuH6g2hTibbdseSYS5xKEqTlsUkq35RfVFGM9qfyFWd
vGaeetPk8PYv8VjetmvVQpReDtdMDjqqjR9BAoNIizKfyReQmIUnoJsU3RMePujl
B7RITJ6Ih5p00f6QzUrrn3oLHsbfAcb13HxQmmbFd44FKGkVfTOCghFPFNbU9scR
HzlSVCoAgwPbyjGG/QoZNFg++xb27YA51K4rBHpGEr8Qsn2SQHkE13JYlk9FXEHs
vWIhVKj+QX4HfWQZfzmvOykWcrtG+xdfgsAKD0eZVK+9PB5TlGq0wZNHjSSIwCEZ
KAv4MEoIStkqPfwEKDTsG1jXoZLAeFOrAUwGCHLjGmC54DpUg3uHTU4kyaFa8c9Q
Oz19orKDtrTUFsfi8YFwK+OtAPflXgb7oKbuouC+qqFH7h86qPCsuV++nyLjJ4T0
XiasBiu7ns948dWNOue6q+iLgBuYLbRyvSnKICOcWHgn49v1RlEL8UhMKlnXFOia
N/KDyYfigi60rQAARe96LTHPVd+tIk8gZjl1Y4xrrrITgqlQ4KwQd1vlgSM9Dsug
zRHWZojHgPiqYRGmSqdwkyGG557ejPKHNYufzQM9RttuonFMfJcxDceZb5PGPxHg
wm4kKLTyF2NAZZbq9ePJLqQaYg5L4mMe+W4c9mniZ//5z3PQEktjsZyoDrFtaCit
VS7G+R47KvMUbFp2LB0fevj3B03gvaV4pWCnDGvvts5ZEe2Sj5+8XqRU7F1k0/lz
zW71llHsx4c6ddiggud2otldNucJ/bR4wvjR5GnVoqfgbgYk6qp2cd/F18hLNTMC
8OI1hGwGMWUTkB/+BunORkOjZdL2/RdoyuU00Zpk65+i9dL/VKtzFLxm8n8DrsvA
TrYT42ViuZ4dRH92JFW1XKf1t8WC6tkjbQJLC22luc9sEgGeHBZ+iFV9NrM58PR8
QvlydJ5PCLihUynVE4Z2PsvzqLIeYOEsks51ifn5mQ+q9ev76ftXl+DUE02Jwhw9
bMsA5v/zuGc2VTwf8sLP6XT+BThoWGOugOYZZ0/v+Z/uQWZN9lXQez9h0MHFFXy1
XLFPCZvRLYencixiShTh/dJ2e5kl/YMoYlzQpg7iRt0tdaXyj/BdPhaDQwlDoIRu
voaxtUyBT3n0ntA7VpXgBDcSPgzTgg/LhlYLIIbbqEMQew9qPQVoKAwwe4OfGP3t
szNIiorKj4QI11ePjvakDNF0onQUS7G3NPy7Nlwpnu+QoPts+yr/W/J2RFePTi/k
ZeRYSLj+ODqYlxo2NR0KFzBA5C8oJ2GfJ8yyVFM6HB+hI0k51/6Zt3WQ/mGubdXR
gXk4+f/K2rCY/qygDU+M8znHOQhqZz35pm4y40GZDexLRi2vR6rWUmqVMKZDKZg4
BRramv0oDb4pVtlvDAirmaqHArpSjGEjWy9WZEzxH2o1iS6cx0Y4Dmc6dwxr+SYA
pyUWcOfARBt7XeTsxNboKJgDBE7sNrWn1PtsHZKrIV7obNuakBl2duPiweZiEfXG
U/iC1ygsJ9Zg7HwQu6T067NjUDIjWic+nplfiWIMzcdDxc8EMi3w1zjj6QVhAdAJ
neN4HOl4doH6pzx+I0ITI/dJ/dzLl44GN1y4I4fCOk2bC84DP47TkoLTK4x2Cj02
7AjvsyFsZdc2IOfmMB/ziicLeaw0fbnz1LYmQJjsMbxLI2ckjVZAa1VW6VHnBmlw
ZJh79f8hb2f7jh8rds8l9jqSP9v49ZdU9SE0AcHfQG7wBgAyMf+8q/j9n1IVhbrx
3tvfqF62GhABt/qf8S7uH/D/lWk5oNqtoFyn0GOYARXcp+0OqbX3T/cHExw+LOQb
10EbcZbWpoFaUGcfGicVP3OvOaSA0DuAOwhV6Au1UUddGSesYBdoSciVtxAWcDKd
pp5pyIrSBePraSRs67c6vT3bpoSSw7Q2nrfqOpydI2jViMbhiZwdyBRsU3kmBmB1
/elVU1nn4i9wa5/FOthVg3b46JQv0wQjAoSd61npK/WeEjg7CnLYD8O0FCsydo4u
+75iW97mbZ7OYsK/IUOr+piBVDSplReRqzHPRUFHWtAxCrzH8wNGPcUwavDGy2ts
lRzRfaF/anJVC2azFvWaqrZaatBPW17Bpzn77u9OozcecODszxDa6EU06sIIoten
f6qsTmxNSAkyn/hIAAIK0zN/TQFMqrPP8j29DpaX/uvJocNjRSQSfTWl7J1qwr/8
cVfnCg2gl2pivKvp6lABCu3Xaj6V5/bIh4gGJ88MEWLDNwgkDGhW4vrm/v8bG/O3
pLUaclhSqueD6GcbL+Tq6nNkhwWwEcUan7NKPCnmkm5cbTjRhXE538r983LaCt4l
M8yr/9cVpeLCoc+EP2nnXiOqhv+YcfFn5ACB9N2pyT1qG4TQB+F4oAFzn3dN7FIV
35EgaiD/4xf5gsWLmch7Ci3pvJVkFLHxvMuh9E1i12yd7uK36qXRO2U3RtIG5/3t
t9vKehyMnGappTW3vsDRni1c+K+2TQ/LzPo6bwVdByrLNGkLbIK1F1EKXTBShBi8
xRv0nwCThLMICaAIsyzNZq/FkXCwi1BdZWqA/wYEgyds6pXLyLwCORYce/VPa+9z
/at3oNp+MYjSYS4w7DdQ/at89BfETwlXlwn3Bc/0KflESwfzxjOM5WvKjDgyafYG
hX2LNGmh/Xsxgo1Nlr6BZZw/lX8Y4uA+JCA3e6/A7AeLJxuXoHQNRSYp7u4g75Yc
c5R5ihQzhCFk7SciagAeHaYwbOC9gW8DGB4KR/PVWOhR38hDAgN6S/JXqoBwOArj
vfFZY3ke4V4DPkg+h1uJkx530dtSmFH8TJ9/3iCad1KjWl8Kz78catRfe/jHu3ou
VKjeFVHAPAyFwhMn+LYOj203ai9X08axHTytTgobSSLDz27/SbZOHdiQG8JOGUpM
kyLb17jtC4L/nDWwrOSCjMbPMKCsniXjTl3U1HBGxjgkutkClawvE/YxUz+e+lZw
QqdKirOwZ46ZHAkYZehO2LZVvQkb/qO9pPvx4yuNYoPpqH6LhM20qoBe1M3/f1TV
pQsaABcfkg2G8CSBxhdAAoFHiZLUe1w6dQ8ZmW61gAq/rIlBw5mpQRFWE+uyDs+9
36bn6LdOdVEiti0lh6miy13iClc9utnl/HPFfOztJkyvhh7+qPNefzhMYzYrp9pU
1icLOR2GWrQ09FORTBottK2yeEgE5O/51coUXZyo00PyUUdK/qni71X3KN68Lil/
+wIpMNxi+DyR2/6ja2F4p3H0uYWAXZFfs3P6PlF8ZPSlJrzYTgK4Dx/UNgjyCjgh
cDSmZxSQqsMDC40194ayzvVpeGaUXW1svC26Uv+/Wo5RrwSSnmBcWKCvw0ptU1rM
twAovR0mqft/HhGWq9qwmOCJerNsiuooOYl9YxxI5kSOg/H7W3o/gadEZR8kFtUe
h2JtYpcUnC9jgK9kzkERvoV7WnMtK5uM0WOpb1zKwhwng7KKDFXOA+cIfa5lRWqX
E0+zuyTZdFN1u5NPPeoHNPuUQZJidx/t2FYTU+cVbByTKcewptQiRAIeE26gl73P
4du/BcrQFM4sLIkCvWRDtI+bQH4SiLTNE17+8YpfEKXOkbfHM/sYZQMldYqq23dX
ND6nwNJ7ZPAyhqWqjiwvJLZSxdJuINMPn6n9bsSmpT776L1Zw9NSZ5gYaUIcN0Mv
kD774gCSin0suIMr8p7M0qBZN1PahgBviJ8lEh7ijhDoUKpP4qUNMrXd3EdgIOuS
kVgNOpgBGGGVCLkIaA0mOvQbBF8i0OWxDrhFA9jNLqdb/gmvs3j4GqS8yS55ql2d
ugUcM+SDX6MhCAsUKYPrHCi4aUhfJK/K//J7zprreK3b3m21SVlDoDv63aqO6y0k
GBLDqr2FVPO3PA1kP6Lw085pOVYQ4ukP+a9wp7CURjZT+mV5sTLo3hA7sB05IEqc
gRVcQd5tGrnqdDBJadhOJG8VjJ4DQCW38+GMQF2GB/V2GNZxoSLILpjb93ww7wS5
JT+TH+L+NZyuQwolKU2HKaq/l+c0ZgIPLpWa85sa07Hq8Of+TyayVOhyabevSBH8
kizj1ARQWhhYF6o5DaLUu4aYxcCZAjedkEWV/Tc7SADO8is6D9i91Y6XIreS5ksL
IQrki78cXoThVq46MqVWSwZUX83CEvVgpvIq+aTei85GH6uXv90p2pSfnYVgwJO1
fZukJOS2uOMreRsdnHQlmfhPXU9rdE6Va7Ph8Mr+L1RTnuz7M0TyMim26lzU9LRa
8xKR8al7pDMWM1kFqEDzElaUATMQ6F0Qwh3uioVf6zTdr3MSssqlTo71z428EnjT
Zfx4SqHIbred96Yy/cZdhqmwKgXE2kQF8RgGGbSzUWlMLOaPDEQ+aKCuY1yOrkEQ
hWnJ9A7ZyzY7inM2fe5Qw2xMEKaYWDlXEVjIdryyDEriB/4K8fg3c+D4SMhShzh+
vbtl2i/iQEXhoq5q0QKj3oBdmtU97WMbuMBDVJbECMRkCR8yHl8zXLTu88nl8Crp
nE/PKJ8A1CLqtzLgh9kNzFD6e2rUXo5/OFYt5z7zDwmtYjQ4qdy9nAru2S/+BDNi
x+yEQsp6OVvK8vrfmujlIug9Y/4tir9yuqFgILGxd2XvvVUKxGPyQhL/iXIQFcz8
b3L/v4njVYIpg/BuVm5eHfZMJBdpzkX1+HoZjyQ+YZYL0x6MUMG4JRyL3KHIEQNj
0msqPhJEjyCCBOSOqWB4KmmRBCbofRMKVOifZPU2JvAHBCBzdgDielS4WhXO11Vv
wg5VOqna+n6M5AwwA6Cy5Ll/z4PxlI7o52PjY+ZdEBuwMXolj+nRNWrOCymvrSnn
TsCG4qXpEa/kKFC5tWeshr7vn4hHYaoxlYJKWU7IT8XAJq/UEbX+z4M2MWsWh4u3
2CqMh40IuxFutPbD2agPvqi5rwVhl2IwxkEcwM7jRmPx6eGKRqLgSgQsoNAi1DPq
sUGvsNmG0vZuP9A/7lrtdIdhJDeKZeSYtB4KtKioqa01YuTzqKTjoxs8TYY5c29X
d7pvV2Ee8uyte1o1LdvYPkwP+TC/uaPbPWbl+80Wyzfd3yq0I8uCAmPZeBmAdJbC
ZxUQACntGYwdbi5qeFcFlONXiA2AsccC8XnysXvR7lUQO3cpl97UOOklHclfvW0A
I3BCpYK4BxV10WmFGBzdbb/JrIaSdZmvsdgo6cZY490I3XSy1yYE6mF2xJtCWSF7
WH5DK7ZaxpHF4JRd/x7xXc/pkVdAapGjhKQTLPWGjOwlSVNLSUn9q69xUcoQ+032
3EuwKeKjkGM031z6ahSpO0jk4U0ckB5HyPsTHRiiFUb17nxqjWZBHxasH/yFheEZ
d9iOLgIVpCQhBeMyEuEVoADDQ9Yi0rtVGlazBx2mxgmb0XM0GhUgtvah42Tl85dZ
M+lYVf1/x8EYqwoqg2gpC0/MfMJBzR9DL2yVVgE+HQxPy/Wl1mu9SY9O/aUfJUS5
hWqFfmZIyTCNl/wQ8ttjvdSVZC7vUHpZesDrvq3dTWIp3F312sqQUXFuI1N539sn
b7JEUMOfhi2HlarfeJQQT3IoDIvSBpUX09VwaJKyk5ECcQh2Zx+JLcttH+2epz6G
akNcD+l144I6qyTCiCjL7l3uB3tibZK7LgNhUmHROfOjRZnMaYolIWFbIfSL5hiG
UvcUNnJZayokGqeMHLqc/gRUZ+1N8uve/URC65gT+M8N4UgZ1MfoXD87wMBTLd1/
UPJhwHJvSCbcSm4WiNHq9OYETQDTBXRRAl3QiXix51yaa3OPOJR7SdziKddYb0Kf
T/qD+UlgP3zIHkL1SDnj50ir0Ic4Ha5uH9NtehNQnucIG4jQB4skaUUHO9JePxfe
etyplDtSY4Y1gE5dkW+E/NN7T7atcRRumr7t1DBVVjHXsi+4w84gkE7acDym/2Eq
HLsJPUJAnAkdY0bKimNqATbeDAipR7oEdWl1wJzh5xFGpxlQylaibLxQ8kDvertn
Aa8toXsPqNYWoBTD0gWe6QIA+nrVcOVxSDGm6QMeYokHZrq2hBaX/D0uMPahQt2f
7Ce7nkdUidyEw/CqLF1rEkPTp+ZJXLTxKQD+WsQCUFq8WNKYAJDAb9efBAKdkKel
CdH5mn01Gyu9G8zL2mi98toWaNeSLk50B1Jcn+3/CT6SXw8X6xhfAphwJQS8xyZz
PD8LqvwjgGi7ts4XpR4GDS67017nkAHnLUSVLMOraYE79HgMOF4JNALI/5MCRsch
qwEOt59fu3gbjdJpb16PhbrDRDsHgacsvTXex7n4Pzb4sAtOcrOnbwfmpsuRm328
43hsbipp2g3fuRh9bmEjxhV+C5f8lXwPsxy0s1gDxGNzxJZrXBwMGNFk2/fsu9IB
8he1mG/aJ6errbWgyZ4CQm/JeEtfr74T8cLelJmV+VtDkFrZCg9HlZYSXH2BmAbb
3mqzpaB2eBTPLiNnuSLjnimXnTOWvWHVMAKFy+ayEMF+HBKGtim+Ddd08gvx3ewN
Oq4eev+2632d4v0ozp4PQtY30p0YDDR6E0iyR/UNgIk8cmUbe4U6+asCXdvfcw2e
NGA+Fqu7xq1JwxfGMmLxorEROJk9WB32znpjeyj/M/GRbzrNsO551oJo1M5lEhlx
UwALDoiL3TBzktik40c1G8ZWUs4jK+nflcek5UneA4x82RkAE2T2d/fMPpXpuDwp
gKjkZ6m3DW3cI48JrxEmWXGg9tyVIzC1d2R8QzwWN0fWNumBfK7cXnw3Szz7KVpT
FHKLPbr9tDaR7r57EPTQ5N9ULL+37ttDzYZSwrd1Q1XmEX0gAN7Ak31rgYLwC4RW
QGIpnwvYw0aKVrX59/x87NUCgLn9CxhpcjrTRXKHPGTlGUMU4HgCgNRpdzF9ysEt
94+M3ocMuefLh/ePnTIqw19yGdsZy567vOYiu6HHG1YSV03qHZc0FkxSFnHc7jr7
IASvG6CjXKIEKcxXMsJnJaa/goyB7kQ1s1YdBbWkm96ChaHIFksB980lY3KGr8lv
TKoBhifC99E/Rf6R333oZHtk7trZF9sTF54aNWs3EugpHG1QpftcbPNOmaZhzjJw
/UFtbIKiwZ9oMw8bfeGIWLMWNHuswmciEvyW3QrhIEE7SRDWhnqGkKdoSOMjPKlT
5h2ZQidEEEZHDtGUoIVu8hstx2+nPWu/Ocmm22NnRaGnwMeks72DccVX+Y4hunwW
2tcNa3ULjHK59pQDnbtm9YCWRSUrYFVGBXaIlcxsLjc0DM0cOgmG0m9aHoZx0O5A
vIK+2D5fiS/bvA5Vxq9QzLlua+fyYbpaML6J5Hk4Yks5XdBFSixuWKnllK35gwRX
aDaXKkMSZmmV/Vovi0BhgxNCdGKlqvvSiEjLTSpriJ1fBWI+/UBXeKpnKhsZOOKz
ObCaKASq1UYpJV2SReiV00I9YTaf6AYPIYWkFTZ1krrJDGdDKwY7j2gY4WW36Zyb
kI4OK3DujkqyRgADv5kyX9s/Wvj2mXPLYvZYgT3SxEZsawAP1KWD9w8FbkMuOzt+
Z9DbI38tnbXH4r1UpjhAKiknW/JXXzTW7dC28pP96J5mJai7WPq2I7VIbL57w8yw
RWdk/gDEJVgeDOE6Wl7UZHSvwuxeyPYerBVD+2AReCTV6/YSczI72KsCrc70Gl7M
7fi+IOLQ4NH7JpiAnsYNKcwXwd+J/tPZ+2nFiW85c4ZlEobnS5gjCwE6zwHkXBG0
Vd0AKv3sWkIqf5jidZzPa+TeTer2h7P8afwXlTQaSNwpyEzvk5e7xOlchUimsbLH
62ZwWluoFV0ZtK50IN4YsizGbLxwiZ0fnA4xMFe6+VHXqM79zVgRmwmY8EqCyNMn
LDuSm3ofdcEKVrse6vETgxdCVGR5QKim/NE8KDGPD7vdbWyQxPAB3Blm7XlqcOMS
Nhj9zIX+BYj++y7jEFKw1E1S4MX6ksyVrX0Pj3O3WSuwJfVwiYVwjwK9vXLRSbt1
ISaLYkH3v1v+LhJmZJuAPlljdgf1Do8kbsQzRM41nCPq6girsO2DKQQTihRuLC3J
/ZSXRcUGM3BLarK0gHLi5tyRk02+JAhic0hDwk+qGJHmvP9bw2q5ShA/R18yv/4/
wCJJ2M4adS7adW2a5zewAmBc++bJqc2uCU9mC4VWlVr6vBrDRIyPLu/j7U1WFjJG
W/4fD8vlggTxZ26kp9XcZavE7RK0JClKad4B9AE73C0AwVy20FdQqs3k+tmbUFSr
JXgASW+0aBRaPdttL24R1bdyQYvRH1omAWSQ5dM+Yf6wRw7f2+bsDSHE1GacN8LL
cgwrQCQv/a53XK3OAaLMVKvFOnedAgcsBoQT7vaB/SuKUPR60Stxgyb6RAWixP+3
SVw27SLBUfRPmD+YoIly/w3I3eiVrJo8wIR7Fesl0eJ6hAKpb/T1cAYuTGLKCaVe
QL0yFPN/avEgpEGmODNQNMOT0wxC1+02oHrecPBv/vbvo0rFAip3AiNu79gYDLEM
nODNgzZE2VodFtYolbh83gZdl+ATZXjNfSbGIScQ20V2TyrLdjTFr6yOX5UWSy9E
kQZa231AMA1mIfbwsw6iywc7yNs53FPzk2uBcSaTEcPk+CYvw3l7GlQqWZ45anz+
MFU4dVK7Lqc3IP/gt0m38k8r3mpAIUUNUruFnUSaziGpM7KjAidCq2wrJPHTOcWO
r0ahWICHGyjl1y5W6X+qXNLbJjW97mIhRIfBwLZRKl04TfKRtqSGzUesKw1Xa9U2
cx5jxeviEvZrwiyqoLAQh1E6LImHInrxocrTiP5+ZSAn58netMzpwdIJUEkGFnVW
xV7B19s1xMZ3YhH9ecsIJtyV+LY7l0f15LQAS6D3XKZT3vY+IIvz/t3PM0ZNqoOP
nGHdIyLL7QTt1iKQI8r07qawGY+/daKIR4VcFPV0v4PSITtwZVOnHPOuiQmAKtZl
yP8xFChQjTicE1VcOcI12+DoBXyH1GFb0vScFolvEtbSTKTuvk3jQhataIdrERrN
lRG3txe3slfzzW9VvanQSsOghc30NLGseJUxjcUmc+Q33BylFdxltN8iP78vYZA9
5LlYAMIJfBoIExPnAYH3O44rHzyiTvFCTRVteDYXBZ1G6eZtTAB7bvXfiH8ZamNS
3AhQi+VFShjtNGcPu22TMgtWK9n2uYF4Ev9XHVabycfMB03QrGNAQD5O4TQKxavU
0jAVPxrvdAt25+CZ+FOWRpLqwpi09xguloV6n0xJYDT+OxfjhOAhhwX2I8a7/MgL
zZcS40x8U5kPhbfhizvF1r7McXWJdcCaqteIkSj0rF0YpCZ2FwD01Ajb+HvyGO0g
sEH/p1pBIDiUYnbq8ue+escIZoGcWJsjabtLu4B0DHde0bi/pkG22LiuLSi8lBt2
g3ooxYWWK6og9MUfoZBiztN/I+FMNVK5tMxVPnDEzQeDSs5CQIyBO8Hixj6wSRFQ
DiZ3PPj6lchwfcMrxM3c3+1aSDpf3+8C6zC/I97a9gMuz3qs9ZkOhiHwU0IOZzlb
OR53XlrJjHgUwf6hMCYgJ9VP/shVloz1nRYDyGB/50g84TexvgqH76dkrRfiVc+E
Aysh024OcQBTj20VGydsBs/MJN/Y9qJXMa/GkroCRBl0qM0EX5L535gZRqhPQdhV
PMybzcJfpXgIGeEjwKlJqEfUQX/zENL8hqH4OinKUZMUZX2mE28T6w94JiiecJ/B
EVmwm+PzjC7JdXiTFV9oi6e29SLTqHupvxQu0Il7Ib4gD1FB/zNzDazPygPefVJK
3/jils0YNgMSRWMXIAy9d5bV+vh+isUHLQeBLJmSmsY4jJhnkd9gjC27XzSJGz9r
+l2KJf5Ozi+ak1NBhBv4RgVmxD4VsqoyHfy9GW9i39tQr6rIbCZh9BPMwUAJba9s
2D3zKuYn9Mth/KXk65PLcC8SYBcjjX/l4FQtVbsvPxY/UTHIsRF3QqWV+mVwk8x8
AoXV1fC37ivXtMSH7ZgZpL3oizkwoz2/TOj8zaTyzvbAVda9p5+TIvho/uQ2/LhG
dxP9ol7C1YczEwKdQ4O2rS3f6Kgwiush37zT2Ie3g2soK+qs570fTQSLZUuWZ8Fr
gTcI37yGtbAtm13pboIvaXhxt6xZwEcVAmvuO2/3IRjiZejLglb2qLxIb/UaLuVN
j1yxpkhxJh8MaD6H/61vVXSjPoxuWUMcsnsD6rwaFMD2vDYok4Sxn9ddjZhyBqep
iqR9phagApzuiVbUlRehLlyRRD7pzmtfqZBqwhYVIJEph1P1/JReTvjs/qxc29AR
wKX2gwvSsxm4ZHYdNEY8y8gskbndBloqpQZy6ZNnDvLh6G8esl7P9cn2xRoLz4So
Z4Qh39EXMgcicr4lr+lMDmSZk/5khsZg4vjfbcbfM2+AND97d4BaD5g3y2iSQsv6
gNWhvYk3vYVaQNfifxbLLMtyDki/C+OJZ9xXRExTDjClLM+o6flSRv0ywy0bKSAk
XlhTD0doAaIBJ7vHbwoFt1P3YVgxA+oUl5DefJW3PGIXd4q710iKNFaAByZzIKvI
1dsqrE7TK+Pw8APWpIvgagTC4Uoj98bEVcuGlI2siZ4xPGM8vYoO0NeDZry3Cs5e
U7j+jzGPJzUUhSQ60TLPjVK9pGTUPEcdKCHU3PhE5HAQcBi/YCw50TNnM0k9pq4F
I01ofW5z5WQEdf2e4jP+lNdM4ohKUAEY5kQlGEeF2LWQhGBDiysHFlFV5XHX0JXD
w37QS5qsmSVlnB7ZmTd7EK1DbrGwT1Qv4Dyl2wJ999+2eiBGz58thj72FVSxEGsv
p0D2lARHYsZbg8HJ/2V5wGQo+AM+WxXI4Xc2GFYV5TVfdcC0MdvOTeuncL4SOWX+
6ceZWVWe4sY6bk2ggqryHwlxCYmT7TxG6x1ZrZ8Ud1GXCiuyjJmOP3gY7Das9h/p
NJacEJgfz6nS1BAMijit1rWZkGlEJP9EA1ms/KEkb6iFHHDxoY0Id5T6dl12y7tY
VmeFbStjLOGN0r42zRTFfZX/1Vz50AUySo5KZotbw6KHy6os6q0oSXCnUxGPNAUH
HE52PU344ohO+EstrIvvQkeM7/OPYci6kqiKWWn+Lyt7u9GdXdvJowyBv7j/XmqQ
dJ9qjUXhY6mSa0jE9OGkOPM89Xv+tBmc4LB/PibCv5zkEjt/bSAjrY/r9ut68e/t
LKVpzg8Cj49YKA2Q5CUj6PmiAXWGqrEz78I5uctjn8DzaZKAY3CPdktoNzCrHEOZ
Kpsjd5r2k28yi3043PJAQB+XqagxLS5Aytuh3+aF/Ct1l6mbQ+i9xVaOzRxHR0Qr
RL/ieQaydheb7/W52+5ecGy5RPaocBHSgQV0cZ++I8H45vKilfVkLDfk2eygpDdY
KLVuy8+fNE0K1MGBVNWMFBeQM1nAGBkCyAWX7+djuqH/SYvpi7b4SYahtwJrGfYp
ZL4BB8Q7X7rFDauISD6OH35BaNAVJgTxkH8FUxS64yOJ19mjlekpSq4nsfOlevHX
OA6Ps185Kwj5/E3q2ZIoYFe0s+DgYuodj+/sQNA6SUKq/blP+p0PGTWj4xIayZOm
zP+TcbfUlMYCVvSdX9DG5F/rG82npQOSQGLZwiVT2FtX7LPCGl2ONCos9g+AMY/y
ufad60aIv58EXDT34sqpYru2R/KxJYkCwQYT7iSy1YP4RBGTtj7o3tmKojKYVxt1
E6vct6t3HZvb8Jdh+NBmSSUUZxb/DQhW4uHikpSO7oaiMAL/JHQh4UGFcze46D4l
jLSSRpSS/1tt4LPXnDRNbzPsugYwDRLZtJqwoJ0+7qkdizvsRtmNajbU7QQAFaqm
goq3j77AVBps3klT+aFXHCe+tdNjvFojpR2dQ6GteRV5h7ij18zsfDV+qc7NVcYC
mFyQqZyFohOg/zZeLq6Zie9f9JPnKbBqGnsWkQ0fsvRRheuuhDKt5zA2pFyjfMTB
sranPEG/80yv3UXvlzKx6RYBivwZUH2zho/q3kYU65+fPGloIAukzjWpujZ2twGD
ajP1A4ZZZRRvDRVl5PZPSPkaU8vVX0L5ypzNGPE/CuEbVfpNEMgLmuogCJBUjnN9
D/e5yc83Q6XdugNl9aWKYtv3FTz1wPTBdtzYzub6EbGVXkgryiU5sf68kabsk8nC
OLh88LzmHgcGCQBXT4VLSfqaq28XmZUzoR1cUqRSYZpT+xqpF6Ci5Pr5v0ch9vB+
9T3m1RuQ/XRDCFFdV0xgHCKPtvxxjdAfcdau4Q+HyG5CIHXuzTreKpgGV/foQxXS
J7IUVBrTR4akW6ZY3sW6rvDj/q386ekuZUo0KecfF3r//AJGOAxz6iWsIPbRVfWv
dKKCgyxnFImTHeJW5q2t0HY0i9JPt2Me9MnkSoK+nVXBoUVViPSNR42peYMwDBAo
yV4m+gaa2sS6TAwHULKlLenmd2RjKjHHGZYYoXME7ElidKs2Ql8jogL7qUOgVGcD
I8edcHk3hQFaya+1tPovx/uur5J/u4hS3Ig/9LF7OrA6DxZhQ8UxAbAdsSwnKeOD
sP5GxdFEUHXFI9fQFho664iYvOFbW3bbgV6Jk6Q4mwmyD3k8NvwJUJf64EYoE85k
f1IZOsxisU6KlLHyd1nZE8keywoQfXAaQdmxa3kY/SXtjAS+O1Z6HteKJ+Lc9khF
jc/SKT93WCGtHMFdwWJlL9enQGh207V7qo6LIRARvw1MYg4qQ+nnl7JfK37T0b5j
iU4gb167HAqJ9hiXzCk0Dx7oQNt6k9WJ+RyyKDNMOHAnYXvf4XyYyQ71cIDd26WL
ah40wifp/4Q92CdmhwWLCZUaTi2GAuPk4PhrzNnN7/tNxQwmVUuJSVtdzA6aJJ/1
/iMswwncqnuT9TCBONRk4hGDM1SFAhA+wQ7GVNjwMsxbHfmn90JiOULJk7mYFI/S
Tq/LjmCrftKCbJSMu6T0BSk/lWN3uxMiscLC/O0hSn+n/P2r4kSHLYdEEm+tktHr
R8QVNGnejxZMlEio3rXalU497nUoZtRGivPlVfuErz2rRukvDsH84qSXeyVyfbt2
I7PfDg6a3P4NjD9690AUX74I/QuYvPLm2AAkqKFFvSk2n+x1MSZv/vrHyhGXWtyi
RQ4kb+ndLAf72THf7ne+b0eteeWCq8tvMXsgY5dF7VC5CBmm36/99Y1F0jaL7pQQ
aiHi46hXAeHtRVDlZqX4YxEv3b/aICX1M7gkCNFoArW1u7xorb9yYLCbzD3cctgJ
ApNdh1qHCW8MCEP136TrZFHiDQUXvOfMelanQErHD7b8P+DHpLVjcHulBBpSJClO
IN+7d1z7A/cE+n9uKFVA0tO/R1cwJV340HJNOipqqnTBK9JQKOE802CAB/KCLqKX
VpsnUOCFZczGLtuCwPzxYieUUCYCpiwJWuhElS5tssd/vuKRUaYPKtvwPS3Kr5PA
DB2TWrVTjOXJkmfKzzxGfKYvAA+GMLtNasRm2SykAiCk7FJ0eM1sZd6aFZRBwFFB
d8ZicYjUTzhm+XBuTnvLD6HvkMXudKrpzM0bpf7wPOSRXjtwLAvzD2erMGmdfJjN
HgF3OxxtERbrBNK8w9LSGp9vmX5XkJWOCbqVRR9VikQIvIBIKQJj0cqIGSUI5jU3
o3sYEyRIaZs8jsw4HeEkLg1djbpyXJ3r/9ZympihvzztGcStE/sioLKqvj7/HII9
sWJc39RcBCEMQlw4zc9f9NBc3R5ytj78S+HgxbodxX5VdOn0qxE1J5jntAPyKekN
+azC25QbmRmF2OBrdVSwNYiyKvU4YmO0RhRhGJIgUE9V72qsjmXmHUgyx+p2hZMb
Sokvg1+oj8P0LhmvdBNYjTTq4wIhAkWcqOd3PnHbhyo6gpj7OoocNyC5gWQpJ/F9
onqnhz4x1xXV51Nh4OGw5CuMoaYsar43msWhqDo3ofGv9KdSukFyc+npqWZw910/
MNcVZgvHm6sOOoz9PehmvuLfmNd3vC7Qd3Sd7Ioe+nsQP4a49ddEKQf++Uo/MpT7
Rfit33xbYUqCcMBU/TbUCtzSgmfbGJgWATj2zYeJcLTa6svuBicAL7EubYqH/J7n
SXeBcjzsNfgXa19ZJ/hdLQR7/WuCIIoyRE93119oAvgz3qFXt7i+2EBY1WH8ipS/
v18z5V1DZrnZ6O/5/iFGqOPmE+hBjntDFgLLBeroIfE6v1tPeTMdqHDgSNRHbZ0F
fCrp+jHMT/tXy8PjTvwqk/6iZ6NtMRymVz7MkK+GKAmmCe5hBO52Off0vJhDuym7
SakjBouuUaN3fsPiBg57xCOePfnHLBiYYOHcCafa/we5uFPLajTuTO9F/1+YiXmq
5tars4Qwjp99xhXiXVbyu232vcKXidoEwmVj6u3U876BwVdy2MKveQzIYrx9NIJO
6ZSCCd0sSAb9FoaFYVgvJO8Y7zFUUGk9Hwr0zwoa0PN8xkNzdrm/ZiwLLNHaCt8u
bG4oDkS92qMYDDIWq+2KH9IINt/UUkuSYvBnizhYOP/oO5WksftyLvN61U9WWmNp
2MvWL7Ls/bckPrCuuqvRlZDHFBkMsX9D3S9A1rTG0XBLlJJ4uWSoaqHYcshbJcjv
aVKkrnY3Llpo0C14tpSGRpivy2ughA8dFs0jQ6SkxYvoed2iONZ/H2KVehbx7Rbb
zpb27PnBM/S/II4Z3uz7+WhqOeux1OVBUj/s+dW89xD07m7CsdpsxsrNVuvWLGr4
qNdeyNXzK84/IdiUDvt9l/U0AtYCdyTtfdRGEpkNed2gRWlumrQ0uNeelYT1KDSW
udY8KDSS3wTXACSHCQQL317N7/y75cx7jF+ZFeWUDZmQml6L7t9Q6DkfRqkdlaMs
IPnyNrO/S/mdWA53foUb3413LXh4ruhHpRurC/xISLI41UvNyV44GKF8JgYKrFiq
aYFkQ0pdVtCu+gpdgSOSh45xxijP51Zshp9Wi/gEVCJxjsu7iCyE6X4IUzmkyDLD
KxdQYId5xImg7cbxVmHXQuZCpuyLuA5ot95h/L2aKnOxWKUnbBAHy8REDPrGjL+6
QEycrW+JfucOl+58xcuyO1kac9YgX+Mv3Rd0aBci5zpHvWsSSQGQDgve8xpD2PVx
R8RoTpjmDqe8PqAb7GicWwb6vxkfDB0KY5JqBbe+kiuT6+FI4W/Mva2EamWOTx0U
ih/DBI+PaBFh47JCcJbwfYZ5FWvf6Z4sHS1M45o8txovuanac4cylDQchzksxYkj
dhEKLgCNCZwumFSriehoZKeIBgEy1JlqNXv7WuPvb1K78+RjZhD/BLu4tsu7pUAF
qiDpSkm6JVjFp2jzmnDjG2cdcN/lpswG5zMA4TzAQ+bho/UjsR6A3Pm3QxRoGa5m
xAWD730A/vkJTsk5Vikq2q0H/YWMw/6ITsQoHh1A8Bb8thszayyM9J3cJd8HmFSk
vXDZ/KwuB5TA33ZbxOelsYrsOmcp/48aKHcK4AHRu2Cn2kePZxvqq5Bq3UPHGoXB
BIIJDHxRSxdhjG1I5wlkDdNCZYFRAVugLdZrrqPKGIt/DFYzrouss6dAAgSjGUlQ
wD+d/znVV9CkznsNyzHEkERRzrEhlrEGo+IA73CkCL0z6l6PJz/iRdyMUpnP+jtM
ksPasoM4gAaO6CQvWjE1DlLc5svokB4yUew6OtCg1p8+cxn1lK3d9RkCNkI0WFHj
/LZVR7VvHe/sRScqbrpcfvwVOF4apj0yzFkqSO07z0YLxB4afqifbX8CEkR63wHz
tJ2d+50e/uV7rD3h7i4rTfQN3v4mkiBDMs9FHv/AmQnb1YEDESCjbXBJ91SjTKmc
/wSzmlGrMRDqG1hSTeepUJvdfDVBljF4pj+EvFZ8e8DMnk2DPuvBxi3/BrtGQrds
+Um63qElVmziceMWyyZjMVvZg8iA6A0Hue+bB3cdN++mw/IH1z17/+Krg4+TSGiw
ka46K0mPVHXCRIv8gO5UxfkgZDfUXNuTJ1fUvGHxZPnYw4jKvfBONZ3AxJpDYgje
8p7dPSw1tQdBf6/mnA1UMOgNb1FebpmXf67p3LvutS6x0d3j/bQ6kVVKRdD8pmN9
xhEbD9NQc5FG7lu/TqoraJ447NVmMJYJFOKTkht21w6sWbR55oh7mk/m0O0YkijM
HyEqJifdVIh6NpXIB/P7eH9UvEnpO/scG1hLQQkRFHC8VNW5rRBVi2AgyuUrqtUn
/ANDJ+mjxTLRkJfgLdTt+vv0/+xG7J6XShxwOAob9csChZ2I7a5ywWbW2kGkMpDP
MmhhYSnngtbiVKy9VGovNDuYoXAF34Vl6ByoHhw7E9Akde3Yr4sm7s/HW7QboBf8
wlBexz3n9rAvtVOvffU8fRhZbvHeyshFiejkumbB3Gd3+6KIPmLVbwIoZSVyYFsJ
PPMgb/m36v88fy38yGJPBkctwA34d+aHShhoHJrapklZgEVQMcphrfbQkdGu3YQA
7XbEsG13EkmoHI16TXh2Pk51fZ41KM7UjNIJySF1BlACH9ZNtS6cL2qekiZVH47O
L+D/MfyXGd55JUo9fAU1s0NM+Su1+QUxBoEYuPCSDNTbUCvs93TTwPvw/bGePptn
x/vWqI+zCzQnKsWR74LLSaoJPqNLfjfhcOY+Um8e/B7vzhshIfIxLcUMNUj3pJCz
VwB9QCVVpN64zzUn14wLjAsQLO+1CQHsxoI6fx+Kc5oekubxGQoNG0jcYxqpTLVo
yoRj1RVB6VCrGZ8YPySAO/rgZvmJudeYpxLPU8iDthfVNPzUZwQ0cxHe8u+EXLJK
Qi+e/fAResEI3jql2ETrDcBsw/Dd6oIUx9WbIFHE+XCp1evJZD63O8SB6wPw1OnR
npuGCXmma5xDxnq6HS20I2e1lerYapBgHzQDwjZbHmWSHRevD2ifCp5A50nQ9doE
93uAuedXAILpjQoH2W04NpEeOkoLhdAW30bSVlzcXdaSiRB2L8U0VV6XHTUUXkxn
QxEiw4T5Nn9R7ArJojafkDB3fVeqXXU77hMxG4TknWQEsW3m4JfqT5KbKSmX1tgw
xScas0tlxnfeWfr2eU2m4YJVNzg8ZAjODogWPxbiTDWlJrztiG6kIcRg76aD+RQ/
aR44L69lkedH6sFxllWy7KUkGgqttUQpJ6d0dHJIyAzMxQut9yfBhan9bF+8vFeH
YLHxZTIppZB2LlbmO8C9dDInw7I3khePjJ9vFsZP2GjICkq0A5iT8Thh2c5aQgBe
gQgLzrYayZ4gDNeids31l2PW2tTmhwNP9eBguiqNtKU+F1zbE8ftWPQlQ/yZ8Lm1
dkFxzIydXN40aW5+yuekFAKll7ddl7Tzz9sCKiGDmsPiIyl4KKx+x0QsjnmBundt
h475LaFDtb3zW+qg5l4tSGG21A9FLXH0KD2MbcJzMd2I3jIFSBPc4FMP8ruVD50U
lOY51gtfpmN9KEeofXw7L8/kkzErqabIhQmBYwi4roQIHAyqG3gXJ4W5XhHYc5ZC
fNBjYqfITGshqesg6Lh3xWaKw5Lde3pvhJTMci1BGv4gcnkVlANLYaV1Pbn3kVJS
IitAbm0vNwkQpq0emwea9v+43nZfolziiVMHFTmCPD9ygn+0hI6LO7RVeXfmpIng
cdutof/KsxvlAsWd8Ef1EHrq9oWhWzFNjZ0FbG9TJKJgq0/jJFeXV5Fk7+4kuWjY
oLD/2XxIScWn+hkeLsHcPluVUXQbusDP1K35a4dFOJSOGHQ8FhnSFRu6AvBxl3rH
WQRZnFaGIv6QvSk05H2B6MCDV+r2sFuXpUI95D9I5lyHlWbhlYZ5MzNrdWJ5v7kD
OzXJVGTdwbbQm7mycyeoaFM40wNg5jH3iZg6jry8JZyRe84XepCVmLDG2E+uQxg8
OLaRzAtFAM6BWa0Djpoe4z3DD9qD9oJA/p2S5idemNh2RpHDAYd6hCooi2wQSICS
k9fjtvE88/vNxrtrhSeipetKl/ZqUKNRC4ZusfNqOgQhmy6b4lcYZO+G7a2Os195
GURm9rnC+tjPq/ebhKIBwV2D4vfL5RQJs+SIjJIqgOozyYROgmjYZSZOMHC2t82Y
U06Rwr5tL48xP1dbSz34wgdz0qI8vs6RaOhhIY/30ZKUNZMxvGMjRiO2jl3bbrGm
8AUhDu3A99uEtduIy+UDvQChxKnm9ISX6yyU76+/vPIdWV4Pg6UPLxfIZX1NvpGW
gBcSi9cg/Tbk2A+NIoLYygQeQREvocnTLY3EB2rx0Fjs9dPIElmHCC7qXe++CHfz
R/5uGUhzwdUF6a0SQ51+tWvePo1iCaPknYSnhTEpNzv35b9QOg1KNXp/G+xD5asY
dEFfiCdLtTVdLQF2zC97IfPaeKbLCbPaRDqpG8fFmRrGaCrsu4I78zcbLsAYQVYZ
IAiFvCNfKx6rgXlo8OP71XHb7DDb2G4O7bVE1elpJFpteYk/6mde98Zfss/oeG9A
dxNbnQEM3PrN4hUQR7buUJceAZ5cxP01DY1xY6/i10iQoU+cCpGkS13uUIdjAmIm
3BRwjmy7Xx6fjnddyetQIhaWyDIWtoBKonpsheYw2DN05NdTZPpJH3v33oG4Smnt
bnkaEFSqAC1jP1504lzZDPz57YtIDWm/ZioY+E/3D3IHMLKA3GgxvdGO3cUd1lYC
wkwp9r9WPfG+TvRDjy7jf1f9aIirY8t30Qk/Se0Sl+gAOAQmDdyXQOO+pM86GmM1
Vs1tYFk71v8rcGjkSLuv3mlRHmIjDEa69sqQf+iGwgmD7D5NJr8Va8+EQ81vYXjt
M0eA3iHGG35/t6F8N38cDMAz4im37gNlX5erD+/NorduUiZZbLf/no5RQp7jXDUf
AnMoWodTHgtBiXr0jyUtZJHAbuJWuWcG+Lur0OIviCEvMQPX+x/VvOFnOIFIDeCS
Bo/TL9jsgpZLr+XoXo10x0pyyp7DPigSWfb8++lVZSeBSLhyRTEgaRuhhSvhvybR
EZ7dw9Xtazu4h6WKGaxBB/TQQ66V4gZLrpVO9D5cP2Jjm7EV7TQsXKsktnLnnIZY
hvXqesof4Ak1Q0l2jWGAvlaIn+9WlmEV9KXhXalwWKo3Ejab/Z6jQ/RyHTIdzJj/
KDcI+Bt7rTKCV6ca+ORhqjMGfZuZGix0vj1EPCiXP2BOnBlLVbUIPOft4+1p1WNg
lJ2pDU3+wFARrgyB2Qxhwp9p/CFz2D4exBJ1F3Xbi25lmFZ2r897F3r+Z6LOEfvV
lDboFzt5Glq0cgUQusAl8+6svgaH90+zirb/AUCgcO97/F6lfMwZC6XrxMsXguut
If7vTug+sHINRG4rboC6kdcFX54Z0MEz155w3X7GP2Ak3alc/RYXOcco2wxaNX+F
wKFP7LaW+47+2NAvbqcPqm8Ao+pc4oiuUWO/jVJ4YUTYcAa6GkAfCKL15hGI0n/l
O4p9dKrAHVvCmJeHFW9haJvlKppWp97kXJQSTu76U2Le+iesHjGubRoYvaSUoFRe
6586PXKzQ5wpaEyIb+rtztbnDT4TJEdL77CbjQM7UTD09tDhOKYTLzVC1IO3EDQw
bHtdD0ylHK9rTuRnIHRsGto1CCYXJn9At7fhVH2m5wgbTjRWgnzarypLTlQGCU1u
9FOehvzVChKU7LG79kV+Xsc/KAjQ914wmSkjQnFjGTVQSrz+vqky2vzPntG+PqVw
+3A1bwwNC8KvdQp0LfI2aFTYzn5H1BSvve2ayk6sgD96fN4tezcvfUT7ac9Jq3Nj
LpKLBga9jpy0TpKRA39KhAtUvy4fLqsP1Tqg5W83pkFY2xCYOikAVFeh/4gv4yG8
sQCYucXc6uM9Ac4WpjoW/YigHDbohRUp/Jw+0rZQ6KnNPFee+yCWEwmNEpFfzXmB
iIX+fyjMkXuw7B4j9IrIzB4WrYk3staNIQBOmthJ1tjvNdiuCpVOcHQFbUlpuksL
6CwN2qIzeDI22Yi4zUNTEhtUXVrrdzwNZlhvANZZg18N/LuQ1i4EYQhgYasrocDi
eYcngeCFzSy3ixeEtsbnL70+sRkKOeWDZFCFqV/XfKV4JB2BtFPQruwjpc6WuF2U
wQ9HrpmzfqtPmDxTjeHAi/pofjUiSTRsUg+9Z2p6BeVdjYfZ2aBIKWa+nvT63AOH
G78CuwMnoXw2orWguVxH+YZ2YPhTa9DPbEivntABCnl0VlTH4/jY1yBXt8tMJPr/
YDPHf4shjo51DTK0nWXtboNOyUUjbQmMdBIqH28qyGkGDh2HoqmFz6i7y+l6gs9v
YXuQrHNpXCgexMXTc9dqJ9HjuGfVvG3xoXi3Jj09v/7usCBuKRi0w0EjStPuUQBs
fvGTqr0A13vuFUPbAHNRgDK0i3PRDB2ZP8AVBvjr+UcDOqDTKLNAQCtYGPNxqC4K
awrkVV2uV033WWRb8q9jy338Lr4eO5jN9L70XHr0FSaQ4yOZyOwzUCW1Hl2FiRMM
DWmTGGprTnzrJAlQFmJoCZ3QfJqcTE9fckTWACbOMCbMzY6w57tZTHYQh+k9fcMP
9qZVYUVSN75PKIux2gnVhNZNaE4owcqvS09Va+xbrLUvudlYnaAmmUdl4V5t77C6
UPLEiOKTqoUwpJ6c/L+aaKtzHkDY6tMBR0X6ssT0s8Lb7Jp65W2IzNg1i/wNeQs1
dBAVQsLInYZrgq4p4lodSV4OXw3xX3GrIDG56SkouVSuggYZowwEVHOmaRzX/6CS
aktMxtlw3bjH5ZskdeAqbAX0mRrenJV3YU3JrqjAT1XW9eVA4aPlPjqUOoT/CmKQ
dbI4sIEhM7UIK3kGOj6gj21/JUQO18Ba1UYs56+io6QkrTSzjy6nEPkqgHjgtp5U
p+robwLIcQ/CgQFKWtEiO1QwtcYbJMU7C0NQeyPW6ZRgf0ozOWDB6ygQNqL3sc6f
6WzpZAVWzNq5EVGLdqlOcLUxvvlbn2HGbKIHt/5ScyIh5SmxtHvyzC4uAvCDqbMZ
cfJlb4MwwCbFO1Qw9WNEmfUp+76CJYZcf6YV9IDl9fkzxQBoQXEoRcP9d/HIP7r1
p8wEI//7Me6WkFPLeyzznUEOgNGpAPicJz9Fd5C/2FHs460K+6bXHFQNbutTqrwo
3OeM0sNPT2j9elbvGjOPet3l5+EM46eo5ErH+nBDyTib2Yzrdlqp2a3wh2WvfydS
SXGqKu5cff1tXSJh8V+40vBV6K/MPx3xSy8SPFSvgnXeiJDEHgPdoqJaVnkJNx4o
kDDH7WuVTas/GeAqtCnoU6kX+euyLMpaX/dxq0AbGAqhSGhoRlEquJHjxE0SiBed
nphwUAJN0BiGY+8fUdDSTNxiR28i8OqbAscU7vjcJ/6TIE6UqYD5fa92Pg2rI3bT
whWInBVtRQ8UTzBkzLPijcPj9PQ7SB8rx3ftpyT4m4ZRZaJRCKgPrwgWvcQw6Rft
jUy46WiUdsSOg26sgGXBi9Ess7gBX9sw2NOk0wMdKt5+o/745JTpUK7fLIL1lmzh
TgeAV8j2jm/sFdtA4Et5sKManvSWh3LBy6AdwwlixQ1ycPx3oK7MYTa7OqInykG9
GejvLBr70hzrkp0vX9XO/ji9cJxeMzeUYRyI5oXpCr/720sQOdiITnCEG3aBi3ON
J9NPnEiCBNJD3+yvP7qF3OM+oKOWb3XdEy/mwd4cc1VmiWbP80lhPsr0R+SpFbCt
vbDWm4MoPWbHfrH6R+XbrIkQcp6TqiCcgq9t2EsevB7/iK54nSlkxAm8Ek0nzh/W
abK1QL8vHsOUZaOG2P3gnuzyl6/K7veu4t+NhLELRjYQFbi64bT3A9nJI1IIAhEl
IQ6gicbzyEAY2JqWzLgGStjDrGiyV1UuqfEjzHGS0bR38ZRS4vYuhcLF7r4bxPAL
zScR67k2j8YC2itSC1vam/Wafwrj+H3gGdl3cReCmdZnN0ZSl8lpfEfPH74viS7G
sWBs5LuplQon/I7junzvmAlLlwWfHw+mjZN7rXlLDb2EHvq5KKEqJ1laNhm9nTj/
j3T51iX4D6MfgfGztn3Lw9L8JE/BaUeuNesq4Ms/uCg5f8726nCR0AE4Y35g2wBq
XYd+FkS2XSWRcOWBfm/an7RUo4PgWNDIeXNHp28OxwP3tV6A4VmLuLwu+e3obYuA
7KOAw2FdpHoZ67JupSDkvIVIz8I5Jsk+31p/YICeBP1i/aWrrCI4RhbkG3VqTYia
nsVHUTuk8KAzVAsrb8+jRPi3N/LRjfxE5lm0rqLZ3jTOomVe5HlcHfTmCxqtv2QP
tfawtcjFs1cFwz7LjAoZTQB38HVAIZxNVC722+1kGkSykSGIVTslT5J2sDjyuTZD
Nef/RBeZ8PnroLZn6eeAe987GJwLEjC5hhrhN+5mN2/A0S66TcFKNR1WkT//Xtjl
0EoYP3ujGy6gDUe+6aoMHUMZW/p7ABjYGR8pugAxg3RaAZruuPGHLKcQJMpLIn1G
OPcMvItcmGSU2X8vBq2Gf8svQjg80aExgEoLtZGmX4ghtmqqjH/iJsIvNQQWDLyh
G9ZzLAl+SBUYpe6NXU3hsoom2a4eq0X2UMeNYz7HQrWynXi+AIlcOb5xahL0DMH4
vwzBUDQh0qsBlSpRMJfNg/4D8FKOZk85fEvvMXBYJnrSfwznKw/BLxkufR7vQmzl
KF+lmXEsLyt0ndynTKzfg7+IP6HD+eW1OKx+zG716ZJDHgvvYiLRtXpan9CqyU8k
NQoUje/qpam9vlY8UUGT1C4jnxEHV9xLpUbBwRBcnNdVESYGulGcmV9IWpgo5GRL
nTXaTlSTCIHPagDBzWiYlWK0jU4S12Vn59zBHIMInKoN50QPPaw9R4q9gJrqZ4JO
2QaejUIcaUbjK6d5MmIJEIz2r3YeDHDFpaNzihRFUnV9WCXcwNE03crqkSxrOY9n
JEhWESEozZemwSyrmJRffSwiKKtNpeuklYGDu1f/HwKXPxRmyNYGntMI5C17ETzU
N0P3HBz23LDNLs8kBYFxb5xNqUJcLCK9cGnjTQyHb8ZAbq/ZGoyuN4wzSVrWWCe1
hnLXlN783sKS6Em1zPx7RthMxDNb80VleTOj3eFWc/sw1JQdDydhlEo2pHRIN04n
Mqge+hWKpRt1tqTtIQlIcx08uExETvEf9cNk3lUNCyQMxcfKokwHt9CGg1JALtGY
EwvyzrVylWDZMmc6AaGcY4jHaSLGfsa/O/8iaAYObTNkpq+gqNCnzGuXa1JmqK5Q
eKhfs6Kh+I5PxrxQ0y7xxvByXQ+d8M9lNf2qfeKIh9S5UL3a5gE+48wZUJOB4Lqu
FCkuhXvAtr/Bq0Ziu/+EZueV9wfE0/xILk7LQx/sazqfHe8ykDn3yElexFemdPKS
0MGO+tD0l8ah/uVQC0BzTOxgihiKTz/Qpj/9ilUID63gSJ4HnO3Yd0VG+Svk3nnH
ScI5MX7nd3Z5s2noFgJPcQ25Aq+M/ehBkvD7zElW635EBgJlkm3v4KAsjNAbdnCT
nXnyul01S6uJFOeHpSofLhwLys5AKx0GQj0pfEeclg29C9ffKVD2z6uBkBPeJL8n
/sstueV+rAlx9G5S+jZBO6IcSWPmgonerNiRP8mE5lPkyocV5GDrM1XQG5UDQlqD
sijgNP8gPBzwZYbptaiiKTarSOPy5OMpqWcZxEP3K2uVfgTZZWW2Db6l7a3UCtaN
gYz2CqK9Qc3Jjcv/tLAMUmSwW9uE9NT/BID7yec7fJXydwsrHwXQ31MhnjJCXdy0
yLOej6+SOlUyiM63Wk2olnXeP7/qKaS/Fv90IP8iGNDndKXXs2CvaQBWX64Z2cKq
ebuxdCHEkITrJk68rGEy30C9NvloorE0vUPUQdPNo9p+4ejSuUH3T/OJ0HoAgsIZ
A0OLyOHKXBrcxwt9+gQJKqsnEIaQGfZVy4Zcxy8wBogEI/36JJob98DZ9jvJCfd8
RKQ9FM7daKA7slMaqQqL6wE0MQY6dAsN7T5yWApcqJjwy++h7cCv3QSbAof0aqhS
uvZrgoagjFpmGm066fLtPBAb3CgAUHJLGF7Dr6SnNWLlrOnBZ7O0ujg5i/PKKnyi
wkjPerRSdgkKdHG+aG5YekDSm3EvcC4ENlP5q6ByBKn5GyjqDf2KgiqoY06WboC1
sI+5O3H5I8ykTynSxYTwD1ZzaNJJdPvb3aqMkrxCiDT2f6CCjWgYtk5+0MX/Yi6S
m3OJRj+VDOouBR4s6TDqQ4w5TF5guZ94QoanRC/pPeTr7siX0iP2tx1rqQFtTD6o
yx5i3fgKRavyUsBB+eKi2wUH+wIplJmxT5ct2/orZW+aKRZQ7jKP58ZO3R3HvfQI
7nZFZ83sOpAn8+T6EAGoB56mRpjLrLWrfkzbgKbjZCK0D4r7x29lTi6yEzJtXvRH
xbOdkIuOQEic1HPZe+L7g2nYs+C+6rsZx7C4T9GXyqAE0hYhsCjFEZB72VBjYvC+
FbOymyWZkXZ3/TXmspCcy/AnlLyHzS/F4ZbczGOtAgAOfrOjzAHypS+bOzXjDLuT
c4ks+wXfI68bFkzG1FtJATXkpw/BxaGZM7U90UzwMXwFZ69KVCvADcRq4+wBYQIo
RzoSHy9i27jrhO5ilJZ2FQCfBKpvnWNZJakaDqHqX10jXcnBlhT6enzDlSHEDQLs
c111KU2rK4WYfhJEDZaWHTQz0r8LSeZyN0ZohJLl7Rs25FKaaY7oILt4OGfaSTmI
r9rt/j3NS+W6u/q6leY2n7Z5lcAm/oPCo8n4NoWFbnzeR4LBa2Z9zT28QSPcC1es
ye/IzmfXpYbqaSD3WzsEHYYrkY7qneitkUY0EdURFUV4dxXmPccenu9EQ+uaBMMU
T5CNUv21AD5KL23WdS6z1BX69H0AeAJBmDiy891CyzfXa7EuTWrSLBgHc3iocf3U
JC+2k6XaIUE4kueL3Gfg+1omi3a3z92TlIvGeSEFe5YuDkwv+qpbLbY3Gnm9xd3q
4jgxBavOUZ5yiBKu87NFQQS9N51RVrnIxQHpeQp4Ut2nlHGCY6a/Xl1fW4ad3pYA
Qsux+mOJ/SFfdBai0R+38bcJKsVK1zLJpOfAeb9USh5bZQuukDj1nJGa/cs01aKq
oC9W4Hs+XMyyxB0hOub8TofafQObauhQP/K8xvjaREgnkfO6rdyAc4l6DV70MGrg
GQqHplvSOIKRSYPawYUuFQc9OvYtvao6DXDg0wjPl4LpfbkP329zW4l3YPxF610b
x2g9Y3AYvCvjA/gWpWU55x3X0r+l+/oiPNmMjVBqhJtf6AYHp49Kkc2+oJbIEo55
lZbYjBNtb1jwGIbth+K8oo+C2j1AvtJbXj5HcWDY0/56vMDujzlWuXBDkzKwgvnt
jlZ7VjBLQcLluJ+25o5XBCKmy5L8eMkIQNZtBreV8Iw4/Tp6fOBziGrblpysQuuY
vKyp7ZGMfwNFtO/Wilaru6eFyHzpC45zCB5X4y7CrHD6WOaz8UaCQ0+jLv4adPUO
p3nNOH3T729bo/f3fBLdIvsNNdUp3bb96tZPp8hrSSEMBzvJHeQWnpJ98GKSwm3i
lkNGumQSa3FaRpjIZLx3rlNrwPe61aai3OE1UkEVqnPy2HrmxSnMmxlkTT6J8XdY
y171ba3pFOBhni/7kUNxyY6FEkuz+cX3+3gFccmbwRn8JD/R0Lu9yAibenKBRqwL
DrNs0FO19gmFrkOt/Yr5NFeM1PyYRkQv7Glb1rnjxombGO5LP6TTxWzG7yM0duv0
9QdSDfMc5RkIjrOCcHTwpK4qj2QXCEb1eYjZgxsrFoAQ3I9UTzkK4TkTbn7Sx0L4
kPvCxpHGHTXkJ/qS026ToTGUxlHhPGo7fAKFXLrNhX4Bf8dq1w55ggRqx0T8T4jy
38Dvg+54Vs3HZgEecMkKrgZ0gkBP50tagdSOe5uhtbeSHPMvAKhBA9tc2Wa7i/pQ
qRL/0ENdUK9kXjM0tSR0u8byuhCLfdFAJ6Q/TX3HK9nKeKUHD7t3dHAByQyxPEuc
qJ3DBEtwgpunXazDcpoc2cnASRdh+n7HqlDKA+OLZflEAx9LamrawyEnWrxO+qJl
Yh7klCw5BQwotlgEk2JShCp/mtxibxuy1DjiIaafj2KXQGvKGPuE5DEpBcdNhroP
fyJBZlxTdApMIm4Ly12e65KyprlUUAWctb1c7UhvxOrryekHR+cUr3lt+RJ6lEWK
nWcXaF+GyfdRmlHuIKnLWJx571eq1ruIxmsMqL1SzZSRaj84hh7pzXqq+OPFg1XQ
kiLw9E8YJVWIQlOT5voh2vP9BOKeCYbeV/19snUluQc2eosJSUMtVA8pAC5X2JzK
OLgwhKGFqFLFOiy2rFmqeCjtjDN2QrTHd3frQ1if3GXWwp5ITJ9ui6FiHIDYNAbt
4xY7M6nfz0wpVEsDgQtVIwaSr7KvQ6Bm8H3bNwN/KEFsX8SbGHKDwii3gzEIe/x3
4OxqClJ/+0JB37fXtiyh75fqW3LfqFVxOJnOxt781S6YABtTqqOuUjxhY7gc3VaB
ooes5/ab3URLtgIX21S2xRI4uSi9GNs74WBVXzE7fsXJ9XhhLcOD6LyJoyKa817R
kZZYQp0NK9Qr0ala6rFTGN9yxi+8qknLkfd0FRsGKlgX9tvqDWOvkonXcEbUPNoJ
8p+ADNyyBA+fuXSYs437IUfMCcV0Sd6NPBlxS62T56Y3bN2HFQjOoy3hbeTp6V3L
W0uRtB4XFI3YxrDoaAJOwB4E9K9N3jv7TZu0nYew1Gsl7z8bOrgCpnH4O2P/wsy7
5doKWtngrOTZ9aa/Qp0SqhkYFLQrOKN2rXfk8SRlnJdogOYXq/mm16ddTMcD4u74
7vKmI+QUF8v3Xwxr3evEC2kBCfLMtdomj+aJrEjCSwGjSZzrbktYq8VhsD7EKQS0
JpOSlznBaoU4S5Uc9JgeAqum0Ct1Od3aAzYsQDal9BNmRgIGp1LWqgCc3mgyg6ui
wbmcwOxIN3NjCg6h8RrIUqr5kyjC08sQECVdnh+m1uzRw+2Yc2ixadAFvIrMhfrc
eDuKbiXPJSXvpOQp9OFqYRJJo9WA2+r1aCDwWu0ttRurh+mdz03i6YuqoZkNChfg
rYTOl0FfMj2whR0qnSo0Ay1lgqtEPrf52KfATczVE0urS1ufO43ITgG8i25Z05Hw
oWBZUqWr+etUrrGaVcTyyqLCivHqDotIl5rty7n73s7oJpp2AwIKcaXpyzZ/EDsj
TpWF8U6R54wkgMRYcer55IegVJkyMOKXQnG/f2fZgP+a3mxtZkQScHIGu5T3CHvS
Dcm8KsRn02vUXpIdENfb8CYBacALZxCp2koWjV9PBKBUX9rRX4HnskFDKpHssThh
vxrPJnf9uDSy3rhuPgwdps2oaQkimVjR1Pi7RAgbBKyw/tW1+VDAh2Wd1j/nIDcg
oMEnNV8CQ0amluVJg+TvaH73P1ns4plSezSwpafimQtwlSXnXvemuLYX0OTQxt3N
ZLPPuyUIpCu3c+IZ2Z5IjrRlwsuAtjwvbgLBY5nmFXm/ZUpV6snNHCGlf/G52P2j
U1KtH7/+/ZYSXjGQgOLo2+VUaXvLrgnc8YznESK0qh2bhQa3o+w4sOzuBxVdKkHn
N/sxjcobakfem74wbg0jajlAw8X/CDRqB8ZzJuyawPhtYK3TP5h7pbh7Zkl2hofH
o+YQMghtccNxA3OJs3aUQFCuL7sY+7pStATSFSJXUDeRpEMA7CYd1GYdnkkFxpif
KskcIga09bFuJ9KTXDbiqm4S+crRqeWkTf/84ZUhO9Y2xUGBrDeM3lOWqjh9H515
RNpNkr3bvzt8P0yI9K5Gp0yL49QC6xs/Hboi5nnaeAzkL8CBl+ln/RMt3gDtIJR+
zw/7aMDSVSqTW/uVN+DZFAZRKo4LS/4YojPFrWtCHl/Z7t5T2bePfUChPBpg33ss
ai8W4AEEIeILHNjp1RRZsJzLKx10kCjvIgG+6j4vVF3wQmyNNmjXEH7/f3Y2OgxU
+kmP9LPXCAN3APa3N6jv1VoIOMNQ82S4lAnVQ+j35tmt6jzuT+00p4Z2GxqneOPv
B8kJ1aqk7rTjJKvRm/i/mdvCtjrNGcMz5m/hZJc7ANIVGZ7YgZ1EcLQ+t8BAz+P2
e1oTwXkw3or/8jPfUNZU9u+bXeoercubqAIZURMuO3jTfeZQwUqDYtRm/rs/iN2v
jo+/vlWlwsi1wq8eeiKwDDeqy1R98nlCOT+3Cj6YQq8HBWSKUqQnCzFm6r1DCBUw
sTTwr67bHX2aSx3EryRsy3Bb0k3jnX3L4DbF/5CUl+PaNVeBMWzHvh/nbgmzkp1h
hnjawHkOE/0435+tc6eEBFTrWMZ3aD7h1JTtCV2KNA3pUnFrXmGONnpRRvVEclLp
ch0/2pEl8bT3G6n3waBpuKcLPkGVhNhsJLGIDW14SJ3MRB/vHi3MwBTZ/3zI5YVz
wazUFa//FVYkISFgYn9yo8fG0NqtpWG3jDCNHYJmlL0tmKVLXgUFwXAi2He3myQ7
hlNEa03OoQGKey8da4j1GRaJ8czDTdUzpiW54IoabPGIRPfXOyTffhbqR5pxQRNF
rCkvGBdk/w7ajFVWSx7L1A0sdtgUWyAlRqxExK+AGiZGiBNub701ghMfXWCGaAZw
pNzLShJPamEwyfuKOdaBEwBHq/gyFy8iGJExa+NrtqVb0rL3CeeecFh64Cx1SdUG
LU9lJiXBnKQVZ2DaT9aZ22WAfY8tFO90GFgtfdbFsXHR86M/bbb+9T6nhluTRPc/
Sva1tI3n8g5bCokW5gWgRGKkQeWT53aTWvyTvI+ILCTCNuLxuVYixxND3SNM1h/u
uFNDatmOEW/F0uIZOuVoGZu11ofvKzJ72Y8dUOOHS45HpzsaMs4DwMizKZSTOad3
9Tc72RGru5stlG0eacp32Yhumw6p6/hVaNo654P29H/m/Gf1BZANgIA5HPaKq8zC
gI4/BQ9UerzQz0eCM8mCtlo5UzsYC8bgCo3Yj0V5jrR/6Pih1dhcX0AYsaBPRwPp
fDKzXJiSdOLQgN9by6S04YPKSW1l2kG+D+FkD+NfMwzKbOko3Vl4aIcsxYdwigTo
rJPYkbOEUB4WAtLDtar6yg/em0r6kpl+Tn7OHsN0FJROnQ+iWbP7FMtVkqbDEwAk
RjlphSFeAyWBSx33ZPw+3if44tB+icjeQNIHyRZobMP4Ol1GHiEMRD4QZLneoYO4
AlKh361XiPn6amGgfgWxIDM6zXvHmUtAbng1x9MHQkk0Mj+9nHH2S3FhNgiEUWvu
h3lF9H31eo+/h8azfG42wIIEAoTpG272Qcd1LQMUtcANDvcTDYLIJAmc/jNt8Xeh
PCiTzdi4fUEPvuHQJvrWE/rCWeOIZlqquEcwBpgNxS14rXmJ0+6zj4+DoE8Cxz/l
UEg41cV4mmMvoEN3QQxCF6OdAaeGCKkao3C5AK00uNSb77vnUQKa/zCYdsgTDqaU
5qyTFapjqYOMVbTNf2vsEoHKWdjhz4UO8Z/s2wUKI0+fdIQm302nlpHVbeIUN+PO
amN5lX1dyTOD5KWaLEvu3+fDqUfKAgqmD68RqUPUJXKNyvLiuK517uh335NSZzmU
eK+mvQnZb2kBEFOaoh5hIohmcidIyiv2dG6VClgnEx2hKuiUOTz+LfeVgwSl6wEs
2CIwd778p+wxzpkjV+M87m3BQgUqDzGBjD2YiQwW+OK6m67gdAtYn4QXVnpCcg5L
KiepBwDZGYzwnCJZfidbr1bU/GMfpdpzjm7qOfU7yJXxUaLSIWGLUB4RTuh91oNf
TO2QGzAZdY+tlUB8gEJTHryorHM5Aog+6xohoW5dyYrXH65Z4zNl2gr45r4zquzj
TSur5o24Asb9o962ebgqIwjReEzFwcWeC+5vMkuKt8EJP80pl8dab3vqmetF+b2m
7YidT1N0WsMXrjlphAycPfUExCKVMx771TXGUF0FrdrqKGK6Mm/lzEJjC8i+ALAe
CCsAz3Roc/QbY8SVRIfBu7lZQuLazj57Hq6rwvr8K3Hvsr/2gRDZH5YWeUB/uk0K
mAp1IrPa38eYHbmvh/4188UoPz6/eUWEug2j98ZKF8+/gqCJm6W8TKsMS9Cv5e0H
ASw/Ff1xwLsfoo2HBaauWEDM/UDWflEXg/dSnfvrFg6GCl9K/vyTU8kdQJO5Vspf
pL76Nn691BkqopGimJLfSMUPuGzRcVmrYY2gSMH7L1GOfCLF+1O3TVLEIKvXosSu
/udK2joIw0nSBd/Dnd0uJc3vH631NopF2CDLxgzDQSlp+dzXotulO32gKu/WMAwr
uLTsqM9LJ2+2TnM3srJtj+T42avRZK8RpARU+Ed2hzIbIP/+X4jkOWdOmAk8j+Qa
kEfsFa9Cr2Wfa0uSjyRGdYEaNjT51rAJCnCHFzXdtXtzJB0SrXNa5X+6OmUYWoex
r+qgiS9ZkiQED261LNvQEpFPu85wMCxVzSLCNR59vJivS1CRKiWM9LOPjxM1/1Hu
uj6NvnABlm4S81qZvGOOoKRrxWxSdoen5l4mHvAQTppT/QUyMqP5J1frF9/KoRT6
2A6i/PUiqGTt5sMpa1BjTqZt5Fvm1o5MLw6hF6LLHybl/irpEhp5rtZ1Et6c2bN7
kLtuPHtRX10sD9s/+GTBZltz4j3hFA5LaZS5oSe0+mmjzxIDvZpZp6jXQrvahL9U
jXrANcamDakR7FSkGudYnjV1q6jWLDa7g7e/BiiQ4yd8RFnKHoBVlwlSF55Tose5
EGujMW3r7TbO9gighTBR1umP6S0B1mAQbxgGgej9XphT1JwiO7ZHNLxH/UVkIGN7
gaq63tn17rGfDwX1HZJwc4eAtNVdsCPxOPA2E9S7HaLZEKaAjCTlwlVEF2bvoUTH
1myOK/5xBnUgStDyKReHgQ+80J8vWJN/RX+cbKeeEeAwrxUJRL/285YGP5gGSet5
ZfCfUDMVc/MRqjPZZcl0XJR891ckfksmFfK71odLdUe9SdpjwN0KGUU8Yvz/q5M5
BHVdPxxu4MT8jF7zbBtQSQTVg4bguCcHUCVPC1EKsZJbvhfr678jTxU0A+C11eEH
RBQ0+rbrJ7aqwy422eY+z4GdXr/ks3Tzq0wqKeWT2NAYg+J4rlKdMy46WtnTGiw9
q/WmdsGVsf9F5/Qhfp8X8B80/yHPy7/DgWxwlmq8/yQXyhR7GFs2CCrHR9b+eFDw
PXJtreWo9yRkgXs5AFwFuVLwVpl5xeAScUQ5Dtt660QeFy5FXawoIoAYiKoBJL9K
AfkV/+mpuQDoMB1FhDiyp3Xq0xhPhGDPJPKrTn/1RpM9pU75OWKm7MVd7BXsnt+u
D1Mi+t+9ixINs5ySXIOBHuAHZRL6KJ7uLXLGVZ585FjXsv9VKgnhHo5ozv7z5NVJ
u/VUOzUUOgmiykH4I5x0CciIjWjiapOuOtpU+pZmCz2Yn29CIFijQJIWPy148xeP
iwneMKkY9ndTuRxjfSb6/gVaORqsLoxunvGWqZhPcRoY7Y1stzyDLcBrUv2ru/ON
VTbeNKBphrbWy5eqEsjL99GLmE0CCYqzGygk4eUzJJnNwR2yQam1v3rgbTWJUZAK
+AP1MyL97Ox1zmSfdpnvpg6MrSPvl+iVucUOL1oHWINeU3JSm6m6u5kt6nAp26J5
SsMdqLRQUkzhzClwvLtPiDhACYDodoeAcjtDtdrNYr6NMRT0GGchwWn4Oyg/xDJC
7XA/E0eAtuCuHCyUqCCEiKVyHTC+G8SB7oEAYoPkqQnWEoduk6kIDRk6FUMdaZoZ
P2kQYatuQ4J7Bks2gwDGCPiHhDULmxSF4hMwqWtLm9JWXiy6zrxFSrJIq4srSkNK
VuZiA7nwzETRTRAaQ8fHGQ8gpbPteoq94xGq0luZtL/BS+et0xsZuqCT+PZf7tGW
GpxzkA2dLsiwNhGmrIayM5LeZGuNtwVv9eKOGtnkaI8Sr+iCwyYoy7HaH0gujJ4X
zPdIQRqvTVmCXR3Ps3y61u0xPHHVqHMmum4/1JRnEQc/Vm8rDlGRiw0B79R8eKnC
57vBcp7JkIDudYm+ZHgoupzX1+alQgMdQmsAlVIiBNsy5Gd4aUOhBj8wFG3Bn7hK
IXYzMCtChE4M+4mrWwNGWwIjTAz8Fl4a6al2SQsfLPOvvNwjR2asWhHb94Sc5ENZ
aCJe5KqUlZeY/InebPKmIBWel0yLR5ruAlCBUwchyk7rFalImHXTagBJ0fX2KuUR
UB+gNcHIWqIy6tjwTw0NBSDtwNAe5o6xz8+s8OK8c5pj1xnUcxwFfz0PEKR5c4wJ
JONxi4+I7AWIg4BAuk3J/1uU1yQp/uoUd7VTzyFxE1tOxoS8qls7+TamTZThBirc
HL5nnQ+AXk1Tvw+4TlKunmaQ4qVcH7UmxqCrzXeNJ+u9CDLP0ApzXTncdcQIfP6q
WTmthtMANEpMiVMpYiBYjfXcc5S0U30L5so+WU7KZXOhs0eiZbPpdRvJqA6lFGD7
arc2q/qBzYbDnVOGat2yd81e7EC0hj4OHfwuBr5zl+Wo331iw6KVQ2mJVbDQj/8c
MaFUrGzIS5Z2wrRJJWpztT0wwvYecTnxhM0PIG0mFMuPewkC8P5R4quev2UK6ejB
VTv4du6ld7EThCjM1CtxnT0F88q0sp/aMG+5N0YEt3lkPqIM4iIPNwu2RVIbG6q6
ToyHeIj7LP7wWakshqlEE3zLRLtqNsTa0U4qHIcwUgrllhHtE/smhxD5WZ9F4LYL
BsibYP5hA4b1lyh/X2mJhPPM9wq9VelxVBwP60MbrBMju2HqI7ovljQKvJmlZx8q
e36Ty9l3kybt9+a23iGg5/Ei+bnC0pauQ9mmO3AjKjgcjPSDFwLPmzGtdCJQIzt+
+pW7MzZss1tcbO3uzuN+LRHiUl0CiqBtsi5wiYDO7ZA+IwhIkmsg9yhnBXfyAcf2
VZPwaCl+J7T0PiRMHit1+OuG82ZkYL+N9DomqcjAonvFegNRCBzMgL5p+YhoHKAJ
mZbaje9/99hdkcbAmkf0CrijXNI4E47Hzki2qdVsuK6j/U7krYmkfFHwhZFZGps7
JgeUtmtTb2jyxijk9c3hkpTM57rxaBUrjLviEAnWumx9Y2s6im7E1iuEzvBr8Vy7
jluudFXqyei7oDE59wZ521fNYXhpkBcjlDDKk/wM1O4AVi+9WuiQMnqjlV8sRHjz
O16CLeZUKvqb6laFM2MfqGNoaVG0wD6r2VYJ9IC3CBUG+8KeReddWOgslsEjgivt
OhuXWX0Tt54+pyn2WpZM3kDe/1t2yY5Gw6cGX2fzT1iQOpSIXgcZddjb7yWmjSI2
eIzG/BR3TWuCUmWLgEnTZeot9+gO8KRDW/4sfD8WQkcsDAsnT9ftDFwUAnhcV8jB
YOFhgUTqSx6BNBn2i3UqvzeffWxOu5Wg9WATizIOnd9S9q7bRf7FFFEASBmjSL0K
ejYI/NRbhoX2mpR0bkeGQ5V51LBoDnbamiQe2WkgNpjuQvXtRXN9Gwh8TFpQZVPt
Xdlc7AzG5LwoPnVMTNAEHbWONSBeBLEUcKS1uepNjfJ3aDFQYJllrzAC8OKajT9d
4UTrWYU+eAO9IzlEQRfnD/fzYWrp6b0Do5sV3zj9edQdaoE8MVP9qqiIt7GZc/PR
xjH4TNSrrpmnKWlkIoxJ3dl8seTb0NLuAW/qM9LF7lk6wM6f53I6vRSjTUYCM0p+
fw0A9ICNNVNZ7ny4+0Zjr8Rw5q2q1umnFoMFcpKrkCL9OH1asX53J5XwIe4TJ8W5
V7Sfj492hdnN+YpCmNh+hVyjfjt5W0634s5Tt471FWkiVSPROGN2WmpnFU1E+2Pg
fY0GkhtENOqkwkp1u92et5rbE5vKxzQjTKq0AQou8tJ+xnKD+13oBJBqdJbdkZw1
yxhLa4jAvAgGU4hl/Prk+kOgHY+zEakfDTE++arDXlTvAlV+xkSOqU4p0eXLCQFW
n/bPyMrTcJ2khIrOeJPsx5cYzumXnhal71O1gny4WhpVe80GbQEm2azU7yQcVy0j
1JBLat3STnf5IiONfbCCDZc0z05QeZiWDNzGFydHiKUhshfxfehN/UWLKAe+twCc
1xJxWu8jN/yR0/ye0OfduCWJxS9QAce3hFbKTZFUrdNubF1Mo4RRxQlp098zK9xt
hIzuRx45TOOh1Ts9+IJPzNqp0jL2NCYTnYQ7l8PhC1ITzx41Dj4ZwLpiCJrno28v
k/CWSQfMxVmgmEjBfKfVKuAm62gieqk+NfasN3XdpgZQ5X+odHwldYm4uMAO842f
+Sk1lioqJCReWWCzZHF0ykjb0M2Y23elC4e9jXRl0UZuLijpXxKfZevXquoXJlBp
N6ZEe7818pMNhSbX4MRmgU7illseADNz7oo5SUnQoJkJUcqe756K1cH0oaKCRF5O
vkQmjmUAYUlid0WOEvtnxCJJSZRqBta1eDy7kkUStXsXin6alOXCnGjNK+pn0WEx
5qW8BbVe9tEY5cavPrqhPgrSNop6QMvFoDyVpLA+xlrX6fZC4w5RXedRWqvPbRRo
yEgFMNwmNxPx4bN+1gidD+UYM0DLY3kMDIZgcgMbJ/VH8b9m6h4lqj+4uR0HBAZJ
yKfB1AkqmuPzLktHZGJ95iIfDqNSp5W2hPtl4CO2uARMqs91oRFf67RoAPCS4lIx
N/XoxxTDI+xEdJ2oRzAKcmSG3x13eMTyL/JkA+xWwMdLdUVxwjH2TSGIMuYd9SGU
ZpSfNGYkeYNnchk1tL7wKb07YGsP6CVYHMWOhnLIxPLn9YzPO6LBrQIIIaGVfco/
T7JErVuWwce7Lkshk0KupjOQfl6AcQ6DlTG0asU7Enmego+1vs8yARGFlScvd5CY
gc5ThI6iuNj+fUp7d35X3Xp5X/+N4UmOO/zAY2rmcFshcSIw5o/O7cFQXfeyvRmy
m7eUC2TTua9biQHj06HdkD51r872uut4cakFvLvmcIfAXEgwnbtS87HSTChw0TDG
F6TrP1ysQnu4YuKFSCLlEzyC0K2hO8DvI/5nG6gkf3Lf+/hR/zEuyh50JJGwParH
79w46AgFIzATYuy6Lxy9au3B+xEa3HSLuaNXDVcTew0sQ2ZYpt3bFGwqPvA+a0nb
nTXVXXGPvaAgODmWAIG90smcqm0/TI/R0QSyxDiwrVxIcJnaILD4GiZb+zKMOsxY
t/Fi8f7Kx1p5MB282/vHvbT2fEepxQgUnz/FWtQK04JZovZ3VAs0n2D3QxO58bkO
xBA++ZaABPXCZ+tucTd4ODRLN5mnDiLxstvIA1mh8m2GAPp47kFmwBkMI7zGez/h
g/47puCV+yfE3TnfHhuLeoGYWsAE/VIH9ILDUuvW390i0l4DaCOSG8L5aiLmhF30
Uf1lQDXEpicRPBD41WJqZzjRoi4OiO443sKXTpFXK28Dy5Zsllx8Imli6K6GhIzn
oOE5hyL83o8n8AfHkLKp0CkgVA3EXmWEqJphvyakuZgxRjc/Pnz4+vdFrK8yvWBO
8km+QJHY9VxYLd98Blni/pcawInNHaopX349g7ByfiGCpuujU0Fp7zzXon2EpRIO
7O4iXWAjHbJnvnOQouPEgqodCUBMXMaY9ET7Hu/R0lfAqBMmxzHTnHEMO8RYAeN7
J56/1Wp05zSPb/m7PW2lH/QNXKma3Z5bUHP7ARmDwkeJA0wTMjNkDAsvvuX9YZT2
lyVKjzPR1nk6U4v+Rjh6Q7ZkmtbQVXW6ytcnrRNeJIRZ6rsA3cb1u2fzlvcIepwj
fwPa6+0nYaj6xBWNBhOrgLYiB8m+wQ5SeEjDG5QfVCbRBl1y493NkuutmGsw6KqD
J4tChLd2NMnutOZMoVXOm/8IuxLQkFUTFNPudshKNA+a6LA9NexuccJw0o8ww3xQ
GP0NIfL+dECuVYyF6GqzX7qS3Z9ll328bLhfDgsvvymHhjV8+vilK0/tmDuWlEqZ
iiI/PSFO9Igx1dwrUl6NZ9G6u6s85QrnrpctSBtY438zlIICm0IHhk99zm6u78XL
JVxxjIT6TGD0RzPaO14LZSY8EbfqERR6nz8KpBJ6ZHTG0K9PAdbGtcngOb/KqKVx
lsbUglh19PeEHQerQAK4bdFAjeS7fb2kwOEoaQ6IBrD9v+6bgLHy9mvrdqYNSnWq
MvFNGcviFCKALHo8Z5NQ48QiHtMZiNJR36mJ1OwQP3u4lrD+PY1x4ry0WTFYaljj
7SYw4mVuPvcPQJqic9pZKZOprh3QTZKMktf0zeQ9IW9p+xoqfZMDd1yMMnL5Iu/g
XL1Df6of6FdTIUNBHfH/b9NSFCFQ6nkrTkcehNTrxZZ9qC9v102MC/Px8nJioibl
cLQ5Rs8DULO8TGFKhVOv1raZqbZUAmXadiIJDJBm6G+VWRZVTZctgiu4FvncejsV
rYlBQw1uSbjJAvfdTNUVxff4iF/7y8ZgcB/cfFMHayAzjiROKpaT3nikxwUuLrKm
M3XYM88WHDZTDvzOWMlQ84RWy91HTwmvfKgenf5nFC7Qy0gbTtr/vKKsXyffCKpL
IGwX3ZqTtAe0wLQk5WKdLwKSw87WND1AZopMkYNaUeTIxHkp2boE9WH3sehWh6V0
FE6T4iRQYGw/F51xWy5zVvLfUWKXCZAA15O1xbyXcjiyZfdpmRl2zsqPPZZ3JH6m
yLqlbCqMA2XOnzy8Hyy9JEP1y3imNd/aux9t7981i5dhZDpzsKwFdlUJ7Id4WnMU
EbFi26AcheniHMh5lws6a3XeuBmXYLSTHvloeFSlFTmQfnEzjMfRgs/wUiIbPort
/MOyWb7HBIAScngImjmmJ7nfUWuXHnNAY02bU2f8HxRRNC+8H3dfJyLc8UkVKQRm
ZrXQkN34m3LVhMZPxTkrRHXSENbVDBJnVMoNekY+HAJy6/GKqqiViDhAwYkhvij5
vTUD/YAHcB0EE0s4xI7tr7tacc2eEt7jd/I6u+ZupHOm6DCKEWnidZy3wvnuJ6xM
n0/41d4iqU4JdEpRxLcZB/Dq4uXk0dYFFC0LP3TES89JfJWUMzRe8xnbInM1ysV3
ejsHpg8DGGHDUIgG4s+lIUcUk5eyifN7Kx1rWRRrWI45ct9+CAWHuiwHfEaBlyPJ
BGnFk99kJqyr4werJBX+gvglpWcwVirUV7XSfMJ4Kr1DIO20p67qFWspC2ELJ0ti
ql5nunDrGpSh73n7LzVylhS3/vmjQcNFrVn8AenGwZ3md0yD+4hU5YNNXWtlk8NN
di92CEps32Rbdkm8hnYgatRtTNRJKYrCVYSUFJpzbXXZGn5SdmH8Nhf1VToHnWSb
y9VPu3wfm4OemMH85p8kCK6eGiED4hRC7e3+UDk0QYv/wY2dQeClbOQAVGVjFebO
NVGF4gf/eKRT1ynru+1+gvFdLrghOkUKA1FIkhGZaVr6zmUoQX7espJ5uZsroPIq
gaT9nPQ9nmxZYBVuEq7fDirLG8EQF/vhIiV1tQxE0DOJ+fMOLnen4MWEwdGc6gA8
Gffk4JomRrjVh4fUkqfYmqbc9wMDTUR16W25aGq+ebkzAfU5E8NCmEK/jJukCtCc
8uPbRc7XbcCKWS9gllTmaEf44RBmxDOneBIwsve1aAGEERNmI3cVY6uT4o3mt0GC
6Qs34N5q43cIPY2TEKFlOwaLqxfhcxxqUT2FBs6OUYFqwBw+AOWLqIrOhN6FiR+v
eqFYbb7//IRxsupjnHyM3lOSASbYeJP94E33XahAeOJ7ieSZezw0R+kT7ovkKu7S
LcDW6cTWPGYbDnBmnwo0wYCEpBN5bzZjqsqSUqMJ9rVsj1exZHX6Xk59gd47Zc9k
6PROLYsa/yzzrjEMN8QFoVI22e7U3IfLjQdIMTorFO0mft3+pZsaFGRUXQ22cBX0
U39QBo9r4fYT5PFODR11gZQ3JwQTYKidH7KX6qA+X3+gMJs2IRXjTjupOenWQwdD
uk8tkqAJURch36s8S8dRQ7Y5IZOsfMAd0SU/Ne6uYrB4bUjkC5aNXDOuBTwToeGI
BUo/cxOGLol9fetac4hOyGRGX9spTyjRCpeQmhRl3z2yPZCof2c6P5IOrIppnqAg
Dm7DFto8d1q6S5fixPsE4MAwkJNO9d7QQLU9WeKKThYC4g3teGu1M1D4W1rYeZDv
K9MF90MofQyThDSQL9GqUxzxdi1dgTP4c9rCZ6VYBGv2Dl1UYjN1ncN4XKJGipIm
e4Q9oKuDHx323eTg0ajrQaaxVa0LKRnzEp07IaQmDbooqOe3GALt1NMifhZ7yjVK
MqTohR2C513U2xUlxQxTI5Eo0VSOtF9vgrwuqaLi3jYa9Id9560KXrQweSOezObz
4OCIAdsNjCAYIeWsTUBaf0LLWglsR5rqIuBP/3uUhekiHUv+efo++aG7wwqHYnXf
uowVKkYw/AdpQjCefbpqYoURR/gI//8EI4+aUpHaLLeJ1wmPvciE3jXE+hGdOqq9
J7xgb5I+iy97lQhrz3lK0wuSkYsGlrvwga96pTkf5bYidiIqGTOrPyQvdqYsNH1D
4FKuMPAj0v3TFR17fcIuWRu02swc35MF6Po+ygRluY14vnKrmqP/XDNVj/Cr2TF+
K1OMHC7OdaX9O65L/XeWiZeK+D0MdooiCGtux4j3w4ruvuYXOCEy9kPVmPBFu3T9
pDxnpGhJ/sBcI22CdqbJucz5CHpEprqpS4GtEMpulQf1tT1wgFNGsrXAuFJ0j256
7jMjiEecAdnkl0uuYa9y/WQ/pp4dzGyvbqBVfT6KPt4VAxdkNwpFIO4j5qKQL2kL
vX1P2B+1VADv1j+NIC/QEXrupW43CicOZP1i1yNcYzTqrbf2SY+UYH/l69cZ3ovT
3odLNftGm6S/HDxgZv2nUvr6QsmmP0Rg46N2/WFTTa+fksMFX7kKHcYKkeMc4m/7
iypklE3Y5wRvUDKYYqWiQoV0PAjno5nE0uutgiRNbP/xiLPzP/eOczEL31WTOD2Q
4vk3DL4vZZa0gp3/fzYXZ4xtQzOa5DAzf1aI36dlaYyptahAKilyRy+unF1QBDa2
6TF4QsUl44F/5MRwUZ9fTKZIQ6hX2YlO55V5hv9c/q9pcsnK/SYoC1POWZzMbple
mud+qxZJJ5mlAAaRYOhub0clXRwXPjbU1KE3AOk1sAZNl/k/xo0XGfS1iY6sj/EX
BTcg9EiQtECGlDIRz2AVD6aryU/S5HK0nurYZthzMhiCEyBH1To24MW3a1R5WTlR
RlH3pPmlLMadoLSaeiNV7291PGI+5Rd1B/sZ9hmp3XCz0rCtdgTCtn/RKNHuYUj2
OkREzfAR53NKaRG3WVAamuJYKzQ7jjHE32HsVstHbyE2r9BqgItpbaArXekyV0bC
R+IaoC+PZloyuRNjJK6yuB+J93DJbOd+k5t0VQzpR3sE1tbf0JRXJ3uj/t0BtEdl
A/zbYZNqE9A5tLxFkrChqvky4ls4TyRlkLaP36FWh7UZR6bj0+xr9EHyFmYTkVqu
vpWyg3IDgV+mlLGrLYTeY3DI9d9/u7kD5tKLBD15P7R2u9whCn9miAm3jkji0mQW
BfOgM9qeFzZa9y+5xEQgQAvlve0x3tu9TeAIpe92EEHleuWTgPZxtlyVdI8EnSxX
jCZXgNNWl+alHk7fCHmAi4fQtt1L2R4wgwmAoYwSy4gVBgGZKXCeVvUMXpdfTlGR
V6pUezBY+kQgqppj/5opqnKvJZviocXK1w9bwzlxeXiz8aCL7fcCVdhl2+NlLs2l
tXAmgRhX71F6tyci2/QdUGkV6rd97PjJgerJi9sRscS9CjMqJEdIMqPp6OsWa9LH
qd9MDkLcM2QCCxfd/wqHOc1JTpXEmc51m79a9vOL3XZchhL5vJu0k8xx2BJZ97K4
PIhLnTY46Vpx+RFM0a6a4kiEQQn0T+eOimtEWCMR5fyfGm/g+I10eRa1SiguJGpO
4rDGyL3uemMQAYRQAVjPm+7f0AdeEIsVvXuUVIFyEk4ZxzmoI7MGTAEQblguoree
X/34GVbolPNGBnEJ1YVbjAyAmjmg9cUUAqR143UBXb+xkc/2IsFTuTcfSdlpt43w
HHJSN/DzDsVK9iTOEHIGwGGMhmm2d1Z/AH8qMae04L5TnkkIl27X1DQU5pNpYuBW
DdqUqtpXExM72gMUJ94wa7N5JsYoOXoEBmMPnro/IsBJBdPH7dPBAvWfe8FKytUw
uQz5VgBa2YwEmajR7c0odxd13rvNZye8nk8RhXodhfLZWD3hAYENP7q/9F24oJ5b
IC5Vnz046TB7kn/O/rz3mrIR6QJGerExdKx/iU+0MyvYT/TOVYBVC5gmMI3X3KVO
gIgGEHgb0WyaUvS07oeVwcfU5mzwUQZkTKdg6aqI4ADQAHu2C4PKgpUGPD9ZLDMv
dNYQUJZ8W7RNCt9aZh8Aja4GPggEXbyGvdJB7D1krbBoKiYYd/qCmyeC8c+eOwxO
KReErNRQUqDkoPlrd2ehtrhcNDtFlj5D0l8ri5T6pKuw0mWUhII+VX/MfwIXCa60
ZsRftCTDNL8QZLomv27/PxnoAvB41QfCJWUDRgTOFlnxy80uQv/W17OERQ7meXG1
Fb/z5V5kgW0gijpd3ygwY2mWSRnWvcJmMgq+GxOSuspPKT6XInRFL/E9//3seByI
O4nLEKoJBa4MUMc97M5booi8flw6vUbpmI1R9X4NRolhG6V+EWkqPBFbD7FVYXgh
50NsYFVPlCLoqhii57ez3Ur9VC3Zb4fRjGnBN5lMWcj6EHGp5XAI+UCC1CpdZr3e
spt+jLuzNlJNmC6KGcn9a/TLsJ0MIG/SLL/2rF7WhS+OwiWL+J5IKENgbjtIpreR
/G6nG7RkyKdCTDMdmZ/cuTeOfJD+cbReSpmxWfwrbCuNSivfeeKe9wpZDZIMMm9s
f7pIyrz7NbxBp4dl7enY1+lX6w8BBisXC7qUGnOnl5AfWriP36fv544lB+0DAKXG
9F26G1DsXENJPRtOsQAOkdEsJ6Dkd15uP7ukkz3zYSrl9ddOuC4fEc8alLooHrXj
X8ZKsC9rbzQYjkaRgJw9VDVzsQmW1TNeIbyW6j13Hpd2Fd68MJyNh8WjIJJLvSHA
x1ARq0l5lin/keIx3KOd6+Qu5ASVBdsDYYgARQPGVLT1KfVCSWhgvZ1k9T5ttvlH
fx15G1cafUrU2EngNRxL8d0/q/kY4P/R1doslKNpMQnIny00VRf2Se0nt85F10V4
qPZGxUlO55yf2l4w3G+NEh3VNBmwdIsjS/qwYaRAG/q3DbTv3Zk4vckeWZXmNE73
7NMx+UcKFrYAOHYjwrh7YNrEOonbqZBb3Po4fwEoIenAQQnxJYfW8rGtVHOY0rUB
eCR3UM6yGAEfiG3CX6aEE1Pw7rCvAtODEKivl0TCClIjkhUlVg8V95akq8cQtCg3
Am+/fmhvMpwL35eVpzLLkgq9CMyEAcyJak675ejpZRyGuzSKG6p4loO/eIOTLzIx
FanqdX22Z41jobHwhcYvRaR4y1iSE1rHRQKpgK3Bnd2bx/HyxktytKmrnWERNTrb
kTf0VvnVJkjHS0MNKkuTGYhY4kIZajcDYz0oTjddW3WTZBffMnlH++OXY2T46sFj
vtaXscmBh4jDrIVS8rX0/8CmB3PMegMje6OgIUgTx0yyUsHKh4yRw6d7OXisVNUD
WZhHc1GTdINONVXIQkFsjQ8ZgkGbyZnZvLjwuZ7ZfSaRDXl70TOkEDsJoPmo9mQh
AIAlFluICDTl0tRFITK45FhyYttNm+L/Fe26IRIMH+Xv+rdYNnT+HNIfTCAC+jbJ
rnseoCbhlvB44kRWBSa4i8OGEZggCUJun+zjmH8RsRwdjJ9+VdwyM1rJbcHcbRCE
q6e9qCgfwUsY4Y2ekOVaZ2tYivyz1LSedL0mrneY5JFO21z0BMO6U2oPVduR5JCx
57zKkR5T8H2hNlCEViLnhT3YSUTusdCTqOWE58BRLRbPey7G6I9VtHVwb+P25GKU
067V6b7nVPAXk//dxqCfssO4q6d2vrThMqfhwNDS3MeYaSPh/DVQshZdXHPP9dC4
IUAvix0nYeMgVyto26Ynz3p8xVcS2qYjJxvAYN5PHQKy562Y5MBrBCpkSEGv0epg
ymhqVVdA0CjcRt7CvyKD4x0Hv1mm/jSsyvSE8K+gsdmu8FCkdwBiWMt7VC/A9JT9
cAKZWSSSelaMvXDISIT+egk52NXeSuFWnirfEGhaM4AuOxwrdPkym4Uf6oRZf8XU
tnNQY2jvx0ivHaynZN5ZwiLPk2JvpEqzltpAFdeANyQ2YzIt3hWhqs1XkEhyYclX
1UqyuK9tLnD9dsIlMhEuQnYw6DCmrQ5mOf8FAF7/zm2HkGO+ws1K7/0SlwZ0m9ac
qYh7VY1G4p/nK9uPp5rY88+C0bX7RP70qXwTPxMraijrmgSeJNGJCG4Q4ktd/LJm
kETQMpbE+CH8YZ+yBNLZLyQU17YCTh8gjY92S7txKVBzh+Hw1EiBCp23igulmjlX
7zFe/WcJIQAbcZ3pcDyzRM/sF2Ue9F3tDKM1V1OaY3F8AcijkUI8EgMNm7Wx/gKL
WiyTQouiXBBENhwGAPoaOEE54xAY35WpOfGuHICb0MQGL/O4/cGVHzo+FXYJOcWw
vkXIyuO1u6rr1r57aAi1UMkr6di45j7wukVrDXAf/mEIDN/FdUDcBqCQcn/nLOSS
a4TexavqvX8HSK7BjylXOxlDOhVpvYPSO89Y2cfi9DnbLdQmfpDuO4HOY+rK79Kh
YUPVNfDkqYZaaqu5U8Yk/Pq3h1QRLGP2eaa+tKtOyhTMVa7MtMxm6jOvHvTrH6bK
8lvOPQm+Yr2cA//vLoG2tcJOSokKPqZjU33cmxWm+C31c7V/GHSs2CpkVvuc1Vep
A2UL6flhuz86miwZZBEhVy4bgxOEzEHZa7YAx9CCF65hZRCTvNfKycSJiTrbFVxE
o+5tP2KXNWLG8ej9388Ih6fUk7VrQRKEvF8qAumJofAVdC5VRXSgLBqf1mk+FRAy
26oz3bLkd8xnZViahxlT3sfi62XlZmgPu9U/99/0KWUnVpZBGSDFdKuA2eWRdLPy
4alIYUHXV2aSY0oGAsQAoTYwIBnO1KPkdy8zg3ItEGLRyJoL4qXABc5VE19WdTgp
7t1m7IyDz/HlqsgQ5DPI5ZsjdX44VvTRp5Tp+KprmCgNGIcjEwJHzdBLoIyMWufS
GOaz8IROaeiDmDlXPK+vfe83NhaTEm2m3YpsGzSAwv8C4siwTkWMpusqAndLOwbJ
jUXvNbxugb3Fpfbd77+43RnwsMPn2zfut6eeEOLQHQRwQxdml+E3Re1B1hhc3/6H
3Y4ypl+q/rioQkTYiH73jW4UopjooAM77cbgYiOsTbbql5CJFUknmnPGj2IzgIIK
lb8ObeEQEAlZcQdq5PKF4XRXltiS6D/sfB00wq/Jkvi6b3N4IHZnagQfJ7ySOZ29
XmXeyRWOQpOZJoMkDBx0E4JL/lEOC0lW6PpflnncgiAZ8RHogbVLkAUnAZYK0GzS
x+O2PDLuxffukqWMha5/p80MfWbJ8KZZpg3eHRccpaKoUb/4S9R/441hMqBkVXBx
UrLA2esC48AX1e29JaCLZySJFa81RR9FxbULx1uPvcpYwr2wPKqm0UriURHt9ZiS
qmzYZLjB0wqsJP+cXAWxr2HKGoyz/fdG2vx44I78h/3DdPCrLLZoSah9eeA/Xmlq
H38hK3JfNYlPjbRmo7vLxJMy+ao3BMH8opOJ3TlinGwgNAV/QLumeKjVlF5QQpZa
FablrU4Vg4S3VmoI3sdJ8dyBAz3rvnztiDYfQh3eqCBPdYSbeaRNlAVaelPIv4sP
qK8/K3g1J9FTGbA/Y0iRMQQMcuhjQnMbdCG1yVDILwFimMm2YCPu/i7Dd6pMVS1M
NIn6Ek5aOp2RMAgoLBcqBiuJB0ElLyq+ea4moXsv7d9au7FsDC6pYS1qOIhph199
b6d2HbCvQ/uBTHnzM2rVVmMI+A1kSSINSLyFKntWIpC5LfGnO9LjsF845gWm/iOM
yCytmWffH0SaLbaigOi1jTG+9AjnM1ludZlyzhmQJN845/lkL7A3/ufFp2AX5Hxc
GSwBHja2KJkBvrHFufd1eHZXiPjSUopevLEu8E52Gjcwl2EymwAh2MhTL0X0BC4Y
xyTdokKInkBuvEYYNSqV0AGcXmEy0JdO7T1GSTf1GkKPK2/dxhv/5S3BagzKoT5W
hgoZymLmTo4+V4Za3hZlIwcBZEoi8uXJHcYZb+gC/vtOwD8pLyLesEVtmdYDnFi+
+dcZFKtSLqRKvRedqMfKi2fhA15VWiffmVZYpbwHpwaJAMxwrwUkC/ElNOeNZj/H
285hbnBTYG97UZwKA+lIE8AdHNssVHFG2dVyEViBU9Bv48fIEeCbuKQVbZWmbsrp
tPtt2jU/4v+yKxUGO2eVobxX9SefHFy9rLf1CITijxBlYatpH1zmNt/n3UDUtzkK
ui2Av0aLnJ1tBCWeyvvENKiI5/IldBbVIfAhVpAJdNhyxi1Eb8E81gH9Q5xTC1VL
STvAsI1W2XEnAeIR+5NCk5r1tJAJ2NVwEZDBiDf+FZwLvGvgc6hBaaaDe/4tRjbq
JkYwCqstJSExsjRJzMbrEH0Qd/IFZOElSjEwDAxr9VwU+mfGTL/B1xve+8ubWrHi
uk8u3LSO6YLw2bmUcYFvQxo8britvJ+P4VPsrAGgPwjAne9yLtWafNmWxa6ANSnn
W8UMh37wihF+i5942mdvquiOvIZWfLDT+oyjrWs5sAoe6GdNQkYEdd1FFGBaahtX
eL7/ko9tX9hKGhWcY11qaKvDGpufZhMmdQKIleyDttMivbMXKuWug8/0k+Ly+pbe
7IVEznGwSGozIE8CeBTUUNARJg3EHQFZSPNuRf+7XO1KbE6x5VyiaiEl4MY3/a0g
MCNYlh9eJIToJAuA2cDpcMEOBjXNXyzhc63TBGtobfBvwbWs8hw0H1Ev4mmAnRkn
eWsOc5uhuASpQYRfWBi9qm3K1+oKA+IALJe4g7SHJyj1dT6oATuiB6g9Dy3R/cjY
4854XhrgxLMqyEEk5V7kiyyjlDLpk02AUCuLfJcNiOt3c0rsurEoizlViG4MPA1q
yTcqwHhyA/lzCmAtu66i2qfLDRbB5fjE1RlGxtGusKUSBsY59WZtUnGHyX9I2cO/
hpFdih8xNCp/lS2ZFkPWqbHWmXhoEvjEZeSwLB1c4wedGGtUJMSE++aDMnyYwY1/
QCNlf+o9tVlrmGKnWxeauLPfgppzWrLWPB5fzcBqdxwvJb+tcclaWQn5zCqCEoZT
CKTWTqkN8E8jV6F55k8UyGgKQIr1cXczUtTdn3a6Ks9/jKOVlhD56MMesbhYKWu+
OZ9mC5SPkM5mdOjgtQgF6M6f9Mokb8F/1Jm4yTs1+mNL8z22tZipN8qKBeuuvPHm
Aa4URPdyuswm370jVASXY9R29lWnioE3scPe84NNX4KlYaAMLhqUlIWsONxkQCfm
s4u/4pY46RNkrYLATcVD9d8r/7lWQx6CRx++LIk2VqS3YdappgQ7TWC3/Yf2u3DC
WMykFxmVi/Lq0HORgsVZqZxaEsnsCGAQi7isUJ/RxWiGzg5SCY3kn41K144es7vm
o+oc+WfBOTnRiiGl606efh/K7NNmROO6ojJo2QPVEnOoA2ThcuUkAuGcHVPZ/FWn
ih9jNcn9RCT2DoDAXtZOpMstuABTvZfF1/+7BE7C7aoJEIaz39gRr+hHFF53Z5lw
suT7C3eafNRvGQ/rRnfXjiJLyyWSKqdFkScDShMXFTxbXrOFYLhdnFJkEDfTo7tS
60EMcyw3YX2R8K7neDB0c50fTleG9auMqnS9xWVgB/ff2SBzX7MKvDCb6c61PwYS
kybJhWm+GKhf8uz+7PUwuV93m1mZP4ZbczGYDL5IFTFSTnrA9WtJj3br++kYFlZ0
kC9RIXdoV3udmu7nyrlIDYCDtGeg+tM81q+aG4G+taIhx+xcQFkKan/useYCD70f
oVhlF0CZciV9O8GEPkw9T7CzRXGot5qZ4DeVXCY76cQ7EwBIJqvrMUKUtjQBU5no
ADaPLEKoFsrP726vu94S1vkJPu03QPDuaN4N+v5qPdEqu9aSu8jRXU0c/rQ7jWpV
AqYuqlLcVsPtXrFA2kHJsVE+oAoQQQ8v7HAwq7XEF9+iWzQrHz3StkokdanFwnLn
eF5koTsA5qfLm7mbrvDRgxIgOWlaiyecQ3N0e91jPBCCJdj4ncZCszTC3b6Y4MTd
DmsoZ0te62mI9K6Fw/yfGs18uSrOJ6EyEUYVHkaxemlVBMq3tL8GNQuZZgbHBN65
lI0oLvY5KY8UP2CwFT9JtHphe3bkzsgKqtRpqBJtLDcvYlZPAqGrSWkcpGcTIdoB
AswaiGawkNMCB0+MnYEgWkgBN8RD0m7NrHIh7Czb637FByO2YFAE+OiX+yBMFTP+
ojP+Ut+2XKOMWe+aVj7fBCbMKaGzTgf9yEnhwB3dGu7IvB/bg6gDiuv+IEgb3zhv
3vEc3AjgiJ3ORu/607H95YbnIyEa5tVOrBR5irkNxIoicvsSLT+3A0/0av/CSYT5
UxnLRkacaaMhn4QCB88JnTqeFBZR+Omk0Rw/496HgP9PAEXmU6Gfi9QfGJealx6J
hPKLXictCC0ySzhajdh/gU1cJdPjP371K3U8BWsixgspfq4fzF7RW+yYOz8mMtvp
XnEj9vMPouwy/9vMNkGcOq92Kwb2WSxVs0wv9fwCzA07IIWGN7vstlUT9fgLxO8g
BZC9/FMPJ69IQ3Elfop84pQHW6Sbg9Xjemf1ec4LAdFcEFnJopummN6TLrCpTJaU
82ToPxThApLIFhiMELmqYP/f89f40PW25etIjKVzRvCtiHs6vpLdTioZLUvrUwDE
WZyaQDXCRZwM17vwxwDKu3HMMs4G/S7zCeWK0JUk8E/bl5efQxkpduAU+CVHe/iW
jU62P3rqgJz4xNPCiCextJ0UX756mbRKe3DrqHWAZaNj9/l4o4Rtz9VWREXBfmZA
D6Ttt4qy8y/myiCPOGNP1xRTokaKp9Er702DzZEYqZIaxwpp5kW1BvWtz/0JQUnv
J+AZxSPyxMQx5c/7veHg0YH6Fn5NuVhwIXMJUOkV3iSshF80RMc1vIbqjjHqmy1t
HE0Wq9ZRVNjIxmJCBUKOtMJ+CGCThwLHYRHKDQfP9kOl+fOjeCDpMkWfWiFabEjL
Hqar62SCNWFOi4izLoLc8rkaHKKfaOBVNmVzXzj9vtw0SKol37TcyMp4v+dqAJ1C
KEdi2hM8VpRYOPeDJl1yDVor93TZKf6hxHoZM0YKe5CrmKWh0GMKN27cMthuDZNb
y++7ISlhSvFjHhPwInsZGLhsirO7lAn0144kBu+mp08D/TCnFg3DpdygFXpyVxvF
AVrrA5TTDqNfbceXMXCSv1Dy9InVHSahFdjlv809Qd/AxqOoL3sBGc7hdg/w59tZ
EesSLlYeEUC8U3OO/OjEMiTcrMhR+3qKWsGvUNXcPDgKMt1DQ6qXylQtYwMVLg3i
JMdiWVLU4TuOH0PVIytL6qZENrdZuq53vGqUb0u2EV8VzZLse2qos3W00AN4pdvt
0GuuqmMaf8hooS7mEFLzlxVgqwQhqCA5DZxUqWN97w4HhhE+LufVn9U6oBO/PUHs
FXCG5KBM43CC63kVvE5QbZWoSZJgt0h913Rwrz179PCeHhKMqikqo+SlaET5shQ/
wCatzg4+/tugKt+q/23Dn+dKB/V2MGEiu9CJQxqr8R++B/bRd0nuhyB/46XqiqEz
dX+e9wwhAvvHHBNBBK2HO4la0T/r2SRDYASkjYf8SUIyQyu74EVhL2EeNvb8aZ67
lsuzj8fc1vKuQ93PIEg16pH+Gdr7pTujWe7ElIHQuZsPc76wp+TDo9cERC6eaS58
ub2tJS1rHuYr8SQDPe7hP4lDKkIv5fLjMbNUeKYMu7FYDcXPdM9iT68bZ1LmmF+Z
BTtem4ZYyZXEvcQmvtdrEb735XLTtWhDvKQl/yzZaVg8Y7ZyDXc5zH5C/y7nEZXk
XLqWj6RJ1fzNSZg+A54MbJk7AW5pePzpovaD982E5PwsquBFObEXDUhS0E113rot
2rdhYAYOxdL+2ZE411O3K5AVnI/VJdeDkFeINME9GwMY5oiBEXAQfQpmtSa2VVNN
kdOjwp78MfMSlnK5Oqs9Fmymk8MbQ49lM64FYAYYS6OtXQF4q3GstBSdW/z/6lum
5vueKMFf3prbK0js2ZGnmNAABamvwnUnvCtBDuD/Rvy1R1GrKIR73D66UXKauSDT
kfP8GplskFx/RL3zJjXMI4q2wfL1Z9r+7MDKhB7PdzTnrA3PYq4i7V90+OLam/OH
ggbPMandCN7Jz2MeKiRIqHP5ASp9z1whkgwAQpePcqAQrVjRZNUji1UH9jCsZN+W
vDFn1lT30WVhcMmtTb6cqvA9yRJAH1UP/JUMieJMpYSfiYc4O1kRTbR/YAQ+I+ep
O9B6aIvRhlBHZoSBM39A6swSEyb5eciNj8MkS1ZYVnB1g+ZFb86BwgeGr8JQSiLs
qxU0B0+eShyskEN17VeztiCNWznm1FxSCn4t42Z2HkHPd3pZOgx5AU94ZhBpUhWm
pplqposfX/HO8TfHBjAekH35EMrnu0U3ER4rOkPVLUO9Z49oDluH5GT0Zyozok43
lr+FS9ZwYRzFDSs783h6aL6OqtYi4R3qWBV/Fph8HbcR2Ggxo9XV28/JF/7sLX3e
7FR+pEezjhA/rMatd0BGWQdP1N5n3A8VUtMbB79COR+NBCxkqWJAnivM6jm6efPR
cYON0mNEHgZvUjcXYk6yhOgCOK7KbEVrNqWrThU3EjN/eLACrmLxDt1PYcjMo7t/
Gi+Nc9Ji3TE76u/CYwoxzzF2bpUQNYoP+pRivbD4fLGGAqoAAMdSdcr02mehr663
9mk57u5ahPznqci/GU6gyw7GWsxFyEhWjLO7ICcu877gJ4FF5yN1gmT0U0W5N8Ul
lGbkmwRKoDpO62ELEby/GlskvQ4mNtyFEcuJIYgl9ZiKiTWGy11vv5fFwwVfJM5C
b2bXU/sklA3PkpS7nYEJOXMjNZTHuH5iLW5WU8C+wLALqbSWf2gdFVlutTNnHrs0
P2icYRVhkONf/tl9QzkbMLbYzUe+EBtA9mARbL6C47efMz6TrBWEQWMNxIQkZ9XQ
c3w7JN039QABaRwgtRJkuGg1VwdV7amyESonFOYruHknvok2OwBoKDNGghEOZbdC
9fvi32N0PAe/wvRKRUa370KFfCu0odJO5db3/ItFcfLPkDl8b891h3R85TB8EMNR
HbrIcdDBKvgy5fts9FzEjQFgshR/Ju5ApW4auiSZKrGlj715eg6JlFRehLOj5wED
1sl8fgW5g35sV5UVJQ2mmIXTX3cK5gFzBmmAiXSlhTkZoDOwbBuYWLwaSKPeqSAS
BRskPyS1+74cjA6n5DTdXFnw7LXWYO9QahT6zk5sUM/8hkqmneSGoz0lG0PQwhSH
tOSsmuS/LsDXODxD2scRNdd5APT75no2I5CH0f5aQVbhnzrEtJXSy1s1XyWKjozH
37LveFz8aMzsquA66XPXzqfFYLVeucpid9SzuTNb5US5L3YhpySW/QX1CoYbNN9N
bLwx5Mq/11d3zvwRTBrIaxi2ax28VwE7nc99ZPDijWRK+VD47s1wpcVe9ly6R8gS
vRw3fkjBQQOZxzPKv1y1pLI/37NNcBOiSkVbQfnMoK3MLUwrd259eeLFxUAHJKJJ
3tM/kILnizLgOCZCdtFNRMci78ydFmascHuVnuRHbLw/m8XCq++B5h8uG4ZmLjbH
OVnsAPyzuL3R2LoUQJhWWHwXvKxS+8Yzffpxm9rjUx1v0I4QVSCXQlz1vpzd9LDr
YbKUkaJuQKqkx+HOi2t7BWvtwNbKG4R2qNdMsLJitF8XVH6ij3EPwHPmI0Aumvgj
PS19mmOLkPOEQL7dCqZ3corshPIzq8Wc+kp86FiK3i/Kc/iKHceNsN9TWZsYSuh+
XOesjt/i2tWIMLyzFxwfJdvzoVyQFG+XTeBQSiemjvkMbwCi5lp5LTI8ri4d+d9w
BVmz9JB+eshXy7hX1Zo0VAxBn7ZWQ9GrphxyvpLnxCy4ZUVPtGOUoS7SPPJOpCqi
+tYE38RZYfdsBBihHXBlIpOUQp/q72WJkSvCIVZFiaPZDHtDk3sXeD7IPmwaEJU5
HB5GSQdIpHgSJW5IyFzWE6KkmRbC/SAri5FM9q8mfWNW/E3NTJOkroxkZ8jS+UYN
MojkFntI0RhnjwAgxnjxmirIyADzlGJKwuefugu+R4tT2saWvBDR7DEMGDkYYpiY
EpD3M8cva9I29fcgs9T/OKZUH5AfSztqYTlq9r+ZcS3XLiFus3McDcgmIfQiX9Nw
XdlfE2HvjvmI1+jEbhuPvdQaV1eG7T/kAeRRmTwf7kJ4fWWx9WtQKj/yUcPWpOem
nIK2IRj2f+gQ1bZ6CjqcpK0ASK/VdYGcrjB7hreZH8uDqvx7/IYZE8rLmsX0Ar1u
eVTw8+4ernLfXgMl6FU33HQ3MCEkfFFGu72kuoVuJwcKen61gLxZ7OBGcnIZTBDH
lh76/FtpV7I5DE4wIyW1P2zkK35Nfwl77MKjvqGIElbF326eEbJiDBR7QLUlolHG
KU0Z9A04OxIddQC3P3AQ5gjrGIKH/PzxYq2ClBOMASfJRxi1Dv9XBhF5FINHuIV+
CEpPXA6Bi7f8MOGzNlyXT4wesTCa5BBV3QRKAk76T32k2S/TEtu/sc1Uj5bAxo9J
IpFOT7YtdUeqwDgTvYIE7TQZFp95E1ElqEFHLjocLWKKoBVX0eeTwdgPtmtj+Fmj
f5U67ZahoyGXhgRtY3csEXI8LSyv6LHmFMxlB7Scz0CFi11eINYkVczQn4x2u0aY
an4FK0gT7RpYJYEsAvA1Lbt9zOKXcsJo0xM97TeRcXE3LqJ4pCDkA1rNgWwxD8oI
O53XpDMTCymbRaGb230nNjXeccqSwI5JOc/2FnjXBDGvcQBzcCb5RmVmndURBIMm
bhdlVacPxC7kgDzd3Bp7S0OMTm/tlIz0KG3Kwe5ByNuv6bq/sbDeEXAz/h7HUXj3
B8g7tzCfYwZH93+mKN8pd7+mGcgQVWzgYbOcC4Mz8XV2u5kksXfb8fNkz4HpvS0q
tzN3XN19nYtCtbVuZASTMxHnoLdPVcwSAf5UtXOrvfX58YoBXaI2ZpTFnk307VdJ
/wWZ1z00pfWKlPfp3u56DdTMZw/qXKa8/devlxdv48J4TXeGpfA3+DnuG24zRyGL
PAriyWncclXRGwIJ8rQ7YfJyUPp3/ZaQJLL6q5xCwbFZOg+MNCbHb1Fapx6YyORD
UY/6nzc73S7a5BxG93aQOJdKTpu99a1AG4WT6vY0yZD27vFMTq7ZE1Q4KVUiss73
RAUhYUerXsHrpL5NxxWr+5JIC3x3KquC+mXwE34qlXKme1uqQeDUQZE5DfOJmKAS
UngWlqxOf0+fEWr8qj1d70SGxcdDZjcGBCLcm+pRU6ExKhYm15yvVF6HX5DgE7TR
wGmga+kEc9DBlsYm++dQLaUKfm/tYwpel1v7056yYo/VJ9T0Qg5k75EDLpKbsSYv
Uu7uiSUA/Z5u1Z2NnmnIOehFLwhUcdma1bG3h5HzqCylEHYLCP9Ex72eJ+n3rBjk
1vFjR9N3rvkhqMM9O28KPfAmAAUwunfHOq7HfNgHMvURgXSh5HQpZd2ZeJhCWedr
XdJvN4LyT3f6exFOwvgsv4Skq7O74nK4rRxa9lvyrEV5CqyEGY+0SqypeMSRNwsQ
70oWF/vPu0LYpIMHteppYAG/hEjWM92QtCA0IMdw4XknqXTEp7skrxnMLNuC2BZV
33yeadvgmjNqxDI+ABq7HQCpNtPu+9t9uU7//Wgv61LpA/YX1CSqVB6J+VwBdNIW
uWUxsrld5rEFVbgrnvzcI6xUhDFm3nL9cHwYU1zlneUsDZ7/bBrcNJA/SsocGHO/
jqewmvwhMXHK5PRSFgOop8PLy8dceFOPZB0on8PQTC9r6j5HZuAwZWRbuT4ABve2
It0zp1wl/t2JpJhfiCsIheNw/h8qaLtSSiVLqzqU7NQw9JAZWSt2jbQcA4emHu57
1wno/9kGs2eUrV231EzOneaUAQ6B+0NUwcHDtJDmHM2snUXKOToBKfaSVyeUoKwJ
3q6dm1q8AIToEoqF0LqYrLSxpa+R3kJlzEifRnhDza87Q4rGcU+CM+H/9Vn587cz
6CYtKIXIs0GriQC9rHesn8RO2/ln/kvo+I9aIODmHLGqxVXLIslR34HGkADanWDO
L6ZTrAnCOR3fFCgyc8lKRwMo+qCFiKqdUDc5g16qY8Smk5bNlithoj77Spa1A0ol
sXdt+frIFC02x4w2scqRqaOCpyXIe0nPXBwq8HnngvPwXgX8fZdsl01d8zelEFPm
sGdDWfEadL6TKiTUujR362LoIoYqUu8JgZmXu4QhYy7F0fhoYAUvuH0xU7CCaQLG
9CnXnSHxzWWW7QYI4eoxkMzFNH8UcutYbB64TvaLEGPrjmg5rkR9bq8aTlaingEm
5owJoHLzcCv2SLe0G6i2riCIb1TxuNdgGAFp2o28vZ2x5i2mZFbG4Retrrmq2X2m
GOJWa+BFl0jHGtT1d7i6mPYWzePDBZoxtpCxepp5iUXgE+nLDeOKMZ7fa07hMeB0
3yU/H7gG8qdvDaIQ+H2R8oL0bFdBhR+yXOyy7ipZkj7hjWQ6kqJcozkdcjyMWgT4
a7B3Bib2Qmsf6ko/H4WywYBg9/V48Pb1B5vo+LodD9MIOsto0g/Fyy3Oi8dCFgMm
XGfj8PwTS9vjhqzqSjGCRt2fIBcs+Rj8WVUp8ffKRauLXc3BVy3zOPwiXD1OuWpx
P+n4L5Tkpfm9lJLcL0BNPiqNuG8Awj0jhXeZH90E41U6jsDWTFhzAOJo66AGR0QX
zleM/tzwRlbh2PsESD6YrA+9+nkJAXQCaxMflwfrM0+voqnbDUke4xCP3dcblTRJ
n3aPtWZfQ76ZTnCLKY7BN2sHs9ie6PfRwLuHgasd4mAVXj+H22WjAlQ8jPsDmlCV
08ypPiBrmXlMGD8UL2oea54YwNo9F6YhKVzcl9ZhHphTiFFpfInH4h8ePBKgW4jv
d3vtvGt+c8MLFwuyKaCHoBZB1VAgCpVawH/1Tz7AmOHemiFdYmGRkxAgdg9/ufdL
btGkB2Y0YKm7TdQrAV2k1V+5QuAaSWfo8lzeuk6uH9pfzxcQ2wHIJ0AIEEo/agOI
McEa55IkBcqKQEfkeg4YhUwWvCpy1XSXHk31krbh51/Rn+iB/6Nl4AujBHgXLKPW
HReashb/bZovPX/8WnlKCLF7GCTr/ezDPYgV9rp+p2gpUu2rr8PJ245GuB64qeOR
dexw1sxRLEqlqB8dK47QAV3vEq4XjeLV09A80RylUM4wCsqi5ZWyzP5et4jQ11dQ
vXgaJDAbemtkIiLYKoHtWWo3Zi89kpXmoSRKQRgdiRu/oUDgciM6INifYzl1PP7/
L5r0t5bxVAXKUMCZ/+7vei/0yM1KunZCg/arrl1S67F2QXib/YuDq4mxF6ueEyV9
DZT7XhLWs3sakix/ymDcTijTEMOrlD05zdbPZTu2SqMQWYP8YwurYqQjapQDJBE2
RvxERltcJYY6htEgiU3Oh7wziGVYZP4HDcj9M0h4XNx2HeDe2dLm64awDYjwHXRb
scIFvOgzpEFBZPP94b57aNElyeKwPrIBATw9h0glmuESAkxaQHOIc7wfU/ae0rbs
cJdVL3i/8kQm38km0rGNV4brEU7dJ8hXVogXDUnudb6oFFzI4+oNNlKPfw/B98Hu
VafvgxlVTmpLmj4opAp/1K1lEvLmA1SZTKu9HUEIZc+3QbIXijtiogSipWSEyvf3
TZ0aCOp72G1JRYV3FSUr3qMFgadCdWERGZ7MUXZp8yGe2UCCAdusHczNma45EMR2
zYckxTu7+ii7bLR1osynXEY2bDCljY0OvxDXlJeOIeJMPjenirZan6bg1/eIG6ZJ
QfNj+iNZs0hjtN4YY4wmUEId9TOJJx3M6uUntllkBEuuVukPS/KY/0LOmHKf+oqO
ZGORjx/jfuLx9DBAnDEWVxgDWfebQiT40cTBDyIuZGhuOpYCqu+NdpbgcFFSvDDv
RsB1KT7Flc8+Pp4rs0kC+Mpqtu+o1ugIMF1s0zj8j+MI7xqPaFoYhMczks1aftOB
FoWyr8SVbDIgX3isnIqSSuxm+zqNVOeD+ySB71GIj72hKOC1rtjjJF7Ag1IkNdSS
JjRB1vJG4s15qvnqKNIib/ZMbtmFsUbuYgg1YTbGUxmx1zEbSFeGjhJ8S55LrDLY
0HkrDtDSlOwMLU4YEdMnOiWsjPWyHu59TeeFN+L8p0N3eFerfx2WqeaN721NQ7cm
opHuCvbF/o8v9yga+hCL1K6oTcg1uKMbuvzxmuXZVEzzIu60TAET+x7UtIZPqqTe
4iwpbXlMY1CJ4LDKPjBQuFb9SOCc8zIwzeOBdgFVqMcsYyf8U8L4oeD+Io+Uc7fD
LSQF1JasAga/BINqY+674v0OnHO0FI8N/uLMJaNwQug6bq+yPjsI0EhSwy717vGh
4QqJ6iIdJR+5X32TtcGRGm7L8dPPwnw4pj8XdHUDXw+hi77vv509eaMuLFOwqXHo
7bjunzcvPZhb85G7KcNclVXcuT2MsYlKJzlwniH3RNhRoBfkHx4C+/QIA0N0tgW+
GGHXDmX4Jq6XvkdZW9UIU6+mBGZQCpN3PFnXVzz8HdVodgxP6Dj5GZ/SqStq4tnf
7S1rqz7P3/o+TEPQlWvktXj5u7YHoJ+gE/Uo0qr1mJhKqPkxXF/5CmOfjkDzkOMe
Mk/QP1Jedg3ICIdXTSRV7KoGIkFGWnhYBA6mHkpIGR66Hx7nKitzogrZOBz/bbyz
vbw2Pk6kX8u/lIxrBp02QjZ2Gle9dh/1gBEetOGxWUDbnv6ccABZrjhGu+nTWiB7
0AJdc1F/iH4XRvadiKjwCjMOO8a0tqT+CP0IxfGDY/EPlkpXhr7Zodd5XxiX8nop
8SILJzurNpjGhYV6z2UJbRQAKphu82Gq4/KHJPUAFrk0Age0Gkh38l6RezUQRic/
6RnW9uRNzMmljbEY1p9dPnAKHN4x1AB+ZHo5PuUhMxTONYKR//1oPswPiozYPEZ6
JLfyHBr0KedpMnG8X8p9V1Mo0uqYCTpCnT1wLoDVOnWMVzXy3xQUEI9mba+/xDM4
dnCEq5lMVKYlCgrHulWDxp1cBdeW4vsHxARP0aIx0P1JNoxkDElu8giLxG5o1dVM
25Jrj/vzKkIpdsKE9FZz9CckoV+MbiPfHxLnpoVjBLxc4VbWa2OWh+W0eHE2Xjk5
eUeXFEdXLYrDGiNDddrb0tfKGc7VbXklhbG4Wnt0iFh4G8XALf+flbw+XOrCMAo4
LE4JV7ZLMqXW34xKfQXAchoPyY74pe8/rhHZg3A3AuP+C5MtCszdW/9XWK5tE0Gu
MC5yO9pyjwe29+NiNN5sgqDwwobkG+1dMBkmi4wmlAC2mehwprjtMxxTkMwI8wsR
8fXJLL96DUGMYnh0b0ei5b7HZgH/ComFu6jzoG+6r9wXT6y8hV+DbNNpdlzINZ68
XvfsCn18RCHTLKMPzpAK0rnz8sYz1hMb2VAU45Vsf/y6e2ZdD3oh32017LjnYZQO
HBoCstNWFn7SniX03ONqmsMinM9oxTGQ7kOu/q5QS1oVF+umhq2RChP+GId4J2NH
yZFMQcWv0rDfscuL89N4RE/GlItta5fLLV9PF919d8OfkmrfvaODoK2v5y8bDUH1
UhBGe21Un0apLXyY4X8bGjWelTCLiFtxtquLlTW9P/UbHk9S4T1uMO9t145NRidV
ClDfWDnMNuBmjyYfH0e10fIs0hRxkXlhpT0S60+NywEhlZXea0AAqV82TLXB7RSH
xqo/UE9D1os0UAEWrUNKvBpusgJaD9P9Pp4+g5rg4l7qFgusjeVmjEupPhDsvEO8
oh81XizQg41MSSgrUk2F2D0ReSusokDhLbKNE3prd1KuAOJxMq4rYL9gNE/VjUvj
b2sHAjpBbY543SS39NEKjfiQjMIKoyNH1AD5Ccwv9NhAVkXIhJ8LFd8m7OOHe1Ff
ayCVxL7pEPDj4UX/SZ+u6vSYtZ2eI+/CqDKBZLwLGOBJAr7HA1SD0nAdY1H/CQ1J
BEoYVR4OstI6AjsLQXCXbvuzWlKX7+HT05eU3F2rHPWh02W0/A9Qspu83hsYx5ef
TWongdarrE/Gb9tWRurUYS8MH26TjZIOTF7By/1LntE5lNS3VYPyJRzJEw3slZGK
/814L1ytlVKyPzPJBECAsNo8+MwFbG90Vi6Q8+4xHsdifySypQH4f8gaorkm4H52
RHbzfT6O0Igq//JBe0rKOyxRPMZRwn/Lz5xG1+3mTrBbfFStRMuKY1pI/Cn8GaB3
a2SjjgGVNxYaBLAHMXFajcz476uL/PLLuayyFbDHzeAhkKZOt+sMcoF1YBc7efA8
NAsykNqTQnXzGY2aCo6m+L7lQtUlKaveFII4fNXYReBAt4DhsMTkhg3pd+VB/4sw
VkGGkPBzQd6l+ICPYYejV73LOcYrSEGAtnR8HMlVuTp16HRxh46EsT+TMQF2omLp
CKr5ewfrpRaORCoBEHi7ga1t120v3tzzRz7RlIqQWfGrCupOizsZ2Kv6BPpkaVAz
/KCQohIzObRLkJpuYm+mTY+bIQl7/qXFBycJK0KIolHDf0tZmH694pq5e+el2fHJ
zCSDeUfS9i6F/lZSoezw4mnoZE79pPGCYsCZeNAxJMhuIkzSIC/QmOpkZTUlsnct
KSt2zO313bv2jDm7hqPmBXfaecFZP1g1vFU5qZbyjDIdEYJhOES2qqki9JwmtpPK
C49WSV4tcsVO0D0nmiyMmOM9ya4A2Hmvr0y3iiyHEj8+IyMqTi99mgcm0kM5sLRd
649tX7wiFFjF+kq+wPjRlmanxZWuXQzb2eBLxr8+jdXntyKaRjuayTdYgBdJYiPb
YH2IDc5E0U/Kra2w2dJuYK1HEN9XzzMx1KKfNh2T+NTi3ZaH7RKYhZHsxg6MOyX4
4jsmk5cQjhVNUMD1sCLFz+JguWQzkc4jKa4tUZ6GEaETuG7XSosrSGIgIw/TJ1lX
ZouhWxtsEsWWLOXzFezDI9l69ROazdgBOlzI7AFKaGoinVt5QTNSeTdLrygop7m0
IYPmGtlN/doq5co4hFZYE2pQcNiTpyruKnH91peB5FaZRSuspizZ9+isP7f1qJXD
0Tzf+F/NqWbIeUMiV/hVTramqDog0e+dJ72pYWyICi7JYA+FNp0rppRoBiZu6hu1
HZl086WcsSqFmDsEtcTTXK4KOYf5jE62BIf4H0HwB0X7dbtPdR4f18pODRc0Nnio
HCR7RbeEsJJ/wb/KuJVgKlHTKFd99ynwgrtD3VxLIExrpsWGn8E2HUKAWqhZxcH3
sCdE5MfTBI/v/DCWFtV8HO40MsV9Bdrd9BTZdspIoUTNQpV/MUaMM6yxQlAQNR9e
rArEGlC8XlCHKv73Dw/r0pLAKllkakypEEbTDdWYs/wHmUy1fT0RipVduGm/e1j3
L8AndzOOSP9z0eu1ahJ1LGLtVMEj6vR2SrLSuTT+DvYcbCYnHic34wkIiBBtqc24
YWn+N6OHQKSkt4LfuKgIb607xawDBHOcGg24wtu3T/5ZNUHcbr+wIl7r+1jCow+r
MNYupPbebPut9csi4R86VoTwVBMOnjkNAse/9mgUiHunuLjEAy/dJrZDpqi6a6IG
cwkYuFm6wd086t1m+W8OuCuTfgN4IpE6WpqpT9EpoJoOMQ5hJ8MXgo7TqxDGpx0L
8KdP9nRtD+d8z9O8iJLIW4iplWRbMaEVFuEBI4Wl+ldfXKcUO/YCnzb5quo0WEwO
nivwPxwcBcP1tIxXQurqPe0Cqp/CttBYxYfNTxcrbn6oPEerzgQXZZxvYP69geau
Uafop7kQ4/iK8C+ln4STHglcZahPFb32O2nsCg0aXeON5yGksZGqmjHjhryFuc/p
YA2ho2gApX9c/4QA35qKxJd0ZX0q30paKFVx0TukiVu2SaSJoECDs0CKvnqhRhQy
BNgy7nZfB9rVUWMVIw6N53JinXpkAUMF7jXDDRWIlehFcHRI2+YD1z1oCyvywk5Q
jJ9uThhnk3v5lUZvsfab8HZT7wfa0oUwTVIe8zd2ysYO9Iy+e8N0gAZe8sTPelHA
/DfDkF+sDqDG38zAwUwdGwMVPsJzIEIT4Ox1G+Wb3930nSWAYg1ulRyTzdWAiZYA
U+j6sCVuOyVBA6aqj9sOp4kNKE219IBMCZQsP3qUcpvokPPHUjnqDzRaONnsCWpe
ARmkq+FQ71UsrCRqoqal7pri5wolFkbbzvY7I3ue3ku7tmPQRyf3qSy+dGyGX79/
oX0xDq0ynyfihCywB/qalvkfcX00KdTsvo8qLnxE2zE+PAGg8mCfGNsKwLu2nbOh
HgGUUMlqZhFe2pVlVUAPgX/p+yaGb0sOAWaKCl4p41tayILB6+lqwE9uP/12KvM5
GAzMqvG0FmD1AzVCNblU2lhUh097buR42aH/0r+JaSz41nLtlmiUE+Q4n0Js/+mE
6HDLI3KZltZbjcxsXTjvLb+RqxAsL74s2aqojZcqRtgFRv7SjsflxhFrhiVnLYvV
YCfSk+8knt0zILOSUvxTCUTvzl/JlInce3ifPJCVwUaImkMClSs+86b5oinlDnF6
PdFboaXnBMA9Dw8G8PslYVSpvifkNH4CYsZlkLC/3PmQ9x5cgRpO/ZUnDiMrnbhe
C0b5YTm5zqsLLEkOnobGClInBPoLUGW/XVGCa2hJnz/aeB5ppIXVanBUghqY/pS+
ENCCXKjspaBDQyDmVz2rZY3bxLUkISVrGiZXC7yslOnlf0xg3INlPKYrKoE0PzDx
67qrV2Kt4NDYrdGAZSewiVLfGgEeBQX8vfKKhrCJEUZ/bRTu/hhKMzRcGBK9r16s
mas1MyAa5TdcAO70WVTWsPsEeaD3w/mt43qaKcD9a1aJ2OwKTYG1K8e0DkiHA6km
OUmp12+f7+n3bOtk6jr+Dc3xkTr4r8n9f1MRWjcG7p88PJX3IdngjGQXnSCXo985
kcZRGPjDajrxTMP7927tNRE4PEz3pAp0gea598oMJRCxLQo65mWE+sSL1HncNhol
qBgi6DXOwGQB9L0bAvA59Jxt1hQt49o7KTZmO3b/HCJNoVGhGiQfeXV72Eeuudz4
5RITgPshcWRNy+09lMr/b9jq7PyakC7Ic7zBqXjfBQCp0TMFDNSaRqBcAKBVeRyb
9QOW1OUD8FCtrcGXTcHDaZnIVv6t7ixYfyE7+5md0kLWPOyJwHJy3QEwb/LTFicp
b9TlJWwqzRM8+P2WDuddM7qpB60c9nzV2e1CvXq0ksf9eZYzz6SmFZh3cvGzMJ7r
F7kn99916eF2uRWOqO7QZ90YpEhXpXCZq3ruT8Om70Y87LIfc3Ejj3AXbCbJBEpW
7lzW47np2O4RKv0uQPbQFT0SJHqw/X43xfEZJzZcg/Us4yftHve635S24Fai+ky6
ArZ8YZtQVEnc609q1UtAWqeVvH2pVuWG++cDyhgNQvsbYbd5W7heIvZYmKmYZ0Ye
/rLAeJBHRLr/rVMkrD5jqpeULwrUPuyGodrD7ToEaoBIgZ7nlVMRws2K/oES8DDw
zBVg9A//AB0FWzHRzsw58ebr14Lvf0opeUBndOtjpN3mMXSpRmigamhmCiChmU/2
diFGpnAvtM+KnoqXABWa5FK/hHeMNldBzwUfngub8YobFOFIORJDFLP/Va2Tt/Jg
zJlEB0/oIv7Wb9KF12iMK8fvj8nulMPiaL/NRvbxmjrIAVPdCelNFoLsyeR0awc+
/QKY4TNlc0NKz/zpMMuAx4HVzwMYdKtCnq2aWLmoNSLGUp9j0485VP7bbsZZcBZH
t1fKOJm8Co0gzWJqvi6tpH98f6rNtM9C7ZJYMyKwlnSsOvnsnbg/TZsrE2hHvfh0
GRY7w5C3CGNTMmZY01jNbNQEuwx4SCLLOv9Fl0+GjwCO0q2X1GSv3Vnk11vfv8tH
wgAKr0hihI0wuL/KxDafAgRXhtw7R2IdXciv2Y8fBfG22N/YhHJnmsJW7Tro64z9
jfmjoPUBJAVglqQ0+esUa6G6a64OEhdj77xZ138/fqGhQZZf18vLFxVBuA8lSSNV
j65W3mGfJCuxZarD3/JsNb/57jL3Sls0FKTj39NqBAjIg0kMB+xYLI2r95gjM9gV
yedYSz4a/TRVjp9/EnuiGN4dtjPGE4G1LDlR2amX1+Aw95VT7y9+LB5xRsASHu8A
azcX1vLCs0kHj4UXkP1+8NJz1eFOJ/Mi6vkkOisRhhaFKtRLZbvs3b1xNpbHTXO3
kVVcyvGGV0LWt2b4sydSPLmusfFoXdyoX1ajoiKjNH9mhTj2IcLf7Hrq0DtYzB0F
hDTZZlguaGoICH0tSfN0LHjugNS4z2BQH/45BUxSNT53W/n9J/BRQB9ek9uov7zj
bJBCRNFESwjOQUf/pu0j8IN9kuLtnVKWdygVJNO1DSgccZtW/bMPXiYIN1M9VLdQ
pFH3JogOVQ55NL9neeZAx+rKXmKQJVrVeZ3CvpR+c8aTwWRl9zZ/FuU5QPauFgaz
ZpYMl3PTIsdRG+V8yO9CEcz6XAwZX5kHoyC2hk4IpeWHMDyJIuGvDKCLPy0MhUnm
lwasGfQwSp+F3C36PhHO1OmrKzcCHUCyx3Zgwv5AiEiccksX2OgmXQpJ3FeRPoPG
ntD5iq9wVzjlpU1xKjxIK3TYeiUad8DMEaZHOUoLOg99XoplpcnDHHfY0BOpO5OK
OHjGxwOrdeWJkeE7d+21UVE+8V/wC+BSMKUDrDtKEX3gL1ebEcQWEIM26/X/4oLy
d9eVplS5y9GeBqtEs2ku80Pfu1nRAl/sWNAYicnmJv+472Q3A10T38uZEw8W2HnS
rY055YqZ07hNvZ8kP3cqKCX5G5kaVAWtEtO4MZLhsCyW1p4kTr6tLZroJMhLU99x
qhpi1ilcSP3uJNq9Lff6gFEL64IEHd+SqOGgXVS7rN3jGI6bL2X46KCLMOqqG+dq
FOnB52InGVU0Z4bPsgxUvmgLG/UnGdAt9eMHKYCaIHdLk5+TonMb2axYUal0ySnv
opQADIMIkJGEjTYZvv8N1fq/3iYjB7MyhNowL8Wk9KeeUCxYtkig5dmnsPFFb/Vm
y7/iIQINBkmITN6Xmg5rzDNW7jSncrM8NimQ/3n5+t5QHYu4bihCpLIlYAj3x2SC
0kT6W01zSCuFoWC09BkIldAZb8MhBOtM5qkQZyos5LmuKisXtZboX64W2x/l30mq
s+i3RNQfLGo3AsyMbSc2dX7tv84XSX/TBdudreD+6KP0WUWFdtDKleRuT3smBpoe
AgrLot8/FEim54MjyatLBGrLdv6GDbaUi0LP6jKOIXhyAyqGKpXZL/wLSdhv812I
4zF8Hy/CRimZTHjZjvTTMYSA7+2OAViNaTsteezo0520W+2KI5kbrBCQFdnz5667
uL8Ys8XnQBzoRzxp0eumay80gXOa3SDDHbx+Hn7I/0fn1z576eFgAxmZIzxGzIR2
OuzHRsruHS/9rRT+Q/dO1fgA5dndZMxGDYzkgAAgYYKKWBlTc7TsYe6khIfRNoX4
dP9ZELY9/flJCV7B0InsDkMqVzt7zH5YF9WHMJ6BfdMfhW5T27qv0Uj4eQSMQ89W
tkyWAymLabc+GaG6roEzj/h8Rh6joD46nAvqXFkvrS5Pu3qnme+vQ2v3kyG6TSMd
6WDcqxzxEJB6dbb2FlNYQgfn/hOfLSX5AZlMs3LAuI8LPZQEhjlSTiVrnK9+y8Wl
VvbuEZI/+xyy/RIVuvlajG956rGNemlF+MD5OQC57DlZfUGcGlkQ0o2N8FroBKBf
gTcl7LmDZJxrQx0CkxqQs+p64PDIsdBrRckJy+52Kwb+HxuXcHdinpPZyQ993ODb
KQWh7YRZStcMIGy/YjVYu171zMhiIQb6z1lFYbJ/weBERHqH+rJCvivbSyYkNz2s
l0kGKMeaOHJxVFFzYHzDM+XTEe687sdJjdAXajosik7zo5dVKoj5mB6cvIA9ycYu
lcKdEILlbyn1wDbhKBJb/QeqSWKuBSbZsuBHXHdYSbKqB1sdIEgoOJL0g4wOg7xq
YaKmTY3LzWq1qWBrNb7Z+YdKYqBmXmS3vFHo4Xx9c1hNAapIM0fnkvINCAJ+TlY4
tkz/LLYIbTPG921FQ24G4M5bp7DFjLzVP6K4Exw5B/8uvngjasaiy19RQQTzSbms
dQqiV0Sv8oQJbLCe+x3ygLQrNU6QctlEqiqmUau5PV3IBsdzFQA7vEMry0mzBmzk
ZS3rZ52rbYG2oGPHHYhU7RTR5FpzdkqSUzlim4yM8pkvG/tl5Lpxco8DCZ/SG27S
h7G33hdXdAygdD7nG2Gxq4WslKJtEeAI2uCBcOi3aWQwNu0t+HU5ntwtpjqOBxmV
xsLtf8J9+QoXbSlK1Ps9DaOWmrukHjJYAFd7KIn0m9VoOn1IdKJfnNa02xo5XFDw
Ij3sKdylbh+7DJ2I9TVHpM3OMDY/8s0FSRB/SJWnv5Kam4R7QrPycWNkklxXWLum
M/EtFuypB8DCA3zdDPgFSMaFiEFFG2hhaD3ABXlYEFcf/b88xYoRI+sfqy7SWsnj
/ZWGQi+Q24Lw21ZNuqeNrXlJn7w3SODQdWrRCtYDRCUrqSIRhWfEicurKATbSHhA
HPbJJhOdYMwo1poxnakxjl1M6U/q9M08GLC1DpmRmAk8d3v3I2zOozwxKlXS1tRb
KTc0zA/Lr+uSKo95mKXFjFZdmc1UZhmMLNYMoyLtVRpdXsTEROhYU1Lwt4r2MQzD
kXTOJidM1QAcyS/FpsA9/IUvPpnPsJ4LiLip1vIOyiCauN7WAghjGyJjbf7Jxvgk
AC0hkRd1mpO9KTApsQvFk9XvNLFtnUZOFfAIhPbc3wHP/mtPi8zJxQL7Z+hKnE1a
9fHx6dLh1Pfz1lrTm4dM4y5wTF/mYkIt1BFet/E4WowuHvNY2LATTGHA5nA40emE
AV3cGm/3c9kQ3fAK3gE0lnVE5iUlNM6Ax3yE0x3YIErnUPmbUo38Mc8ifsUO6wHV
s3euv6wELT+ckkEWYX55/BR5/ZHfpBt/bAD/J9WouZZKzfKkNOHGpXQYsQaaSAxs
Qzr9JmEQWoAYqTb5VfAmWboTfXV2fi1HuCQ+kM/2leQSDagnT0azrnQHk6rTg0g1
IRJ/DY7q3+SwQaDzWdwjsV+VpykLeDnwz2DGb1lo48QnNffiQEN0DY/4FsXMUmtC
NOmNCW6ih/Y0NQ7XZBb+Rt6UkjgFGAiDXM3gEyGsQQ9jLeq4fbZPVJaL63SVcCo/
9qf2wTBxfc9ftAcn+KlJyyESSTkoekGu9wKEEf3nvtv9Tx9WyggehefNIkbwn+jl
6NzUi01b2hAYnD76GnuYoOjirUDFjTU8rgZ/vZd3VtFOrA6neZTE7hRrVJRtXgQA
++wgXATwJJFC6p+RUZZ5D4MeOzSBGGqfB6+svMJN+IjRTR4BwHdnecT4ZAI/YDtu
zPHgd9KGwgvNzxjBzexLtvO81lrs6A0Gnlz3jL8fnEKLYjePVC6PLUwbTeIt7Qwd
Z0IolA3C4ZuEnrBmBCKZTVJSNWSVCSqPdyHEz+Ol6/Oo1+OSHev5Kt+V6d6pD3vk
0vBZTrCBVzrH08jLeqd9gPkr5+R4C0TJmlgYQnx+gEH484R1uTmqAIAmr6Ry0IEi
nRUdLvZgX3kNxjPZp3HRUUdld8SIZIgE4kGQn3i75zarRObwoWHYBk5fgxu4Bwj6
ftizFTWIEV3b79deUVunB2oPrq9oLXuSQdq0QJRQoMxN12vVoLDfYvrnx1+OY0kM
KTGRGv8zWmgr+UBFmmL2OaIjSr2X5FT2cMFJiUvSFNu5Ffr9vcnoi4yvky3wT0KO
ddrhb56EyLojzyjAnVqg6oc+qSAcKgfpnRfNOF6Mkp5syRQ0XPhRAhq/UtTfDO5M
q/PfD+cvyIT2VFvU8IN0a0UnIl3xmReXqsPkv0Svgha7rZ4lmpD3qFuiek7NM+qB
HFvnQA/R4F6DjPewqfJCh9LwnOn5oKyZJzAMZOoO74MHaNaxTXXII9EDZgArYu+L
1b2bwLFpvi5aPsxrRuQT0XKYoD/hVIBx9JKS9s1VX0ThP/cHfm72vD6rAs6Znsl0
LPKc2DWYLrpT7DHqEYZiW7dHdJDPp1JZCiPCQiKbbez2rweoy8zWmhj2eHzuiptc
hEhI6w0M3sq2QsriKH3Nw9z5solJ/MBr+NsjWTX0IJ2KuHLI1ntVdKnoG8T6Q/Eg
xmdfL1cARlqcSmwzfhX4u7ynX88tQ/GZF++H6tTu8vpD/KLUXr40oiYHik/ALRVm
Hy/5SAKPwCSFlswC5NfUvb7CovRWj+kS4AKHworkh+mZz6Qv7P/sx9h6MfeBsjVK
RaxURhGjyRQfX1jCCuYsizxPTKTenRSY5f2US6zeQ+wrcQPz4PFRPv17eLAwCWSY
j/YzqasACyTtgwtGOQnvCrWUgqy7zYDUpVTYXBsumNHYIWGBbDd7k+OHZPYJwY1A
vI/3uYPJ4fiXHjDDPwLTA9DHEvviCVXrVdUZ8/ZMOnjYvgfERQGviRJRRA4p0Ve2
+OIQk/lWXDwBvUJhP9Pnuj2uLfMnXopojtZuj7CJv1d9cQk19ZpAdnVz4eCLIfkc
/SVmwcW1Qu9uJi+wu6UMqwZCAXbm7q0mWYTh+pwMQXd4/DVMSsux4tXbaghqqzpI
p3i1WEhxZLV3xPfwsaHsFynbXHlYP5F2QWUj9CmFc8ghT74h22n598VAIrAKpP+B
DRRiIgDTiK0fkayCON53bS9or3WCDI6tmmJxejt9dgEytaHv7Gps8cAvrJMca2fX
OK/RQbWqGS2GwYiU3Y/qeaVts63tWXLLtZGOiAT4oCDktkPqZhee8WvohNYEjQqs
w9hLaRlOOBcI0+ZtHuXxb02r07vaZJlmoTr+aAJESxhn3VUI/m5YDCozJ4IDQngl
bseJLm87Zb1a6D+hBBKXb5VlJ9ZkQqNQ2IR/OXmUL0xwjA4LOEfw7kEVGNMeurhl
wUYn3Q38YqftjgyWLXAtFqMRNhdSLuO0z2BJXxE2vVqc33qVR09bqFNNgNFk2wbD
IokzCJoyCCPa4/+Aa8Eo7A0t0QaYlsPw8PlJBA2XWL27uiCWwdtAgtO8aT/QR+y5
FkK2RUXZmSL8pQ2r5WGwJDbT8s9ZQdNApeZdjjupOMuLKPlWUkGlxTUCCm8M7jBZ
XxyHR+XqXyYsWMnuAqdrkqIrTxytnACQPLGF4MOkpjxPBNPufl1NPzCujX8Jh+Ob
mWPdde+mLHUfWVDY07ve2buY23MVY5PL3SylnDg9T1Jf7OruimBqqgSIT9jUbOZK
FfzA0uhbI79FcJWaKP37g4EhLChSKmLZ0h8ByofCMdq5XsnrVErLxC0qx97uhl6S
bLm95Ki4pTorYT2+fr7Q2CNnRAPtoH9WBzJyUh4GSLA384BAV01Jyfm2U6K/kA9X
118g5gZFegPenmxyvbmOl9XaTVE0zhMiOfy4fmcxMDioffmnVbQA5g8GeEtBz8Rq
c2qmi+rk25AjbkD0YTYi2oBuLYBvK6QqlzwO8GdA+rv872KJmbeOrjfgAEK8EGla
zA30c/BOebhpkMWJqAYBNGD8I3pTI3+IcR4v6Ek/oJm74t2ECEfJqRB1lxay7kxY
HqDpj+e3O5hOxKNUAE4ywE1ZDD8Q9WkPloIpTn9OUA3tuupIr+f4xB1SnrMPUBVF
1E9ND93n+8WweeIvMfz4LqjdBuBPtGC1Hmk/UOiS3AA/2wpcQhc6up1eOfp7baCZ
dKWY5xFvmSHfCC461tm/rSCq9iIWrHVS2mZCqul6eGR5OSc30mejQ4/tEyAoqS/U
L9Ua74fOsfeV52FYaumznn9sQV/6jfemmyqWzxFV/QUCNCveZYKedrkYzeMglNt2
dFvl0KjloO3aitJW90iO1jlKAv4k8vM2CPN3Y1tIkxV1JHaLb6FJsk9jKln52J4k
UWiFoYvBNzJRw6hrq0Qi7Pez72tQQw/SOehPvx04Oc7bxc+dz++N3gM7623KNjaU
XXvKGRjENbvUC1Tnn6+9nC3eOicsV4rhbkRognNsiSP0ixBTAQNyMMG3dr3kErj9
+SnnQVCMqT6uWcqc0MMvy120/vH/TOxaO4rJVEi/fqCarujIYh7f9X04ko/u1qKy
zqeLOkmTRKkbQwCc2POcoKMJ4Edr+YDM/KphMzXVVIfNm4zavRrpLRXihcje27WY
ZGkFuaSF5n/dsugcUxd+cqWEC2pzyyiw6a5Q2b3m3tSBTAY+kT0mjpCCT0tvrmgp
w46YTf/Dql43cVDv8u/2T5RmzBFqV4FDD7aHDSh54Jgdwpjq+LUuMBsUarP3ARjd
qjhQ9jj5r/Dkd/IGo2YtmwnY4PhSHJMuLaMAkxumxnHHA8wKl1uFtwrxaIz9faiW
djiq0VKScl5RhR8QawZtaS6NIMPvRVxqpGWH4VijDfAQJnohudHRAZSI5iRThDD+
+iOwjEjDaE52HY/yqiS4QO9FauqX2AsD1Z9AcyyrfDDP3jiAmeDjWXYmrcm7aAn1
f4Th0HGGuo17PWpd8WV1P0Ztimrwc6pamFIQaijQGVxc55jaQtYEUjKeA+EoVuWP
/MF1urjQKD+1T/D4yhv00XR85XSLxsHu9thhhKaHWAk7VuNXccr40J/DqvlCmvc2
LZbIHAvt/q3nPdr7qvpnEgdDdBKdiz3flf2577GclMcehF/UVAwRWOg4AfMVHu1a
bX3d8SYIRVOTNIuxhOyKnH5SnPQLst5esbXJfPbZxHvDyIPlt5ylU65+DemQvjlD
OoTChTM89N6MSi3DOLPF8D8WrCvrL7HmL54/wKVF9NiEw9ZsSfYhJj5JCYZ34yxN
wDMZSmB9WgG3V4NIYjs8SMKbrkp29a8iqViPBsCBP1wLmIH/iwfiW7TYx7lIb5tv
eZkoXFndemjNqC9OxynFxX91j6dKzpIfCS3jN/2n2qzxhXLvIYw2/Y5qZBseIV8r
7DoSw7Qxe4edthPzNuzN+1PARPHwSCyWuzHGoS82spgf0EEotZeXxrn2pWF5hQmX
QzMnosoJuHgYddRyKDfoK2sAwGq1NfFb6uzjCnZ/DkUFRh08itynqjnBAZFdG5pX
E2XbBzmskIOP17Hj2qeoHV4obQI/A+JDuVyaoFOcKnkuocj7vLqVXs3Ec8QhNMN+
0K5cfqRpRHjfOCEDGo41vLLrBLntTzKrAEg2XdorvqphNpYUxVw22oSTOPwZOfsq
c4IoTggrh1lQk8uWz93nkA5S37CDSP1o7+C+GJVn6Uh/C6wc4UOybvSFspHwH42c
nux3wwLbBXF+Lc6M7SDPAFB5uIjHdAabqFjYGFL/udGiTLZeX5F1zvhV3R6SOh2C
Kmx9v+vXIqQEqtL3MHYcckhAuywuW7nfnco7V/o+szfjQAu/SILoQarUvGquTn4y
R3iprJKeESxYt+a2iiukrPvxYxZPI+xCicH8l/BIqfgiOjxU/c7PXaXC45nS0kU1
I4l+X/BRTgIJ56ec5RpCSFHxPSMKtzRarcKJJLVC7PRvDQ5hfTpGUmx6cJEG0zDD
VDcS73kFHktlWUW+2r0e4gKTZ7Tj65dkOGZ8RIgb8LXJCT2FyfNd3Ba9sdBkiPii
NUGJve/cfw3Tdjc7/aPUjAcB3QMSICm9pcUMAPXzmWUa6MPDRIVvw9UQzo+CIGSp
awKL8h3JPAyGQReR0+uJa7Z6Rwx2AvyNsTAfAoUKC2AExkXY8V9l6kW8auMoEOua
5lJKLaC69bZjsX6iCXwpqnZsoxZEHJwrJ4mRLYlsZsZpI9b7SILqszFbUY6Or7O/
Dyslr3zV/qnQIaeDi7EoPpQ/Z2A+PZLirfk6uElxUxGrirf5Z/B4CcF7j0NN4XpM
iJ0tOcTjl+2eCFwyXtXdahtWGS04GcWK5Qn9aha+jlZQUeZSEAbgWliB7ZDa/fhT
DEM8twoPoCumvJNe29JiPR7oD+fDhbWbPXU66nDlbkpW6IF0ycMfln3O6rY7dFna
wy89zVeUzA5OuuKrkKo8BkH7AC69rL88LCAzfi/1uDLGC+DkMnUcrittTSTARm/p
G3FoHfUYHCegm6+rFnVmRtM3SABFg/lioZMxHXH/0416QCVobjFghN1YbjwLfrLq
zUlYiOqdtAgnlxGa06KIUGjuJ/RWq2kzHqokYUIAIN1aq8zVHL9AWiV+cfPrkv87
QGCqQpF92ZtrHmTUTKa2GwlBFGJU+zd2mnSIvTnynwHwIsrivxgyTgpsug1BknYf
FrUzJpEKfEsL4fV2NDC4fyIIOq5Ip5FGCCrr/ViEe7+8w3xAOGxxM75zzAcCM9l/
Lv2LOPyNgxPsPdrExeG9gCsuptRFY3pKQ90NfMosBZqsAe6XpC9BaTZBqY7SL37E
+3P074x7ZxVEumbINdSRhBqnkUxfVVR3mmaMxf/GVqxavpm+6GjXUWsGDefk/rAH
hTaAcFBkOj82x5Hl2smVerIRYx8peIPe7rp8dETPP1DE5GPWywk3vyMRUK1Oy4Zv
f9ZkXyFr6wEYpUvf50+XrTIfewQHnmG7wNKcpqEx9Kf6qzqu97q6KnS7LYFCkkIE
+IG0F2KywTkg/zYqmyacM6YCGGHcFd+k16Jq0Pe7wg/Jvo0SxKb3dJ3BhYWmLFTC
iyZJJ7N9t7Fc9OqCgysGL2gWa9pU1sfe8BsuGa62p/5SzegoGVFlNGpO7sE1a0iR
Dd757yPMpG23SkwgjOWdWCeoddUp5AA/q7YhOTuFD1EyPJBvqNSP8NEE9t0ZeoQ+
SKRIl9Ommc8QtxVNdnffa9KuXeiICHp0zp4MPycU6DAfIyOzeUKcbcWDDbh5kqaF
ITYsW6EKslzTWYpwv9W/KCdY2hQPv1PbHWCRbB5mFRqkX5Rv81ElcZPpx9+oGusj
og5moqQYnrDzVEI4wSmxDIIxN5aYl4Zs6RHRALfKHZCtnrrBq+u2hAdR8XYCeJwS
mAMuXlY/ewGa3nd3lHteWMWplNkvKs+u7eD0AJBItzVpr70OIMXuDgVAdfYHnoLi
7GOIxB0qeoCj9eSiMiJlLyhXg4TTXgsuDSO7QJPiv6of6mp+qBxc51fUpNqUVtxB
uoxHjEcQEB5M6f2I4OW8oHeEYcluMl/kS/VKtmyta7GxRZMsac+LfKkE9Wm4lba9
jeoDFthCN+QaIJdC+Dhbiru/uJVL4ZTF/xl8YJ/YsUIh6LujJsZnHwKMa9ImD0w4
9/pBBA5/BYE9srr7UF8tmNhzawcxMzXRWW6we0KD9EG4/FYVB9dtf76CRmFtnSZq
JloqB4D0ixwLtdYhVqWn/jWf4JeFWZOO628qTnIIVZIOLRqZnMGVFQJmErQBLjri
g0W8TB/7m/T5pllsOWLWPjUk7M6pNbsa36WXHcFs0YHPjxaIRfknBxylDZYwSRJm
cOAvYVsi4sUOpIJYWzThTrA4FJgzX51KKdYVPq1a2NRa2VWhUm8IVYxXDinliSQA
0nqdffGfwi0iU8VobX/v/WmZumiRStynbcN/UTAUaVvz0LgLI0jmTdprDps4Axr+
LqF8rukKoo1SfMKlQNcUByK85rcE3OfJffPSXnKTSBAZ0LmHbT76wG3okOxbbqQ/
nvq0yZEPzLzCj/OP+LnsGi5NsjJVMLvxDRKOXUyXw9BqCvQpXBJ8nMsko+6VRuCA
6b3bwp1sKnYTnzibvmRaA6qpHcVjG8f6TDdlMcC3Dyo2HMEE6xrYbiu+0v6Jgzul
cnWwX7+DYLRwxT7qDvEZ5qYMHk1l5RwEuu5cgp1DeFj8LkmKYBjKt2ddfqZ35FUb
LLchCyAoD3/JEBG64U9bvyvFd+p42Vsi7b6PIlDkB6p0nENa36kRRWDWEWjJFoox
tY1b6VdRM5YGlqcyrx9hK2iWf54u469dtVcGLAi+DDEkpzZrlUdVLVlAg2OS9Ma8
XT+Lttz9YfkF4oWbJCnpnHJTQIBZ1pG6gp9xxXkU5qrtRFPr4oR6l87jYYEePed5
n3M8oA4hreLMyMpgKlL0+V59xHmwMaJdKOeuqkmU/YTYTw6HhhyRh303B6/Jc1N4
5xQ26j8CtiRziG13UHldA8h4G+h0y9uMpswbv4qROiACGhflCP8cty7ev+Fp/Gyi
WFsQV0wRWVLU8cU/4C6mF74PhpO7mkXy8v4hY9VWZr1gx+7k43ziRMRhNYGrq+d5
rWT2lIroE4URQ4QllWE+OiVTgz6S6OB6Z4aX4/yHPzylYelGJdxbh6GniD7DBaRB
pIBAXncW73XsfbgCvzlpxd2wbC90fRZj69PiPA4WffLEDYj1r1o1cWW9xvARO+MR
iny+7+6LMSQmcCIPUhAw3bJ91vaIHhFm5Lz0GmoJstMbXdpCd36WfL5dh3tLCGNb
U6UZNjnWTyzdYWJKbIBfONp2ZZ57SgEHSAqpNcsGwEX0kLLCItAqV9af9GkcrVVs
AQq6IJS2GZ7BIoicuD4/KCVAd50iLkicxVVNKrQOeGe/VuPpe1QRE/efR0UBoz05
jtMBDuk/2AUZq44WvQ6I/h5kTanOvgDMmPsNluSL7WdGS50Hi++EzNz05OJpGeFH
9xpS8jaZ4e2az4/yJmcu2+JB+2KVQGmuxzevjv1sgx1DbnyxaoROzYaiCbg9j8jt
PbvO4bLUTfLHYOeKQY2ms3Dsupvbfu1h3qU/H5tF0LpijLeFrDNch3C6G3gMXy+r
bifmS5e4AGrn6DsnEEbLai8mm2jslzD9XzD9XmQrVpy8VJbLSFFwYhWxNyVTb7bM
mw89SjsqI2psKG8PGl4STYrAafZZV0ay4uXL6tCLK1jjnOxlkdiTFxLvz6xePPJX
cnqgH7Qv5obakEBacFmRUcQx3hOcxTqOWIu/sv5LMSLc1C1UYg2V71kVpkhCB71e
k9yQTpRnX+V3ZtMpfdOdB/LoSuHz+uyrXhKi9o1tQvH9we8BOH7udOooyRuIe8Dh
0Um3DdFwKytlr2pHsBS2d2jstKki5Fv0sQl9jWuA9KxT3+LZWkwSaL+m65NhMIhv
R3kmmg2C0P8XU0LZ7SYtkBnQLVlkhPMiNH7Sxbfbq50Gj7Kg4ut8o4JWl7dNeR2r
hS46Bvro7y/Ya0orNKHVdlou0s4FV6tedfokIRI4KXtbKlz+zk6r0iLP7/w85pud
n5/FdE4DzQoAnM7Q0OlZ6DLfDcL7cJtPaA8ZkWvQ8/l4prHC9jYDecd0eM1wvQ29
iHtz5gTWNObHxvctscid/WRwNMeD9AV0vvFa/DEOl1V6Dx7gZC9jU3ae5q9D2lUN
fOwNur5ebgBxaZJfRMM8JvyeGRMfzw9oiR/ZOVqwM0RV4TuPYY+czwmS4hbUSP8y
h+/MRXvwgNUWGyHVKvlsOuUPVu7gCa0+KVHGo38S+JgDh7FFZHdpv3e4wTRydePS
UlbOrDDrrQUKarLE+ERb3RPEFvbvQRx1F+kCmfP09lZqDBmtqLS3us18s2RHj1vO
XXsZnjjD1x/YuK4lsGR2bk/xK8jC1WpaOvlKoiI74TQe1DG2Vc6XWlINs8AZuoqY
ZNCAY1Gl8yCiPsJgc0W/RwrpCY2jPNHraYrCVunjvb6E3qMoRAzgPkrGyDNWs5hL
ClcLYp9GhnUOMx7JX1h3wlcw4doJuiKi2i1m6Yxa1eod0ofreJsRrYer0HaQrA3M
q7KlRDY8esvHLZ7MrBLjbdLs9xfBo1XthKCXqok7s9eS3qfD7VJh88RJjenqIKvs
lwEIOIG3nKgC1O7MnMCGr8EFvnPPUdaA2w+36D0s9qhQd8CvWp+Afa9hcdYiNR6T
iLlv9VZjXZDrdNJhBqtNoAwfkuYgD8Umdbyq/47yNxIOZN1ZGKR7ffilXoipnSKb
8/azRFJJamjVAga1Aw+1LSzwd8jRhWQgP3Ip7CkUysmzWCy+kqU+kwY7G33IpLqb
4vI79gaPPdpsjmCFW4NobfulA9lpcqFAhuvQ8ThR49H3enn5egXwVIch4SpDA0+r
aozSftRFPrIsGWkYJiQj2Ylgx/0wz+sRJjulWt95D8pa+3YBbT7ZFSwqnnm4mR+f
kfZvXU4hWfysaoAnwxqbxaJiOj/CXAf1IpB3OLleVs0Ikreknoro9QlcBWUEfqs5
s40CGXa0JsJFjjv/kKqnMmsr5kXovAlIRJRxjp4827STkMWTap5ikI0pNLtTj1cr
Zy/aorfpkZGkoDBzXRDmimRRRgtMFqblUDm/0gZp29o=
`pragma protect end_protected

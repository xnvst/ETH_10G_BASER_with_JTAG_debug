// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:32 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dws9l5275r9ktqTPxA5uwbT1qbKANPmI9yG4hV0kneYykpTOIbhRmKVAVGX0/1qh
ws7Zl92kTmhq4Vc0rpWHv7rqyfK4NGE7L50kpz0S6rwUnS6ejH+iYPSjccGwASRB
3YHDK37eZF8wfm2x+AuZmXGfDNDxpegX94599XVkTks=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4928)
okusHE10HLGsP5YABWoRme2aT1SCYPw7N8D8uUz7yK+YUpNzK5qDZSFS9/MBeKtF
YR9YHbEPIjxzDnqJw8SGj7cYobohG1FpbijDPZTZFoYmE9DfUJzlSg6+P4aQ5Xz9
WwGClAbmwN9j7KkA1rr7naF0M8PbIt8PJWhI5xzTLJ+ianzftwN4/HCLewBlzOl+
rikFH8+mue77CnXnCs8HHShv+yZYCUw+7R5XpqVm8pcdLgYvsYQ/MfHpdKgLpwur
Ik/ZGsrd+p+vEf5obTg9m8AB/wFLFWDjc38w75pxPNHYiWaNKRETbx3j5nifsC6m
Wm8H+nK45AppSvKJ9I5oGqTlphhfHuv1gXza+Venxc43MmYVlZli9V/GPBsHlW4Z
hQY9OV7ZrWqRZ2sZEbBLCurIgUfKmFU05G9vWPm8tMzmhBjYEyD94NgkD3bCeSNm
GmE2xMgL0xplbdQ/Fw5CBcsw++S56TJk7bhqr/DgED2rpr0Bhz1KUBL1eaTyjZX1
0WX+L4vkp9lcm0I5N9cp206USEXE1GaVmcqo1+TpBp6AEqDhaWq7p09nt4BiaRzG
F6FU+ARhG2sQTeDmWsks0bT6y6TftpRRdQM2z0Sq9fcTiA8XAup6LFHwTaIrTOGt
d2mQbX1KvvTei+LBqk/wvLi5wiwxWG8rs2XYwwf5K1vWAYr6y7igN+5axKvOL2XE
GtwUlwyozBR2Fftk3E+PzIOmhcupqDsShGe1WxWzjf4CWVS4cR2rjwq6paMLwY72
tmcEzWZ1h5MwNCvxBYTP6AcSUq/otGngHxrPEmaDeppEF4ihSAu5MTYwOVSTQkMd
zlOkjhAEfJKr08K85iqKqLeMSc9QQqOBR7bVFWXC65Xo1ncT66dlNhh7gO3K/OjU
KGcph11S/PSRzoGSRrzeN3KEZKyThIDIclVmvnkzHR1yLo2s4cajYbop58tUG6y2
W2BVEcT5tvK8zkumevTOQKmQt3h+zkXK5xIBKxvpuP+Rc6sQ+jdLzNjsIw8/eYiM
vpF65vn+dr7xQR5Cw3KLbWyvGQJeuNdP5ou28GSp0r+Itm9orMpz8cp2t5u/PFvS
iya65SsUe6rpOywc5uRTX8T4CWMdv6HREWXeiq27h6rmx8WHSRDfAIoKwK33UZV7
FVYSyD39zDCN6tYlOXhwu93dGBQJQVjCQR3tcBizHZD1KYFhZRf9pjnMsQmE9J3H
X3rMip/6allLpwEqIR72k8uxbpS3+sHfBxRsBYv5AX9WH4t2SWz5Txs2HhUTMNAU
1Go/KlhtF+i0frzWxwK1YOcsukrFleFrXb7r7cQ+YKvETjTjWFrM6b1xjZjwymCR
zrcO5P/FByOUiFPHlLJdKwyguAOriXWisErpWdvxpa3zt7gYkz8oapajjvjcm61e
SVqrVBU2Ot+baX0TVc8swkE5WCE43uDkgBvFEyhN5mdTHbci3V24vyjs12ar1n9A
8ggJ83BTo1c/DdkE3JX8IJBMj4UaX4jaEqqIpJA1ycWrQLqszvFKbVh7bV8GsIW4
V5X9Qf1fxp2LGqAOqKfiA1qHQmmJDnmfd6JOLcQ0Qo9ZaZ81F6R6M/R8upZ84dCI
EOMe+bhb4BZiLTcR+sxWXiqDA0YxCczrcG6p2lpN/6TkHkoqFxB1l8TKj91mUSsU
deYQWqjoA8u28I0HXNkPNaMtPbN0QD2NfiKcrkynUuFAMNvEIRM1xdU0v7BflgwJ
UwbAHfbkxYQNBPsJuLHa/IPbWmRtIC8aQekqYG2PGtj7zVpsXwVPWLiQuRhSNh96
AQar5Hg7h8HGCJSkEDJHIMmAukBRMrRH2VE10ZTIkzXyRlg6aosh2fQBrsAhnZZo
IT3/qFzF8yZpODXKl/QrVCc4pczfRRvj3J6e3tT1nDZrE5ipsI5jUuZCk/toyKy8
gplCciLLgohxJtBdDyitXrvUDdVkbjlTIf04c3Gevv6rO2KXegl862aVxicVYbss
S6c91RVqJq6ToQfkkdvBH6k1O14F4tZAP1hixRyinJpAV3g33QXLvZZOz8degB5Y
5OWkM1w/HRARSBPblIiEdtfI6/algJ3qa+4kgmLGeZlTQEk/1traV/QPlrhZ2xkw
zDRAtL9e8Mgp3N5iTGld6593ts6fGkBGufMMpKFPWt+TwVnFJeOU37MrYl5NT1ug
oERz016oMYfoNV33Bk9iSGe/stJamjHwmoWyNsZIyXUg20gRa3u6uk9AQpytkjlJ
3rsQPhZ4I6fGvEvnRe40d1U19fJG3r+ytMofrs9OBOmSVXCuM8zD4E3lwsOCFFE9
5s3GVYWdsgVUWvSKK407hCWYOfd2xNR+wJWuOzJlHbFuTwNGeMscx3z2z8nTYsb4
EWyYy2wiurDT1JCMYWQxmk+OsqqbWfp9ELMD+BRgOplq2/MArDkQWpktDNcjoGtL
2WSltMUfWl9rxRARmfZCXjko0iLoXtF6+ZA1Phb2SJI/USOYG45tR98xcM4H7bOr
6SgFSmEvJrGfrOguEpkR6PriN+ODDPyCH2yBHVU8DDvnEJi8KIgjR7rAdaG5Q8M3
BkA8OtiHP/Z7iM900sy1Np5ci9htPU9KOcN2FAxbvv/I+Cdc6XlEF/4Gu0GpAE+V
goKp1lmmVKfY/9S6BNVJReGeINvWOUdQPtiaoO9QLRVpkKo1j3MVlqd6ywnWfrYV
BStzBpB0XgnCHkTP16594YPai4hppJ31EX1UXbl7CQhCD3bFuhvhHd890sBLuh9C
uVy06rVlq8cHI5vnnDKDT8mSXiXWpQCW14OgnYMYqWLh31dI3kxSJGToswWi3NtN
6rKKJZKzKDQcNO/j1t5gnCC3YEDdry4+VWRZ5L9eTOcIUJgc/uMey/G0fgMaFwWs
bfZyrwwNrD154IKeD9RiAkUIBodJ/XdB+Kne5wFDO019S3BMKcmzwx2figYdZyZy
hIHwei/Ik55CsjmHE/i5jIHKBUh8NSqq0r7HF3CSTP4zTAhkgKbUqZhsDWCBnsld
dwRrRpsFu7Bqycp2q+YE6LKqpWktYBGKFA+o4QqVEfwKtOihbavlUwBRaRZosfSL
TWgWNUfUG6ZaFpV0BKcWnIH494Gq2dI+aoMeXfA7mdn/MrPTmcekwkJET40TrSK/
8erU/i14En2Wv7i5a9sRMuBG3hW4SWbm9ANSnEKGw+kUu/tUrrI/wN5YjcrmXsfU
MehLRbVYRbRPwQ2puRaDg/li+MKzLl67pqIqF5r7HnHxi2JUBgOSojuS97oy1daA
lPYHkg1PdDPd6E21sbszEdmXimcmXlTXv/FKXuPlNwwfOa+g1ng0nMpdY7lkA33P
Zs2TH6vrd+9mSWZwf3Gfma391Jki2BlYF01Ssv45oAVZ87kZCE5z3TjGGiP2KujT
GQzDPiBJOZjeqQSlgz4Gt2jg3SFQPuT0UjdSh72OVgdghJOran0xF3VTqkRrWpTr
KyKARtHFW9Gy4QIp4jXpawqhb9b8mwjdOgvZxO2fRKYaTmUoM91JJ6rGh8F6LQnl
Eh++K0tpRYWG7809clqvgfVdGA5MvNHOrCY7gV5bhlMZvEuRneGTIZ2yYhnfUy1V
VbERYHaPRBHcizliERz8ym4vjwB8m4EM8qnRWuxefPmypNvlSAti/kzQvENXcJPZ
Er34XbcvNvLLzAnijtwZtSFoNtn+5vCqIdcsMDLgpoJvd8edEGQXGbgqu4+M7FZL
BISfA3RlOZEzSgquh13TEy/cPn7SC0KrYm+6z6aXKGNRajNkNPrgMdnHiynmVokf
X2czH9l2u2N1cj5YUhrrHa0Hx9TDsNIajsXQo3WdPIGSaXUKd1WnjKkwSnhMJ0/6
wbbX6pgQjxSWO9j4ucx8kEYeUqbmbnzFjqUiB1t1IaR8wsnkOziFpzASjSj3fE4A
83uJh0AfGpdUzyEkeRP0U+tS8me2fJ33NqbEe8natIrV1n6mAvC8XNrtjx5Yz9Y1
rMbHcrtIYCwUS3Y5lNuwJ1s8ZskVb6jMYAaA0xyPPllA76kmPsuBZ8mjxfk9sL+N
FNEV1lzttusvvnRcwGrEj84r6Z/3SlySNHsAkIrT6vMkAFr7C+xQAI/oH8YuB6hb
jYDSU4DO4m3k3NCXfWYgejatY6F1NYpfs42iy+BZT62hvXby0f4nxizT+Ug6KDot
3URu4xstAbRTH8QQ8Z7rbhNFDFTPSbNZi3sBQ0ZIEE2W5wfxPp1JNnGYu48+6hjp
ksA+tmAk7Z9DfKptvz7JO9BYnj8d+WCYzYvI4OBoFzEhggPKIJ4cxcepCCSMJmrk
K9GcKHFF9iGM8aWRYABtUlsJrNzFErLvyLXRqOC2qP4mHBMzj8+dmTO+Dz7tZKB1
zp0PMNb2+wm/tUDs1PuPtNB9DhnMTDy8nsT4tckJ2gIUiX4Zo9mBpuJDv6QwUm+5
X0JFGv5vw28rDYRtmGcv5VkcBmlZV8LrcXf6Fnyk5PPRTA8QuTRTzwfCQ4KbdvR8
XRkdMiPQzWdH8DYaNvKxOrr4LsC6gjZnVmi4/cFdamwGBiEcX6yK7/DGKyVFW9Ld
hYvTWAiNnW4NIkBS5VM3lWs09pH5BkViVmD5PzZx3lbFflr7ApfGefFVSIkE306S
Evzpn6SNE97E5AeQwDjnntHLXepfDUdKBxDrnEsXwhTruyc5ksxn+SmCGs2LlGlP
2LFOAKZyIycMHrrVMWFRHlmlf+AF8OQaoJCT55CTjVxnuGZQSIOD5CgvX/rmiSJg
0ka9jhdJN9BEWYpXKMoBIVhlqmd9Ow2tdW9KyAjlOSZiHK/leLSynG9u/XcfE5tP
TOTAaV8ZanTFa4jaIP65H5Y5Lz2H/d7k29eP0oUDCIkgTy5bJHic3gyZaWCajTy6
iXS4JsBmyoqkLFL/+hfJ/KxpsLfPLtg8HIwlbd7ucbLniYEhcfKhmqDmZ5KEVXWT
Wc6TXBQ6Ee3Oa1DKSJX5A+LJU0tGC6H0zfC5NKs7UlV83OgZl8vUcTF+0KHRsPT5
n1pP86vQH3ZixboPvF1mpbSaDSEFHdCBvv3dO9WejAUx1b5rmSj/fvSB1PXINMre
9j5U7cPari232FyKIDBaIk0nZgXkcXSBC40ZJu1ALB1EEmpehMfUMmwmD3vnzztQ
r4vnFVAZ8bkRleLaJIypgZ3Z+jlUl/KBAvpB9ICD7e4X3dmOtNLcFV+nXqpK0MF2
Pj2FlAiJbTXUUxFDV0N38Or5cMcEiB7zTpMxt5fKPpSCTr1pjmM1Wm+vbMItxtT2
9ODsqV3imy6nn7whpPv/KTelyVMOQutbw9237WjAmfKViXAATQ850IfNlI0BAHli
LlYecvhvLIdk5ufjSt3Do0ErFoe1HtYkNNcYebjGveBNteAvoZViGjExE8IMGdCz
iBo9y9F1RDOG4lT3OqbXfNSC49f2q1Tmg44GR1UbpB7je13tQHPLyvavn5/LVtyz
Qqf4q6g10UPQSMdS6shGdh2/6dIYbmP60FZOnb8VTlk/jzvdL4qd4B6R71s5OWe2
Iges6HyljRrIPmx+8BZSZsqr+8R0IK4D4K2sYGqAO8PYEbKjYvhSFqPdeEkdt+Jt
VCXRDwVKMgbWAh7Lz1DSgeY+S88wOfGuapDFpJInlFThPTMJc5bjtPVHauFfUF8o
cmjeilCdSEyxusVif6okYxtgyI1Qid2/tbcwGEfAIlucNK9B/ghFSyyUBMtZxKy6
MU/GKxRGOCBkXM3Z7/9vAtWPqC3SpO9YbXABd2RxYrX4P7XM1TIM6g1+yGkAcycL
NzTO3o+fSzak2Gssn7jfNk767vyeNVJLgA5dn9v/d/3h80g09P9JWdCIHM8SpJxF
ipRarQKFBhLRKe7gAv9X6/eoWWHkrjYPrS06Pzgr78MYL2W6GF7q0WaPqhPk2ai2
4pPBrfw807C2o9QLgnnRNoX6mnfnTcvCsc9hWlagYCysgQJLyyjOJFHhY1wqVj5J
MwRvPlaI4/E7tqHe67DVmsWKivYojVbk9F14g6Q0qHuF3BvUOyjWyq5Cnd0ynlhp
4+RauY7kcts5xZNHekJkpBjUJ8Ta0KfAfCqZtRrAfppQDlvYFf7iRK32V88q7oxU
1wZh9swtwYMWWhi8yZR5Jc8gqHeomYCyZM8ZEjiAzrpbwhDIvcLwpabN4JfqUVVY
Us9tk5blGKZ/q1v8KBRIpFKJqeeQKm21zZz56W3vT0JeDyQc6zTPWQjSNQlnpeGY
cHFpVYpvpbpUSn5jzkyo34uJb+SA5rXpKKihXJ2ZzHxf88edYqk4uqWQZJU/Dzso
0npIOJjXg0xY6IQVlBfd6Ct4D/v8Sl47dfwxC2/TPn53G3gxw+q0TJvvKLwSe/BL
Ctm3mp9bcHR7seY2zwyrlakwj09jrERjzioXVK9lnZmyhqefGnBsg9g/ITsLkPq/
m2UN8gC/mClDF494ljVdq5uWFUpAGJlTD8C2NBCTwVmiwYZDkP+qB9Vrg7hAgw0I
ud06OwgwbChkRs441G8rOre92offOO3aaXFy5TiRj0SKsb1eniOvj/mD6cnGup3m
Iy2lUheyh6paBzY84kkR1Rpcn+PRIffFhUeaOY5+f7c=
`pragma protect end_protected

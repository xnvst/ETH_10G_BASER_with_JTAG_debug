// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:30 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jLMgsrmCS7xGNNm+rPU1SxoOgty3I5/tKVitLfqWmtu/9uWcCt0wfuV3snS9KqMT
tWIZldau/oO3euEeY5t/WV4ztIiPUiQms6zxRFF+y6yoZ6tdDviXDz7MZwHosG+V
yX949A9NTfRGPRmmY5UIXoPxxk4s5jhvIr66Nhx4BIk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57888)
LUolncKYxU416fAB4VIjjnSIro3mgylNnYEmiRXixTIqsC5ZtxlvxkEKn9K8sl+j
9hySnIcmvqB3loEyv5QMPEFBpIjjz+m2xNU1f7XGwhxB0swUh73HHJCpQeFrftrH
Wf/Icy3q//6l8fUsmMo+fHzcvhkGslcbCk82ayJIj3br2QUds08OzboAhAQu5Ste
yhUHQfxJqsT9MbvXabs741d/lGMUwAkBYHSEoIxW++bxR5P8ua6kZs5FeYYeQeK6
HfqXjkOdMoH/ol9V+yFsZXEa+Fv1pSSRYrsprWbV5zpyKIREs7Xl281/3NJAl/eb
bSYgN2HkHYLXNaOOX727RmxF8tXs+NcZyZxfdvcIOiDlaw2o/OrfFZ6gz/TVZvCh
GpfDCfTfark7E9AjxTjNICGzcP4LueWBoGfR51ke/Q/kR9jtpPZTTUxXRHN4PyqH
SPLOKb9JLsb99zXbmXiWKZkFCrGyZA+nMduXRCuxZGtTHu7Mby7MJCxipcNJ2GAn
99Vn06ww/dij+hUEf3Xm/scMJeuXEj42TMNffcJ3ObkxauBg4u/Z0JOaOv8peufV
BwCSC+vflNEM++AGdezIEs5G9671EbYq3i6HQVWamxnzxj8x/7WfKN2b7fhSCNI9
WzMoHdv5utyYLytZbz3cqJpPvHGuTrqTjgmo6F13ZNRlYxwuCt7l7b3omSraLu06
6nQ7lcou9AEoJlDl2E0JHM3KeR4w6iWKCJtMKD9H9gId6nMe0+pUKWYE8MVUYODD
WuKzFyz6cMnoXIV14p50ZUXLBYNAFPPSwH3a+/UBXxiqvVH3OZd7O4ADqvcffcRX
5zOR259ViDA8dlvxRKvlQQ6IqtYNqxvyGCxtYCxKEIUidgJpvcBHOExSAdo0NwWl
h+CyRaY1CJxgQrW0hhBbRhLPBHywW41MGo5GP5QXDN1fKy+oc3tgZbFPXaRY0Spi
s7eOpBdI8lm9UxtxfMLBm6TRHlukd3J/G/o0unLV80KgeF94/AZW5m4Cieei6tre
RwaGpr2t8Zvh2HpqXqK7a+vi4SuuyAMpWZQej43N8uIVdAu2CFkP+5I3xYezWNgM
MuavJCNvCfm6x8UOpBDnzO03gUiYG0JrYoDi7TZi/mu8UcddJaZpwZ7QUH970HsX
s1dtovA58+FNpon45GL0xQ62eQ6poDYW2cxOlxcf50N+9r4WfVdkH3vz8t0GGiY+
cq6MV5/FW3E1azthiRAo/YJ3rsw4SNH4uNMayVwgOLJSsfk1iUyQnh0qnIdoLFSG
Cb0rEGGn54+skHmDpyMvnD7yr04KWHT2D1oCZH6+ursj1jIz9+NHAN0TA1V4YT5a
nEjAS3YarryNUpnSqA0U2yKY/fOEfhW7obe3zzRwZ5fwSAeudg79kNDNG6GUvTcu
6hjizb0VlLUoKGJYCV8iOspE/IXHAU3xw3ln9tCzgHTPYCU9Bb2RkuPL0eMw2zfu
paWOhZijsvTbbdiOFHTedX20U+/wBt/4iglAj3R8y4nWPUVDCdJdKGyb5GB7DJgn
Z6i8hPpSZomgM7744ZRv3TiSglPlVsCd1NGM04Uq4anYxBHq77Wr/Ky8jMMs7NCQ
PcQu8jG6VWfm3n6oNo3oW+OWlE+t1fQldoxGbY/OAhv9J+6H53lQ3GuvsY+NtvuU
HKxP/ObIbnEHfSAu0UWOP76PVG2mGSLbwGbPzhJRyWS65KeGM/OYC3W4BEb9yCjW
zpV+ObIfoQuGrMTq+4xqNd3f5iOFYtUIHP4ou6RRL/o6fCLMfdnJcwqk4RGWEobC
1UcYcHuDE5OUJSEoT2iuIegR+jfmHIx3COeOPidUPTVF5BPgtVEQX3Dzmxmaf1QT
cx2OprZcPPmdcIN4oy3VMHpLMHs34lvQRkgyaS8zQ04ZpMyqANQVyKHQy9YFjHWp
Y00ojz8CGDJt76bP3xqHgID8ynrDPsbKtz84SynvtHrqX+KNOG5kTfrlCuoVFLis
1+dojowB0ILzON6CNHye7qYHMjHBojvB6SVuayXoYx+QQF6epRlxn5wpmZNChAl9
E3lEEqMLs/gGlLJZRRNsuyf3pFijQ5Uv9V8DZ/W39HooDM7NLIh4benPtmgH+n8O
MkBGdq1K9qYnLOosjGYTaXaMvMXFWqyDFSWLnjBuiTXAq5Znmuj2CjWFwxDARogJ
K3FIKU0TbrftX8xZgE7s4HEBA5Va+4lMFj88W+BrDS5JJmTExeKq4SJz88ynTJCy
WbZX+daJ9aKzNt4n3vhg2g9FengyGasaHR3OimeTSzPdB1esS/JH1eeTdfs3YYYj
HEHx4nUAYjQiv2cJoKbSj7pKgXL3XgKmjK4qm7O8WuxYAOVNSJHZBbwrXFff6uXn
VqUKPgGdedEExPvhAKuFde5FT0SpEarJ9M686qkKs8vd6IeVLOYXwXQKl7UpFMky
LYdyTC+pWXa7K8vW8gdZlQGQ6kS840lbYeq32r0fC0rxQ9uMheQeMlHMXnhASgjr
cqWjtzY9G2gp97mv0u7qTXxS9ciKmR0Rjsg3fLbfdwk/t0pth7csmJh3D4bMiPEh
aHsHejfD+BzOq/bnh/hJ/6IpRm4lOsTIMANAj1HA+kPbn50YwOVcoLbKTK0MhvDv
f2+nC7y3s3uVcEHOANOgcCeTwaP4aQFu26FvHGLzlSEbGVnPkG9TT4KogNAu3y4S
anZwJHa6zXRjdiasqCKE/AZLg5ZYUFn8RMQM6wwrQ4K3/B/f38cwjEMX9gM0ICFb
B2sAiaJ/f0lqgKXAQYEotBiz0BejgTtW7MyRI5ndM6m6z003obmrtT+eNZ7fWnrr
e1eunUn/zhligC+jTn3MBQHkXs+u2A8xoV650nF1CZcQwvnCGwYb7UiEGevNVHGr
NjaBFU88kXSzdHF6GlLhoXTOAHET82BvZZvn7+TfXY5/2NT9Uv/28lqXydcUK+ld
ijQtUqd1gL0epRAVhSK/JBE4WRKyGT9hiiH1d1e3CBS+IOyRUZvJpjLjybveqIjo
SKCoRiRe3fGwmayoArCBZ6S9SZc8eObg6XUISaFAf5On7OL8sbj0ExQMva8B3Aax
8YPPA1k0GHTevfkUAavdQe8TgyQu2mM61mab8xL6p256IavMcfF3stRbPit8eJTA
y6GGPAeg6yM0csIVagQmlnVZSzGgehcMmtPqaJ42NiGMOmPCcpFW6xBJ+qmczl/G
NR6FTftrRhDMTcFcKY2GgSP8yreZuo1AvVSA9A0rNgNABil5SRTaYI2mKoqzObkc
34RcXEnUT+L/1Iq+HJk27BnjdWWEURlpCNo9EHK5ypqm7NFpBZylB3qLjsMIzNpw
lilmGCgNBrnQkV/mhUhjdZFnlAc12SsuO4em6qJ5StZ1wr33ndIWkRClJf/ediRf
gmrwojpjVNIi3mTsqX3TI+cOIIPWiNUgIVoVcCsZnirLAAqnQt7fF4wASu4LhqdI
LW8jcqu8zh4fYXRpaePHhtY19y6EPtOCniy+zqrotbwDny2b44XD8Rx1xDELsm5T
azNKdSo5QoOm2PiJooTudUPldLura9v7lxeargP/JyDx6w6/D8v4SC/Gn3oXvDGD
ps8aWEtUy2PK8J+hB0lV0foSEzbez1R0qLyS4OGX4X2JWZhZ9ocqEbooDvSe+Aw+
pul05AJyav7TCx+byypro+TLgMNR+MyzZn/exmyt7ObKdrrRPme7fXre4iYdYMRQ
qYa1RMVzLAn8bPzYFRa3Xnt8rIpeRLV/7OpgM/E4fIj9f0LEU42lu8LLEZWzA+U/
ecxO22Gps2ADngMTo63g04fwI8tuSEp791c9kNuVQwLXaq4gLDOL/j/FqiYqrVVw
dEKraaVAjuR/orKClh96uGSAD2pIzME3xb+mcjmXfs+ye6g0Nu5A5ks1nT02WUII
19Xkv24rOuJ5/k8HcnbALzasNuL2prqyP/uUhHOm81Obtkj8Wl+L89hhtzYbJ28D
F42lDhp9s3Blk0vEYPFjtTWErGJQiNmXVZ8nTY4g6P11uCweZG8gwj4TCx7clhoT
FGvg0W/dJqhbuDMjZoLUIr7iFTv+MeAlpDrlFW/JHZEZMOVPLkUPZxZnrZjhli+P
DEkWIpFcb5EpsuaBzmKMDy+0Ikj2hiwfrsd+6mLbkuXOZjNi6d+i6ObRGPHnVmTE
x9l+HfeIQKZQVSNX+izacC1Eb3gEU+oFVgWjMeItatw9I2Dg5gdjLpmyig2ceP0g
03HU5t5CpFYT4TwfrSDuNcjJYjkKaL+fIqrGilpHuzvFx/lvEVptqtRPE6KgaJu5
7TqeE1av6ZSjz/XR4bDBNH7wgRBqV8Ds2C0HRDGLeH8nWn9k3iAkENIBB1v/t1fl
+GNlfcPiSQDbur+ofB5peQVyTz+HrILr26iu8Vm47LWS6WkbD3CMwvM6tX+GWrua
jwly07UdkwrLNNrRVPk+Q5WQq7i6w9+Kty4AMK1XuekqoOpR+555niV0Hm7VXFHV
BODr7Gd2EgelQh3keei1ZVcJmoz1NwQZdHTCgtQpPzci8q1rgQlE9F5LRWPuHJ7a
A6NbTQmKaBhHesC7GheKPv5+GKDwiXVzLpK53qS351yRMbwdwfBaRv4LQpanxy7E
ju2nMjq6qGVwxwhEUI0yuIYAcAklVt8Q92oh8dluTiKo1fa65r/Ne8qdhAdh8DsT
urA5ierGpZpi2ZIS7eQ/kMTGBGeaRiLW7NSJmU6OAwdk/65Wz0/AgieEnsesLK9Y
dCYREB3bipTDOhu07a8uzVyRjc8nB645SlAHTREEfo1JfbJ8syzy36UvlNuuSHLj
u/3r5Wj/qCqYfubTtXAwu1F2crQC9+KrleJfU2m9jzMlxsO6rKo57aY+6gfMFajB
NHqmiIqQYY+PNmbdUxZ5DIEM4p/ECG3ZjvJD0Y7wVUiF0RSLmI2035BBvCUmTRpd
TdjkoOzaoEVYrejOkh6gvUyQdc4FzDat9UMXEiRDd7GTw5g2f58H0ps0wKkbFUmJ
3YvQGflj19uh9RdlTqt1Z1j+hzD4q5KQFH+e5Udm28lh7U8Cx4b72wJ+/s/DgeYV
pN118rQlCKhKR2qVHgdjn6uJLd4yyIOKVkeXdHyRsDmKSgZGGJkSW2tItXUl6d5u
M5/sK7JrgE6nFir1qrfYaLwjcWTuezh2LqNVNpnV07JF/KiT/cl2h7e8uSmMdrZ6
prV1irpE1TN28y2mI2ppnsSQ6r6CQekS+AqMUvNlhMlskQ2/89uanP61h+CPMtAj
mcB8uYJV4b/iiR2Exs0evrglHbarksafDrB85rdR0Bm28IVDC0LcYdHzYTdhCtNV
2qDkdmQQ/asZyywUQculOBnnIdYQ1VlpT6TFEZus/VLwZ1PigbVvIN2z+mM151Fg
qXz2/ID4WhREOY8ky3s9Z7vvJ5JY82FT+4CavQIaC5WXxNAn9yHLJ1P1M0pjdScF
sqBnzV2lKiyPryx2kcaaAMW590Q4KTn2D6n/GYEhfCCn/eBby7UKTywpF99/Ho+4
V+TqRaSGS+GxJBZ01ChH7yKgpbZZBIyjXdsJmrwYk6T3JpNjlF4Cf3Gs2eXyI2fz
Nr/8a4Bq7E9ehJFqMhEbYMYv5DM6Aosw29m40hOQLXfhJ0ArIeWAcw2N7SB5YzT+
7nDncYwl9GnfUWd7d4JmeVvLBFWp3M2Pyi0bSu2kJvHra0lW44f3uR21BUYYUvTo
HtVdpfv45bTL6treLt1mXigngoQCEDjMeqIiOkpjtwmOqWm9xxBySJt8ipz1blye
z5idwe1mIHcdey6sLqQycjxer8vlFIglfZEjToLueEoZDkF+Nc99NgWPBB1a/DOQ
7PwYnphms/tZyuaCENRUH3CIKW0lA2VV/x0AmgXO5XXVgo5C2uvkzK3ZxGoZrBDu
Qiq+Mmbxs8Ey8NrD0OQ7cSHXRPOT0eIO+PIB/Wi+1klcOXfpgatx+q2jacwa7vvo
IxXpt0g9YGxOGPAmybKPh+CtfL/jG7psaoYwF7fIZaChO7o0SBIgATESi9nsgfYC
9eLa81M1TR9MIQH0jYfLJh6hHgc0Db5kJKEXJ88xKPPSq79VWaAOgqycN6DOJvZR
oahxH0HK3FbUXsoTtphOXi6/0Bjl0cG4x8YvjoJVR2VSr6AXzQU0AvGri1xyI9YB
6D5mjhWBWf8GmG6ontUFLx65Vbn8+wkWmOy7u8Y7tYGlDI+vvv9RLBFV5xK8IJ40
iEEkTKogPBC1j1VFelKpt42GFj8IMyzS6+nX8lX/B3JfE9seWDHQO0HCaGmHeSrP
+AWKeRhAGQeWWhNcw40jaRqgJw5q5q9lRwkAWi7ToU9MaotiWcRkBcSC96LYNzTd
O6iqV6oHqjb4FetuQFUNYgr30/w2CaHmkQkKdBt+b8E/kph/6QgO37KeTN7jmtNI
/oSZ66qtDrXnNkNt6cs0vx5aIoX3mwcPBjPUGmzmzGJ5hmgto1vsiN0a54aLGJ2S
7C3lJnzKFtNfHXbacu5yCyFZewe05XhqjqVQa6HGArsmG9xaE3eKzMTmeV/KwGPO
dzhWmer+WxyVMYW7M6OumjRBi35iOe+z13N/wZsS4eB9N0p9Op4rP9F336l1Opoz
OQb7ai2hRFdiZcOwiQEG3T6E3/j32frHF2MOT5TqRdTPAfWzPnUbkgR/WzvuVMdK
2Q7AkA5JI4tY+psE/VsExFGH8BOtTTd0ceRcDrIpujoWgmPQXWXNk+6H44zNrgG6
dXJ0/ziE4jFRXxwhtjCssoauNLrDjg8u1hTXHexgab0nGEeqggK0eSbVObecVGSA
2vrv3OMMtZKysUxmUYxWMygMxKlqQ6hEnGprZI0mZe8W89HAWiZaEqYb9rt0q2cU
KQMZPKOB2pW5S2hWunqVHRCGjf4HMLOZPtx2Kl4KIKOURu5xFAdexNc+UExl109c
dD8zfVPef+Dg9b6bosW75ODrma8Bo0pOdYxCTvZufLdRXX1BMQ+zFLIEFoY2WvFB
GoBvj4XLfBHQIoqPo8STXB2nP8evkH2IcTG/+d2/idZLnYfvYNwzIQoPJIKP9OVo
5E/IlGZ7Rl78hk6ee8fJ8CiHgDozhxif8Qjn/utfEr9U+cydgmzKRO/xQnDX5bnr
XMZAmG7PegUSuHRU20IfybJPnA0V92umFwaTea65dQwm4IZt035oD7J3cXJiqfGh
jD8aR2QdFTqTQNA3d4L/ScMBCg6zWF9dDJK+vn/gPPtfJ3UVIEw/J5WKeeZkrmW3
kPzNvARdqNEVkybwbSTuzT96vrDhnKW9RoVg1e6YwC7jNPFZG2otIyBfrxb/2o4R
XgOgq8M/IftiqCWJoImEnBMOagQGNAsbA6TMdOBAHq33npJ3xoHHh9g/SKTj4ecp
O8XDENV5GNTshrXjjsa8nnXm4BNUs45C/O2qwFYDav5T35dvvqq8KkAo4UFawwwa
PWSKalpLSb1oCevzfpZXNVp7KZnUYsXHKmqmnXWkey3NQHkdlly5BxmJJeH4J/Rb
QKksx3/9qsIIXCs9f8jeWkgdkNEFaH7ml+uR8OEWp8hhNB9+aiV0d8o8EiiEdjTa
uh0+D3uOx470bxDE1uGLD71z0nj/GcX7kr39aS3uQL/3FCkVXTvI/w1TjlwjVYJ1
IdZbbj8lsalJ+VssE76tNj7dMnvSPZB1v8owgU+50rMPul/RJNX0OfSAxbaQykju
sseArf6viPUvtBv3J/GUpEjJkxK9OGC6iWSzjsimpqifuDLw6B3keN1th86oJ8Ia
qNsPN7ChT7yRH+xR/BYJCGR1qKvDKWc2ENipe7VjMpuPNkj1/ciZhMGYw3vnjvbh
YvT8brt4tAYjhXOthhNgy4A5WHK3bs94UsQMx6QI/EYxmNKiWET0mPIEFpd8vNh7
60yNQ7LE92AHDWfsAEzlnKHRR1z1Foy8S+PY9ffigY3bVKEO1a0j4R86BAG55c/s
5ceRcTcyNZW75tVPgGPtaXqYRmjPENhz8rUM3MuyVXt/k8xCHRwOX0tulAqqHElQ
5xZB4ItZU9vFKYfr5pPp14EQj9b5EyG5SSuQcQuwzpZZ2k+YB2IXaEFsXwemdWEn
bvEFBzb+pt2wSbkKdcAW1a56/pZTAnRe+CkbCtm/qV1bXPtIx1Eht6PSNQgwNmMP
QZPTIEHcoTDqBOAibxdIDrKOouHBRnmTBeU+dbjMD1pbhp275rNkX2+4+O6TmTo/
z4ra73M7o9Jk27p6zZEkVLwz13/x9ixPNfB8iWjFIao8scPvnIUFp3A9GFQwCMLh
UfI1J7gBDTgAHDUJnsrx2kCip7+kiuiaXPqQ/rxVNU2kaTZUvojKk8dGSTxqUBxL
oSWXvy567P8MVS+TeIuqIRegalNGkjk/qfwhqKNI1Uk9qvdFYtyBdAq9f+NXeo73
JRTlE/bHNnGoRSv7qdXgBePD99HV4m+dzbhSaNTYKDdL1VyXiWRfHIfbJC4e9+e5
eutACxOxRk5X1kttTGvHxfDOVcH632kjpAB7gJsNd2TpvkqsoMp6IufzM7Ux1x0j
+nMnrk9Pz0qVdZGwujmON/VcpeIFcoKV9ssAZpYS7U5Ws7XXmKC+Fz7XisLhzniF
ehcdsu6SDqMcDAgXLiHLA9ZjvV2pTnjWnsRupyhbpEkd3mC9YIvbkyG2Jtd1oPcY
idXBIQ4YqD55rwrxSnEiVgeUMYEPSDUWhUwOoIS4Dhb5JCUOI8G5xEi3LrRjlaDn
RbaC6Oaml2BRVRyxhxoOvrRM35hJJYi4+euP/eFxE4BAM+Zu8477o7DpCFEEZubm
LrJcyO4hV6l8BMx92Um1xXS7V/5SgHc16Z9xo5bkNDcw52GVeiRX9x1cZMK+9UU3
mq/NvSY1rddJNUy/DGMGEAP528siE9jKuec/qQ1SeKyzMXiySphuWTnW/UIFZ5Qq
QVMzd7NHExn9d9kmhKjWTsAgKclpRH5LuMMqP7ahAvG0edYe2r7hjhZGzM5HmEBX
Jb30u+q0gT8KoMrVbbJieQjiXvWnqmaWTOcULwf1gQvqnfaKIHpIeB6DKGm0oPET
Ku3PX962/D899CvnVJka61iXBk/Yo8kwekoKeQoIgaabXfTA3jBd53U4g20of4SF
8kWirvdlizImp/GwtnR71qpJr+7RtJu+U10ZyHBg3+jJq8R2ASB1r3lnk+lzMrS6
1lcyzswhlsvleGzl2EjcdiuWxPrKABubFY++2vUNZkYR5SEhnk4BSUdh34s4hT4l
JCiz6hA7o9mlSPAAAyP9eSU4vuHKs0Ae6nSrldsUW3mbmFYXCgpiRpwBvwuOBb60
lVioQpUzQAOVwHN/zkN171K4FlrEzc6QmHhZvp1wqr77IJkWZNqh227sAwGVWNbi
Pza9tRMuf9THCghyFLdI2gTmyoD528TjNnerNh3XRqUWyZEN2xGY3AEH3umEJqWB
KFffjFFhgOwi5cMvUcF8v762Mnh3Xm+cO7XgFz+SYKVi4JNxWmnwuVMWSMAnnyCC
p6cLpg8CIhAMQU9klS1CUItIbaTXiMkUrDB7YTLxwkKvgkvqyhcVsEjSfNYC5Sta
+w6wxcHGfNkxxlJVUiLVIFmF27xP5f6BGWu6vCu4da/n1VP8JYLEtc4o0Ffv7BEE
4VqUTjzCcGG+5ZUKyeyiR1KXnUoL7/zDaS1AKzIa2n46DBsZa7i76jGy+OZuGREB
70EpydRsA/1cuNFqORSIx5Dyxo2ed2pWtaKyGLWcUmwEQc4G588Y/CTreUbwmul5
MOM1d8TtQoZUxs5w1QVQ5lLLB26iCHlsSEys6Q54kXojvQt35saO5n91AdFXpnkS
cKSsY/I9J/Ds6ayffRRQP5Vt3htjZVWg/aSMYxR/K6QSpyOSRLCtNB+/PuDR9xsl
mPwEAKwvI6stdMzTXn025V5AgacbUue1eFQnriNWUbfLT+AHoZy5vbv/LB1vKYgu
EeNbY1VCRCx7ngBOLJGBoqRjE3/2Lg8tmXnfDJeYdfkCp+yfz9WqVsRnjnCjdOGF
FpttIAWZ/TAMwPEFA8R/DJV460qkvJetOCkPc27xlCxQqSNWfuzxDFeLLfLimLLG
Nqp8oIm412c8GP9MwJYUo0VImVAxcB0exeDdUeE6h7l//j85cTZgikX0ds9EnHY+
57BjrH9Dro54imLrR37W4goImbIfrYNJVOl5FYxtQt5ayZC5wiDsI4XqCC3PvF0K
QjMwEMFyEWDuNm1yngwFRO61ofM+JkFnFdMoYpW2A8YZp8P7jBQmM2/ckd/VQV82
vQQrH4swcMUFHgo+DK3SF3otraRnZSet0hrquTXl5ZCR3jBitpu3KGsSDgowNDjZ
IF10pBAEW0yYVWwd97wllq6QZZga3qHtKivrr2g6NCSX1coRk3UnDUsJ1NpBqnFI
EaoHXqjr7PUu9mWfJWn0pqn9eT1JFDByvAECgHM8F5xuoK6l8S2/e/DTFhcYm/GD
qGVX7WL2/MvxPSdRtEXWT5lTKj3XigLnyW91a/+txXb+BtUD7X2OqpSpAgepOud5
e97zFLmnVmvuuJouQfPZ5vs8T+R4phi+dnf+XQv6vgjnbUeQDQBpEc1cUHBN/sNX
LV8+QrWUqG+qwV+VDWiT219BcqMi8fh3e07EZGk/iubofhBxVQI2aE58lJLneYKr
3GNjXC+yCTHe7hayk2zbCt7II6jW3PD7x0u66e07JnbZA+smNPl9BPdFdzvOyEIO
IZalh1A/Pf0ADuwsG3gDCIr4+IPux5M88ih5Ntxs1wSVEZpX6XASk1VxEa/nlRfP
HwpKJirbElW1XmpJs+7uYplqJLVcoAR2PQn6BbcN/+MR7p0UU8262QRaHagKsM7B
pTyWEdZNXCapL009RIG0DatEIFUURA+gceS1rUlOtFOzgbJyr0obe54F+xKHKHRL
PXKFyTr7ZRHSERHj3MiI7Cmg/k6QPGrarcWD8R9P6NNlhOYP+g+6dA4OAsTgExGR
GOY36bPtmXxmBVTlFbJrHGuswU17pyr3QDy+gC8tneBlO9Bf7z1CN0lWoUEGwZMb
SIsc+Yzir07yD4EDAPC0S3bcLR+UCEug2X+IFOcKDJERZ62lNeCCNPnG5HG2g8wX
xY6fjyy6MceVNdvhwvDUtLzZcUpGZ3WhYex+2dKxuy84vbQ4T8w+AFh35BjCzbuw
tzA8+YXJLtwgiNXzyuI+J2XofYJt99jMiGPsRw13wWIzlFMWePEjgTcGDskfwfbD
kxlf0EdOO21m9U0efHQuykTdzinBWoLtXjuOT1kL3kx4kuaUWbdgP+G36kizpSsg
Fyx8wTWA3dDUgkJRFKZ9C0HOjszUCqPwixLC3B3ZkTn5KILX3DA4jkLNviTSDvE7
5JOSZFqcA+sSZSqxv4w666GgQ2bdiwHsozFLKzur9bCYvOhND+2F++WYhLBv1QCQ
pm8+5QigOm2DwOGpnIJslyKh3O+WZIW53LDKsu5Ya3318ibPO8YTRgA5kKY+/jXl
8EnxrwsjJvaXFJaIzfPZABb2m1m7dVirL5OPNKyfqejRuhKmpCJQMi4spu4fwGd8
QckfBT1mkoAAm0Ch3noyCfhnpGX9WEKJJEAxMGAnX/monYIInGcVbpCITnPhIC64
2v9j+ozY+B9oz36c6TBIZSak3A2uSfgDTDBwsdaq4q9H1Y4kZ3yseYb/pFbYHI37
qVnzikpRovnZroYHrt3/B1ch9PmHrzNACkWKX8UITFpL6vw0spm43oa4y2WC17gM
u8/Ea4qIlnr20Za8dCgoBv/osZ1PEDNX7b+xyEvYDNAtplDAWpX06pQC0irUDcnk
CPKfvdkgnYyFYvAbwpmISNbHPWkLmhJmVaIKsfuib6mXxNybkeuMrm9AiKrZIj+h
Z2kxwG6Yd3sROdcfcZUmLdu/YwbOW9qcwph6VP0MvVK2yUWEm2h6Z01CRN54UNT7
pxlqom/aFNOfa75wMi09dg3pnllfThBeDjB2HAdrEAfQUBgSOZmfFNdAAtymE2cW
Dvmt57YMbAsyFuL8au0DlWRhiKVg/NR2FWBIJJlZ0xZReeM8AHCBixGv+fSzi9PO
/V30TJ3X6cYur97Ltb4ZydCWXCTZq+vbTkbYWGf8CjytsPzkthZNO1+eBUBhGbjm
5rHmcDMMQMuDlNcO5PVEMtuYNPzIysiQ9J/urVrW5GrjCKH3Ja4DmarDAF+PvoX2
+w++W8SjAbVElSSYCDh2yLgXL3U4BuG+EnE3aNxmKuXqgFxaeu8NSYoJsWqIm7mZ
XMACIMRBXaf0Jl+pnw9D1LBKxtfuWkf00fWb1n12d1IK4Ctb3jYvkayX/WAVkzGf
0RvyM0KKLleRdCV5oDtTGWK2++lNK/EHeJPupa74X1nKqHqdA6vZ/ptvki3vV3eN
4uUzvOWkEJz8mt9XTP4PEIUYmCZSNlRQ0QfZo5yAnmy9tiRVkDOT58JJ9J7q5O3X
VHITDob4owXwyk4Cbhrvj5O/BGsLtHpySp6GmbKcgOUH/rfsqoWG14TgN7NWqgPN
14gIhC+6sOMCpR4AkzsoMFshqkuNOuP2qnKG1BKEznkEvl4/a66Rfs7zAcakn8pM
JCfRKU7E30CfLFgpea6RtICBvXQouqPpjNwoT65EhLZwF5DyNWFFDIOdpDKVnBzt
QLEhG4FZVHycTVLaMC+kygcbJUJ0JS0IJPchAZ1AF1A456y3Uq1dzPyKbbNGuaa3
LkoIjfW6iYeAqvsIdT6n9+Ktk6ckmW3ijIkHe/RvGIu7gI7oa07ztB3LRDiu9lzg
YVECMVmaAOM/lxQvuNXz3m7QnFYWgY03DVjZpUWq0eniJUV0lDiJSfWUZxz2Yn45
5YqxNaD8abBAmyX7a9PafHYVbmPsJfhG9l/cUdknR25ivUXJUp0h+LwTQqW/sx+7
7qu7pgv59Ynv8XC7eyV93SZiAIkCzECRAlO5mCKEl6oqcDdKMGvNmKhCyp6r7XfJ
AbygcUfoLZcb2BTp9YrR41HRtDEwzh5DY288nW2Pz/siE91l0u0t+4KRj2FVQLBO
pjP114EPfpRCctOxkc678wVoctWxEmXImVAW/k/MTp33mbRDG0NyS8ZtVyrQhZK3
jTeQj3czPWP0IlmAcSJfeD0wH0xb5ZV9vZsQQEaVTpy8uLcVO3ocoorlIKyjfZ65
rEJFCct0pV1ty4repKgDI0ChNy480DX9FNXT0F0yA5far2+31NLhPtOqqpHHy1im
diF1V5t5g1KcIr5JO34ajIlqdNdUlePPvUO+IuG08mbkU/zAG7wcwE336EtTlgDu
jiJWn/qsdAJ35Dyorc9ULi1U/FSF9GlZ23sdP8jN7hAHJ9Vsz81LOHPk81pKeMQp
wcY0T/UtTgJR+CqCJK+GlpYj+jKqkEIxmvxHqPgsfgNMwkqPUAeB+UPKISdQnNTM
V1HrQLCBi3xE9ws7aKMzHpeZ+5S7KgotyrOpgl2YcIaOhGn2cHCqCIicUDus16bY
m3BWaVzWi+tz9apA+LqQeheHyeIKQSM9LOokke/8mHq07PFfawuengYxZ06BUP1f
C97rB08afpPFMipFF2jm7zKRpksgAhTgVhD7X4fRKu0zUzdUKuZOXEKbLDQSl4Bh
t7WltmCy9Rt4mQBHR/umqm1c1IHCP7M4g05qIA0dZywjq1FeZ+gszzKaC8LehQD9
z5Sj7mTuT4dW1WX+21FFbMZuYdteRwsKuV+z2TP+x7GPS9+UB8/akWWaUcdXZsY+
zpOItX5TmYq8UL/+so3ID14PFY2UXXu7wXeVlH17M+nxdENWS+6h9HkK5jMeRaRb
FUUpbTcVEKzg3nCyKYhmTl2RBanlbEMhP1mbPPK6NF4IsAjOzbK4auyX5BPGBDHU
KKsgU0OXbjIHRrzzWXunSE+0QwTHj8nCqhDk5Ysx5QtyfLhCXbWVxhMnKyi+Esc4
1o4URdrdcjHeBjwxXWWIrGtioCV/ctBwg4WS0Wu77DcJBBNVjcY00IfFiSz8LVQi
jGsu5V2QBX+n0j7Ybyux3ws8zp6n0MCOQtOCJ5wUneCPqst173sIJPudlr5q0OyI
ytFSpnEzzMXZ/x84T9D1hFzs7lRrg3DqwO60pRBfZRaHMCmWuuje10qDNCHgiw4X
gSq86LX3/x+aGLHr2R05WTnCv3S4kmjR/Gw5zfmee6V0assUlTbFu4v6D61gb7G7
X3z6GHBoSQ/6+v2P0AHblTm6noS0n3lsv/b+/NjxzT5WAKvSO4pC9XZqwBTc/uI+
WVcZNKMiW3DDOKqHQmfnaKnVyMVY4LheJLtRiUaLsaTAm4KYHWjdZlV1GVU7UKxJ
YX0loeO2ik//HhSAgT1dzr+6vPYdOV0NOjI3HdbksWIg4YHRfYGj/yMUxE1BKIuw
SxaHpGymhpKO2E0nyxS/deGDBXXaASQPNe+1dkaSQV2GDMQv4RH7ZXWv/PEzBWVF
s1u0n2n0qIpFuoDBvp9LLjAedGBe77xDzZ4biZGGwMIIqeJbba6q9yvSiiHp5mF1
W1ENnGUYpJds3jDwXnfnIvrR7UB4cB+9cjGONV6OF/peL8boisZxlsswKK2xqLJl
s89syhY0vZSWdmPc51WoTjWX0keaxjd6OVbJiahT+OGnR1tO1mvAMSMMQr3HR958
3rLgmZLhs8SByCOYkzcnEZyN1CGA3L/FKLrMTv90Yj2yGiZ1PVArT9Z8qZ6QjNvs
9f48bxDbD2GgvYe+frX8MiwlAwrzvfT2o/R1rHTVpO/1JDaR/VvJD6FjnvlUjZLM
H6WCGqIhtyeEvEZk9M2jRd28wiDT9AcoTF6w9AxYQb8EeY2Gl41mEyuXBZEUpgKF
bnsNxd8xB3PO+TsmNWnhrsOLLbq46lnDranF6qwGFM4tXrOBus68nTbTyQEpoBsS
Jsn9QdLzlhb8p1ffJbKx4HqML0vnDFJ373/0OeMjpTI28bTie/UGyKtxyPgNgmeu
sjfIyqSFykWIMiG8x+a+6eopfcKnGBjxscUvA8Y05Ve7xX94AjU+Td3MhhE9UnWo
DcRD2fdL2fsrz5Huorrs9ousD4awZvh/ZSDJOMJn8s9IBRWzqJKGiEkPgHSVuQRD
/fmAzZPIlw4MKJ5RLJNSw5pURZYMsPjt5UaekqzIyoXeler0ZGn6GeXAT/IMc7YG
u4AO/K76NH2vYxwI27Bb2WPLrEWQ8OTmkYOpnwMAWtXGXRW/d0A1gNqYfwG8Ew57
k4okZx8wDr5mxPELDuW6ugh4Mz3Z9IZiGrnxRpMy70E8pyyQtuncSGt+MB/3s1sh
2EsmzmiiHO2Es5U2vRWPH+6SIK0fIpYdaeMWhCI5xThqeLhrPLrzq3cIzqARkgMf
bHhF3oMbEXJE9VlbeendThDLiKjzuTkiA7LlPtVJlftX3T3DjXcprQLNPDtK5IY3
IawHAVaEqU9wJ1VjycZRLff31LL2CAoTcHlZXVRlIOiH9YbDxN2E8wYNPUHsh7AM
5itOpKRhPHvKe3R6RElW0j//dicdLsrp48v5PxUA9syKp7TUkY6NGlIB+JKl9SU/
B5IetzPeOzNMVQxX7HBKE6+zEpFeazapxVfvG+S7Ce3FL/BGU0y8y5z9MxQ+Wn+s
yk9Gmkd4QqM6VDtoeKFRya2qcT7SwC+yvtD682yC6KPJupOj0wvH8FxhVksUd5p9
GJvrmWsMGPhtVIHzJktJJPu05dknD7KYl42xwlBD0dfbi1Ry0Wc1XOA64W2gE7+M
+BBRjqfzxiBWiyqUPs/h9AcBSRXlfAfjASlkF84b2iuJkl6K1+k1W5kEm4XONZMI
LQ33IaueBbJp8n+Y2cqtr3ttI3mGLvpJRg4UmaanTjMYCbGQaNRy5V28zJ2UGV/b
Ge1KNJvrHFz8Dwivsc9RL3o4UKYIa5Sw9A8gfElvoAZ2PMsCMhKf35W/DV86DMKd
82oUK98lqt3tIHAhI09Bv9JIfXzsN37yoly9uYIE6pctr7InKYs2gpPT04prYPOv
2OVbcA8+PL7NBc7MPahYPH+YuVSpI/DcQZUshLBpisKfcFI9xajUfMDwi1Lvcfwq
WoKEw95s7Zb4Tf026r50yAAk2/JTVSmHMs427evGZctYmQPgK4LdDEB1g+PbWgcq
m2rhHRLjQPYMRQyO0RYgvioNome6ArEAhXmP44ymjFutOq/Y13b94ZafQ7fGmGex
FnUdARQnPibkobfU5uioWBHtGtsC2uMSL4TGBSLSXeeKLSjtyCqneORtu6rTo3Mn
ohD2gvXUV/4vbXCjShps2TYcwau5TsXzQHpMQgR893L7UHsdYJOlBKf6RPXaL6RI
tUp9qR+Jba80rwJODT/6cVBbtxkkgGjcImufru7/hwzKFUCYAthvghdftdCAGQ5+
kxtWcR2zm795BYvlV8s8HHtfPvQIMD7vsl8kJ/HQqBMfv1eEDv1vuwi7lT+ACtBv
484GPGQ3W3jEIcx+t81C76n+WS1RRa5SgtjOmBlZvr5bo1FoBhx2IvhX+HKnTNDr
nsE26VZNW0xBaYMxwboqegEruHGPwlE8qoJjYm6cqp0MCGmx0KbtNCPd9CCBIBcC
aJXVi1cX7R6PxfXV5cE98Iyq6pfQZCEvftsnelRsXgIjtQ55RFg3bBsocV95ozNG
xV49D2RISOYeiMy7A+mMpLjpVGEjS7kWyGZi7II1Hjxvx4fWW29uPUxsM3/ELbO2
zKKeWDnf9wcjkaOCvhVtFuZMdmxmIwip1VdkFmCL8NmD9J823u5NiDtODkwRYHw8
tYUtCETICMC8g0I/EPwZGlMrEhkhy8RiHFLjdoNKlze9sP6Z46rgXY3UwRS3YDHK
C7qNgCwCqU3OOYhHdlbltaCJywKxNOe4JTFb75rJ10vP11X9AEv/pZxGMwZSJ5vv
l1OAHnhOpRjo6QUKGudHkk1DnOtjtw0aN5HWJd1gna7a6JucCbdkVMqSbpNqPnY5
qsT2neeG+bdI17NWsDDc+lWqDy4rmy/iHFkdPvITcxn61xtF8j/NHLwJq7kAWKpV
0ClaebM2ArljcMZwnFNKIXH+sICk0xAZL8MVIlO5yw0mBP+Qcq+qZBqjCxprf/dC
TVM5JdLOpqWagSEnBO77Y5JBjP9DITGK4/vaz5IO1lth3u1fu4yS+8utgQCRNSbY
LK4+qHVrj1lChkqUgFKL2EkPInUoSEBFOOp6Z7vDaFzYxOdaEn+7v1bxG6nt/5FV
WONVizwkeUzTsB+64VZLFGoEhwRbJDKjPqCBPpijNwx2j+QCEeSpJ/zfrY639ebw
JPgtyDFwAgHIdvIH57DyEbJJMZb5iqeNNNdpW2sz4BcGZue6oBahrIyDiw+27IBs
F5bLGkD0p3eePS6Yg3sIRG251QziMyhrygRNtTH6pHa0jgEP4lN3OW+US34roTmM
gLe1CG69eE2MGH2a+z7xJMstS8o8x3P20ABZqVmx3exfF55IfZaz6HolodDtVm04
/KPWIEU7PqUN/sk7cHTGdfpImXU5uTYv9Soj3o3iGxG/A8b55F0fRaQ8o7jmGbCL
Jihtr8AamtYPAX4PbbpNlUgVQQsy3xKtCTa9MzLatDE1cCdEpkR4NPQ037QOohJM
RajlNmMIkWAiCnj44Oc+M0qk1VPEROQNc+f5LBpxLvMZQa3iOL6r+RC7Y5Axjidt
axiBmA9SJohQ0Rk5Sq7QbxvbwbAa3YvU7rVozvzWv6lOI3FhOsRj4/3fEFePGpC8
ZGYrvHix3qMuHlvOitV1QdhmPsmx+kKguobS1RqNDpaP2CRTAqq4rRJzTeGVtwCG
yKJwpdZhISoCuzfR31fL7y3nBtFgUokxQcoK0xoMqV1iN11dFoHUQVEBXlGjs+CS
U46l/reSphjdPxHmnmxj3oz8GY/tnJrQyhl4Kx6xWXI4JViecOzUQPyhNHm4dG//
XxFbkVZsZpHxmXLgtP0ZXKKGQ2EwHAU4MDRHmtti4MqLTQPUnvu6SgTXAewBm+au
EFbRxAqKUSs200KLCdFSijrs7Kfak92HgPu/N3XWdzsxWpiFWzMP8Smgkd45sOKP
vGwZeYScfnpdoLJqbCgub5oZcOyZUn/Dvfq/u290V6jQ4iC2cTXnmA6wf2b8Ac2g
s+wzXB79pdf1ud7ANig7XYwoCc87PboMiSIW7BGchcVfFNEcde1sDgLunh3BKCOP
A2QnN589VvjPUr+DMEKDYRtz99lBE1HNp1gRUNesRZtAh/+8f1Qi4Klc5HmwtjQf
6DWDD7Hq2/aJRSYYQkDDJkjceb0KonbXC1VwcCx651G0EiEDQ0GZpNmgtIcEZGQu
98RWZobNSt8LdFQDjOylFtEFKTX21tRNcBdjWXa8SccwawEuubls0Xs/0QFF59Yw
29pYkBHxeSaZD8sHkQuibLUl10Utv57ebTqggiI6kDlpMQvYNE1yyj9Y41HagarD
YloqeNGmZNTHAidcPnZUCu+qgrhvA6+6YYxg1elMCUxphHi3SxtzAVXlxGrlnz56
gROofWAyIzU/TuJtOMdJMD+A+G5v18XFvPIxqUyGVrRcdS53sdFj5eFS32J6WXmd
Q4hch8pCgPJ/90TiOC9V9ukXZCsNavdGsK+bzW+M3Qah1Yoxnsb2QKLMUaH3RVdU
pqios3Yu6OodM0NyS/0rjeyl6MPfI1BNk5whZf8brY3iHd8aXA+2tbe+jJefB3tU
a5HDqIXGJm5DUjavq0r9ZZ1GqToKudHGBhB/2kiF1MzoKLtQaCbnYV3mK+g/8DuV
PLBrqfgd5iulug1D2YW5W+D8gPuIQLX1P9RbOfnbVER33k/pEF5Jl3fby+JltuVY
+y1Idwb1tl0kN/BKgSQrkxJoV+LsVa+HF1iqQCarvQj2F/1l6S3Pwhm8sl0iUl2R
IXLM3sEESCzP1XSmKoYiPrZVfLC7A/iDEA+6hxJCxine9hfRbWyWLcBFP7jnNxqW
Cvnnz5xmpVeUjknxDDEjchOGEW8L4WxxNIEOwYL0JYxD4sM372bBVzxyG/3Q71GU
Mj5rl6AyB3Fr6qhyj7mhrbhjfgvsPDcLn1z4BgCfgFKDE62bPK9fS1TEVti4WSbR
WxNnrurXhpLkRvDwwi/xlcjzyYWOxJvdUcujZ//G814TQgpmo6hQUrhbFazaO0lZ
FgXSTKV87MII/P1+NwAJqk9sAYqPUeEDkCKGETRArPKVCmrbL8ZoWzSuFTKZjRJA
PfyfuY3BSbojSs/+8UovJGvkQutZq9dttNHgm2wYd1HoynDLjfeZF5E3dIC2txS+
tRshgu+17P3LYXjO+cklPZ7F9t7xVhvPwXbshURsxuvT5Kp6qmtAfG1jAttOKngS
brKYwr1vBR6dzdB/OQURyZ19q5IrgC0FlLSbhKMgSM61wyI95k2hPMZ4l2TC3KAE
+UOWCPZlEq22ZvmqVP/k5zhzJDrp9jaIkTzuuYUaWfGSkyjjvUFrLDW5mMcTAD9+
mUYj7wVSo599aPfa+O4FtLu1PO1MEW0VIqIRid1nJiigQ30w0ektQBFL9dWlWRAP
4cqkFigsNZ5Pi7ROcj61iVgzFlKZCWf0fR3GwkSKSriionQmlZaIVOhxzaCi5m/A
WcES7Q/ms3hTpl7OzSi1rCH+cFaoQo5lo3uOCvbMiLRFcsUs6O2qHM54zjAgkZ7C
jjmnxWUBUpfI2bPyottv0215swUXiB6wmqOvcUxNaEX30MKpCDZjT5+1/Hdx+/Hk
dFjnQEHjHoP/tjHnzSb9WBqOoLuhfG49hoJxXrs8S3SGGbzPE8H3XHj3uDfjXK/n
X3ON4Lfqsbt9FsPoIdLLXMhr/nJne9776A5pX8Lm+PrcYdAmo1+qcbq/hT5tNOAQ
nSC9BxxuVlPE1qOdiDBXPK3ze+EJamFji77eY36OQjAM6Xwe+CZ8yPN+/bFtfypQ
vKt9we7HZz2FOYPOZKwngK6g0O7z73Z/hUxoqQVoI9a3m5KnfOv7dJCUbWNO+KCp
mtlLkA60zIraNUlNAsmDJn1ZFP6UMuH+YaiuEGquo272D1rlQuPW8bX9ZrG7gI4B
RiKJOKco9fD4tAXa6XkmgUNQFXmP3gw3Z9qf3Q0HUJZUBoF1fPVakuCm1GRfOoDB
41Bg/dp3zbquhEG0WhKCYGyNEluhU6CLHBscY0FWvNVMYrM1hd6EdmabzS9GhVIX
4euLSQXgenGkn04TLnx908WAKwWYrYtqPOEcbVMdhsaOdqNw2Bfu23f5j7SG33Sc
ftlWaVXles2MfWifLwB7iw87vZrLnppIWIyDA6VunGZVwY/Cx8kp+pc3V5fd9U1q
GchcYBxCLPJeiuvGIi+1XZLBTbCLvqoJzdF61Ye77ojp+q1e1eH9bT9Ob5kLSFUk
r7CWcrTxioIe3jGcfB+E0EIdPT0BgJXzIwxKryUpg7z9ajc7dOnkQpYtz1T/67HL
f/txVyn2rLKXhh3LAb79buWvZt3BRfFUV1Mik1dsetBkXGcHQJHxFIYCCuuT2iKD
ivPWv6SVfvn5dRWqcTIWcBquQGqlg7A5iE8YpZzypPv2ycHUaXT7H7OglXIiMwIz
NuS4fnDwZhM1mPRwleZYCp/vXp72juAFuvGz0+gHxlURaWIcL6ZPYHB3VKkCXAIj
j0m0+Q6aMj2L+NbGTixiJxu/hXwzVeBSPnsveUYqsA8MTEVmHNDZL8gWNie1Hvby
HvXCnoPVeCDi5s8UmIpX7nLwAiwVlTznEvwebBXJOLBWC8jlXFyjSpY0ykOLii7v
Zk8LVz2Vp/3ftsoxEZIlU3QsWn14kNi8vy5vG5+o4GTOOjPwyqETaUKGpkwOEf0f
lOxl7gbQaYReqcSZYtVRoFViw+PbAIqKA/ox+jvo+ite9koskOZhSG/wV0+YUd7h
HVXsez06CjnDa25X0wG7omGG8wfiAbp54v2Bh5iQv1CwQYV3dMXvUKxShBqQZuYb
OFgz809ZND9jUsli4O6QQzekgkHZngHLWK0eeO9Y7H56akJFqW93unHDTeUeKjAY
rwS7sTlm25GKmq0afKbcMgqOq7fIqE7mT3QuMa9OBbN6dKFR0V3pkU45WkuQIdFN
wXxY3uWPMOoLz+rECWtg/aJYtdbkDIAK5cFbi5LcpADYnIK1evtEux6QKRu8xyVm
LTnMJty/qxd6iGw8+GJhvvdXKllPnJ+ZxxsqlOixRzGigEafu7BCw+9tglfCSW3O
CACYAhFD9jJXgIgZEzqdKbsB8LHRWV4qPNjTbnK7MMGiglCpu0CfkmTMmiex51gS
G9boI3Hsi6yuab9BKG212IO5+yYeAOFQyRdam7l/K3/y5vn7Eyu5J9c/HlZK/zyV
yICIVsCnpvJmjRe7U97VfDydbKl6pXM7JPTegIxetm2Xggw88KDD0GjAwq+O34uC
7GfinsyPBk5s1DBTV4znxycqcTEsT1AzMJZrKTZgs4jJEcHpj6ZTfXp7biceTkUT
FcQ+qm8D/Oi3QGO9dCRL73KzO56cd0nvFqEmALxNqqI2Vl7lgpkAwPsDiKSykY5Z
1C7LctwqcwGXUeBlK/FWGaAomBPEZUvrcMLqIpTTQ1WvW4RQmX1kJGh/eGXeivG9
/Jljy+cRUlDTaFnhxwAYxuWpT7LzOsR6HjabGAhvjS9QLjanD3HZDpV4y04MY5Uu
nOFbSR25pJ/LZZgcb0fOK3otH6i1f+66OgCmGfKuLMu/j5huwP7dLn0Qx6yihy2w
EC6KKGyrUgqpyPt7pStIaMVFaTtcgmXh974Au/r23/klu+F+DCUbHSodMLkhdanK
oTCHOjuptIJmCYhlO5yUlYUA6FuAAU1ItGeT/bxaWhiAraCNwIWVvG/8QXzq56xi
hIs5eg4acuNtSLAvMZ6fS2y3LAz6RItLvp2587drfcKyJ2IL3dZ33FE5pjxxDGDq
07n2aR4KBb3Ka1Olba5bUxHTWSstMnZ6NEFvcZbHa25PU2Og6yQmrf4MDMGpcPwj
KqDXGq3aTGbXJianUlxWZUgYCLdCG2OPQDxyz8Xxi0NJVfKpqWf0wOeQTo4tjraT
Y1fuBChRbq3cBqjja6vQHYSHYQn6cRXN7pKIFKhOkOQE5N6estvrpZ95oeGPyA95
BT5wekL/4OGwZCHr/M/BvZEtzgRwQpXlceKE82xZgS1KhZKCjjgnfJD+bauIRMg9
y13+O5J7qYmDp6FuWMff55/2qN9Ols3BF7ug0sE7dv0Y0EngrMkLLB76JYZaiKlk
aKkrHOVsyA0/Bctm8ZdE5XnD2I13btuN2lFw74f4GQDYOmKyRXZ2AtSburUndTRh
KzTCcP76IaPM8j6uM1Pd27Q7W+lrnd42IjV1ZCp3ikAvTQQyIL2fEGlA4lMXOmr4
pbzqJFuVqTTzFZEEHoem14jFlxLWNqPNcBU9SOY1w5ypagtAYTrM1/460gLpvBBN
/FtC7wOvo04J3reE8F1oag80z6Qj+XDjGTcdSxDcPnDzFkpTNH/Gfz5E6bMnJZAH
QjwkH/tE7rtUx+ccQA5rwlwSe+7cgugopKe9Wam2pH9md75vjnWz424TPRc+6NyF
uJ3VfKDICmjw7frmcdkvjSnMXN+yTq1C91d+SqXtGLQcmZo3+dousjXx4mpC94Fa
U5l8aMfam4qqgYx+5PMVH1v11GYBRbuW7/ziZ/eIqDnw4ZhFCBtz2qivFk6kPa/x
c+Ad+TU56J49mi1qdQa5p6cl3jTXg9cW0vcuUz0PSCKEbZQVoEEG9n1zKmxEMJlk
M0OQGbVUdmFNh/hRsmpuDlMJCnlcMR4jTGPg0b7Sl1yoR8pPUjzmbEAsKKc6NCpf
EqCKLYk1uk4+xOzgCBt/GfRbhk9MsG00JkjqOhGoH50xRJ9l5DkIBywkDVjBQgrX
NdDoFPkt0pk2UzzDTpCcjtcDUEAJcfjsndwl9fS7a3aRxCBTopNvz7efi2p6dGb4
jlADrsvTRXlFUgY2cj3SF3uAA78pYEFmf8UJHJKF0YCSAmKPt3uLU9EEYlWR4KyO
XjBaUQfgOiXxAq+jxWXIdFNgsDLyP9nvo9eOkJvgpg9/LesfOaWjVFQXl1/X8ppb
yyQYT7UZ5pFEY7ybAv1OCrYQTiLH9K5feUCwFieXDXrpbnXgoVyFeE13hC6S+XjK
HHyvXUcJPdKdK5GDxafnRobAnp3JGDWv0X/holIOnrB3yt8i284D+7ixepVwcNqx
qcX4Y86xg8VFnv8sHxpbAzwnHJCRTI19hOnBHZzYEpXd8su88QOTSo0cHDJ+MM20
0jphWGm9TH8OChcfhmsT3cK/gNty3LaGYJ/qgVpBovNIT5VaLm5CfXpGxzW1A+3h
e1Bq9icpPE/8gF25d9Ejabye202z2OfzgLN5yjdoTbck7Z9tfAVgT0kF7fAnqCbi
OhrkjY2VmXY7HeCQ8dFRgVUZU5h2Y8uB9rlbOiF9YvBQEzR1OTotf4VEADRw+F6Y
JivU1iy1TMZSq6gLZ/0j8814OtrpPC0sQ3s22QhvvHdeSr1R0uw5YWZjDg5g3mWB
OE10aMTNeylVbsN5IoimoTFFNSSyIcKxi9ljt1gQPICCnNTH/FL0xOVny4+mJzmu
cuRsqgoCH9JKUP1d+fC/oubE/jt/qIKxNse8Tx1vYcTXyjMojxe8paOYSfMaDJ/L
hHEWq9TkxVCETKSXI0j2FmX6SxCVq+Ug9KSEM+brILb5D+ZlgzBqxkvNJ7TklK3o
HAhLO4NJWDMvWO31GuFkHLurCqTMAImCSescIbCBkEO1QlffO2Y3JrV2Vp/s5zMy
DP6y5cvUag9hRwjGHwINedD/f5REncI0lKR2wyn3c3kDwkiA3VKdLvlAS/wGpsva
DNqesdvFDEq6mDlBvrzvFBjTrl+aA/95OrEKKNNyAv/POE5hMKmekjZQmn5jSQo8
FxIpk/1oQtZ5+OAZxIcyFVCgggY81N89F8EpB7pPoRWo62zEJKnnubYffzHx5i+r
/GLGJGNFEaM7ZKmYZoFS5AzSmB4n1F40GUd8P6ifR+3KTG430NgqyiuVrpO5bbEo
aUUUM8T1QNe4uOPTB8SqTxc15aeLhirWO3wS4SxiP3VCAM/x2vtJsujsh+Jk8zsL
8rplSSxNkrnuGnFBk6bz5mYGG31yoYMS5CG9CquqlcIN5ZL2fhubIC0Yn0TE1fX6
EHT4WzAm2TSqpLS0ArYYxglr2c14FaI8OfYK0uIQWseJ7ZLAKMmrRA8lnjQ1RTdI
t+W+k6ZfZWHRlV9qJGC04b11CDdUjbQ/LdZoq5aZMPiaaklUaD4DMuYbhgCvTDCn
3XLJVM+AIeeC6nFmlaxxiva/A2NrSh9Onzn0vBtdgJ+ZJbOEFw1+/ADtjY9G1PgA
kwTFTPIQJXW1xclG7xEgW0d0COJExNx9LNSsqPb/KdrrYR+9m+2V1AueZ75VCSX3
hYAPZS+Tn2kfPm7E4W6ALVp5kJc3K3HW/0+rjiEIjKmIuF/xvctkf+nMuYP0diDW
FcRk1sleryTy+80CLlk0wbIsFzM1l9+HZyaimegisc51itYEZoqpZRUPMu1dS01x
sRcgt07r0CcIon1AHk8cl5TD0Im75U7phBwLJ0Q6R4saRhhcOjDLEQ2PS6+aRqFL
yHRYBysmm4e1Mr5MF2B9zyGXdLpsBapN248OVOC8/lUHyX3OS8AFk71adc+suquu
vP69XLr5nWYxwSriWUS6NkT6NLQH/d4lgaKO2fHrtDvjcFwe/2eKaVpuuK8Fps/P
DMFBzZYqE0SiNArZ0GlWrapeBgWTgNyd0MkM7BjsRpHI5odEysD1IQsIwUFlQQje
bLPP4XckUQyLpjwYqNog+7qO/Oj4Lb7/U40K9AQ6rUJGYF9+efNsBnGttSjiBhPi
6J6IvOp8Yrq8qI/bOv8++O8ODmOcLXtyQiFAnCXVhFGU8Q5vFICctEnC36dZodwg
zq+uDeDILF0ckV026j1FEwkIY9+KIBsjU60nInKH5yBgHJEdRGRye2EoksxO5qrI
1GYg0yxWzMw5Rr3WNSE/e4NrEDwKkRIdSa4K6Eh1KQlZO3zHJ4XrpAuJTMd3LE4J
5QlbqgFbnxUbg3mRWYPTbB3+5SKhVto0QaB7AIDaqDyZSttWh15DDubdtxbUDNfV
MS0aKCosoEEms/XeAibxQPq0TuiA42u0wSS8GcvwAhLDyzGdpJ2f6qxRUv0X4NCU
rUpD14aIKHp3MTQhLX3wCtlKMEEqd94lWxQCS7KQW7bFQMg3u9reo2n+28z1ScTv
MD+Atnb+mk1p6S27bRafNEebgL8dW3ft5xG2dUCyDQKJyDHGuVJUINm5OHTodeWV
cseyCCphzP0nB8YwkKsK0ws/3wrqfZ2HXadiRHBFPQZfMsXZ6X+PlHB5taL85aH8
vZ7uiOWBPlJqzBpWC28l1R1x6EcTPlhFFXoRi2buOJchWsS14FCjIdgWrPSC5ej2
c5C2+Xcld22QS6Zjw6pgVZnWyRzX3hUFASy6FdNaJ84npHsxUFU/zW+mEFV101tG
tNxgKW6U5rEemkbKoG1NWU6+vzRJxanjno1ybEgv9QZO1BPtgDoXQ6LWIy6CsdYN
D+vELi5ooAsgiPXs8NconiZG0/bVEXRS7/k3tQ3C1VQ1A45e6YJGJtAnuMi6yFeK
KziQEnppcZ7ZX9Ss2sJW4jzkUO307ijtS+huc+am5fg65gjh/FYbC72UQoEPAxT+
mFhx7coGQc2vq20RAM4U/0zi+uXg6k+XQ50tfvkDlgFR/AMsnIWkCkFYvSdGYLlI
xthst5brqSPx0aEao3PGym06Xk3du875B+0N9zBywfMLiZX1JATnx+7UUYP4VCRY
05sVPNd71OErXVE5jNc4mAXxfiYWuTG6OoCFVr8RsM/73g3bHYqurGjVv7eC4pqp
kJyyWb6Ca8v8ffP5lt7eFS6rYlckhVAMrkpQ2+oENAyb3kZBkQMRrjWOvlqBMWwS
dKS/7TllnGKrCWpKMxnY10PLxt1X63iOLpgco1ZeGkJ2MRH1F4iDILtjKLsRltmR
vG6EmIJMwqeiNjApMhw2AEr9ZXYYdS3OO+7xx9jqmIR0iMDxk/VBXrSzgV/n58Y8
xG1+fErJh73G9hg6hmf9FPnFjS6loURXhS84GIOu4xi4gxrTSEAoR2dgckGpsDx4
fk4ie00jBEKWiXf8+Gy2ppm6YpZHWTuZH8gdPzARcXUq1gvfOBNxuOAvQjg+xqdY
ItgLmntKCUe2JBnATJq4tdFyINlwnn8H255gdL9kOCKztmwRE0nuPhGMUsxzj1Qx
rTLL84YGKR24dpHFU0qjEr3OApY0z07y7YXOfW1zfK1FFbXNO9Fjy7Su3Lr00ApJ
jfKzJbPT+AVADUmrKbNx2iYVn+FxuOJWh6qQWA4OjyAqnfse8qIOg1o7Jx3riHs/
CnVQSA6wzoFn4eM76KNApI1Dov5Bk4LlXJZJv12dJ9BJV7t9vzX59zn9QQyn3PDu
usdqovrFoMEHZAYmVrGb8kBhBM6IoaZCY/RDZlE95g2LjTFausR0sjU4clvBf1PC
rfngTW09ECr4d1FqTdLp+VKaWiJxL2fWTkuyjnzRwM7rzsIG+9b2xJuIP7ITF/xO
Gsh7dhAVPVeeJXzPb1lpy2vUyZ5XWwo+rbBtSPYxWoao/pyFmyX80ggBCKZhZFht
RvXYkBGHvwOckrFZtJoIDCguWvK0sPn45dWtRvFNXwKyRbpTrmczZxGwZ36j3oRR
HiaEetJX/IyYBMMX0bfOLTsdABAoR19za7dQ95m5NhQnswCR4wJNkBY8XCvpL5J0
OCXFM8pRsYjIXp0hQsp85qrEygql4GappnvP7LPMAf2M+/c9T1SImxMr8PCMCcjW
dYc+wyqjsUk45LsliM0XJN1nQEhKCkBOU1Q4ddm0zYpGI3SRlTg70dpg6rdLrXWy
SyF9FahGnaqCiS40oUbTcsRxjYmBnhJy2NiN4BLU7Tn9cg0fWLuBiIlOWDyCb35G
OlKNYwqhXjsZpSK04WpQm3FUjczd5kl0MqGTPeNIHIIkQ57kzAfrnU5bApqUzYVt
GgZYw11Ra1IasRgcJW2cLB7sc9pPy9WUveofn8qDZImBq++OvSD41x81/Y/ETNqA
jmOOSFVJhRPbzjChp0eHfHnpdPs2C3/70kzctx0btWpSbTd/6Zr2OfSROnXhBGz3
+N8UlkgpZ5iDaXJiEROOrN6fPglMSVaaIv/uBxhxWstErOdcgqfx8wq1h9m0EfsT
Hezb0aDD3mEecANS7zru+8qt+OqvKupBuS5H5dS63/MU3zqigWRpOXVzrr7vmycM
ccOLKDlrXPxmsKfQG/YNA+Dpmz8KnkzjRwLV8sZ6yyal9u76uakGEYFzQppkqmEN
dQls0sZ3Pyp8ZJJVy5WFzG9nlHa881GGZTFZyrbNW6/nRLc0b16K12VeWfon07QS
EaSZ7jBgBb5KF/fR8TM+1Lxk80TVANsq/ld0c0GGlNhxjpTBaGZEjprKUfqYZ5K0
VJDxsnkPHCWUQopIZZmJAWvcUsmrnj4HzzzBHgHuETidHluGPMD+exSt3iiqLvIy
wF2BPN4C2k0Yl5Lyt+fjHM9zn3ty5G7hGvNISYT6W5ajTMfM6pWFv5VMBWW+t/k6
Rl8NArBH57aqN+8vPP2/lCNa8KSCZaUzJPVVy5PzMoN30L9NdkafUQ9KW5HybK2K
Ap2mac93ctQ0ZTxsR0JAerE3Rt7SiVtEYVPBqK8JNnjdWWgPcuHnzUsEJqI+qWVJ
SSxrX8mkJtArF2hu4iF+U5YbWHgSe/i3dmO11LdpGNSKs+dZ9OoiZ6HiGGPbgb6e
gdBOrMsSUoDyrwd3zK9+VV7Dafvvpm839h4uulxcHS+t1grCx8jIFIcp4t36F181
6RTPSET7IFgYqEvZVZFBXtck3NYvpCH7NmVRXinoGin0FxMTV7ustonOSVFrIrJL
HYFDUS4KQVKlUS64BLbKun5FB4g80x2CNqpi0UFyraAzN56TSi6v4JRak2yIF81W
3fP/l6MB5u81Wd0ISPoUWG+ssOO8TfSm8p55D3CsfepWFBALDvnv0ZZWOmVRB9Wq
BrhzksOfxHJ/E27bwNVsmEPein73GnYyDGc3mpry6eYxkG++dZ2oxZp+1qAb+tFs
UuogGHyAcjAg72y/PDouldBGhKeVnhSX3/rakof1v/22avOTxIJJ4Am0cA1Sv6vH
6jUogIeApgWhhcK89iTo+ET8ubUVbozL1u8zPb3v1ijsH0ThLealr3ng9zCbh8mL
eR9ZxBTrJzX216VNgI6xJaiMyuHNVXgtN+bllwCvA+1aXH4VSGPs8xDqR+I7IbVD
AKw4D5A9/ujOahUAR15yUtU/0pKFX7oZuhFsgkeBOpp7Xd1tILUIRnQjCaISx+7Q
vhciE+54N3kaFrtt2ZvDfXTnEx7a5pr91Nsk5u/RyAHZ+275q1NEqUINsml2PqOh
Xn5+BOtCIbvsxbUjV55+6i78v8WA1Zg8R8enIaHFt89EHgWcjzHh/H2+3UXA1mp8
VgV3E5kM3ThU/dkHvxfZK83sKYlnYqLfdXXTg58uFItpznEclokoml2ERVHrJEm9
20ATi64Va1QX1er4qi1eaQ/cjJRIbDokSNHExwDtz055E0rpoS2A7GrOjkst82ay
HBeVCNhW3X1tKVJuTv4Q66jRh3ABy1sAgXXdu1yIeKRZ2vGAxhNYjcdhwxHull2L
lBCxkJDYzeoEt3i5ms1CVAHBs06ktobVKcgMqT8hdvUf2j7oEr+NktxltUpTvk+/
g0aLNocaAze4ijP3kPDrHx60mdfRfmbOnNYOh/B0IuoZ78hWCLflOKvI5+d0/J/f
zu1ydSfudjmHC9NZH6pmTunX+dx7mJLL8RyXeGvMw96fr6Vh5+v0rUo0KUfCAhE3
2bXA+3jJ/l4shqC+/LnRN9YJ5JYvWlodEqf5kSK0Fg8N9UO/yhH4/vHXJSKUeDHe
tnvVM4cvt6guvMvIY4lX+q5XjCE2Mw/+xdgc9W4Hj8nA18xvY+Sb6E8yib3MdUf5
hL7JHaz7SECBZl+QYl6uwf4dyhcAFtm/eHjl+0KGZEyCNM+1Xw66yY+j/tPdhV48
730SoDtbgGLhXg8TmSI9EZ0uFe+qtbW11WCjFe+XSy3gHy0KlLSXb4VaLGcYXMk7
3MIhQ080jxLHUzRvPELQCecy2CAtppgsFUggkJ8LHpJ5VqOumAi87dyDOOlymZWa
IqLXxd94BILcXd6gv5egmJMnzDZkg4lfMzakZHVO29kZuhk/AqhXHz8iuI+HjS2Y
s/iLHESSztR8qS284aG8PFkMGOvogcVOPuGy9WjhHWo8yyCwkcovK2gkncpfpwlH
OYabL5XwKitlAc5Oi4EZj1KRkXbEGXWXDoVFOdhIbrwN/Wl/AC9liU1lh0kmlyiR
4E+axIHWeFbE94C64ASoZ/y1JTrmdKuvhsqK5OS8NPLKJM48nG2/9DUF9yDySvnH
i81Gdhqb5+EFELBAvLUW+OZ51G55/ynStMWzpmUGRXvWFmCMrBlcYNQZ6QOtSJe5
TMtrcdT5tgBhgsANzmhb/iR5qvulKw+iw+QvK1Atvp7ENLQ7k6gDoRlcmhsguAw3
X0bt5lGC7P/G7tMKiazC3GF6NJA2SWy/UkuY3NhLYgbZJslXWnNDbeg50pv7cxk7
8fBVywNLWWasnJiU2MpbjXPIOidKJtJB6Jw2DlGUWZWPQUIAp5p6zwTmul+5FdIV
iOgpsAnSe7XOTAitKB7bpxZl6cFii8E52f/AOoPatcG0xRp9y5cGr0XsbhN9yOLB
7qrSIq8GeTKtOTK9nqafIujmHTw8jIa4F9IT/FB5cILf9QSDsUSD49AuZQRN2Ey1
aIuBtRr0kJbhN3UgY9ED78M9Dw2QXqUJbPdULOQzRnlJNps5NIwPQaKlJVL+KdSI
PiA+VY8TuUWGQSIi3QxVXL/i65sX50abeENAjsMJ+ShxSd4d9T7osUUAfe8JqzAZ
MRPAWamNYKzVPL/yuq/yeZS7ZuX3GT9si6wAtU7IGTae/rInAT7jP49h7G+TnspB
6Z8fyUVzG/y/XLnHTY1HTpMMtt0Wjk2VIId4lHAkJF7jPui3lbWAMqdxbKEkVQ/8
PHaJD/LBCQ2NlLA6Or63lH3KdnoIwbMRY+Eb+/m1SRkl8IXizpLRlyW3VxoNBuUK
y82+Q6j3lEu82mkys4NxziCoX00vgjlKqCGTJGfP47ehSuDzJc1z/stJ+R5mPTgl
eQ7F3FzoiKnjh9y9V3swrDpHif8X6Zt89QVOfhO8DJe2D5qi+0R81r9mpOz6ltG7
Cq0iE997C0ahf9utftuM4ZswG8PUClMw9r5R0jWT4Zqi3addUKW+72ywxz+MOwpL
I5xAr9Jn6nhyBs15htiLHFf05b1+eMGjj0cUtzxOajvxwXcx4XPuDwpupI1JB1+n
J7idwetEhbZQwSQK9JzWocSyAgGM6w7d5w1OSiuJ4MLRsaBRA0rOzQgd6xE3Ix7k
byYyBUkOb8tWPZcsM3EZx1GXum/yIZs+Bf6vVNyGa3CA9EcqL8C9lkJSJKTS9p8f
v5lTVfFgHWGX+LYnbsAM1mgR7To7eApgsMow7E0XGF1Eyyf/NQe+n6LcN2R6ec1l
wfT+taDZ4atTGW6dEw+LuygCYVeW6Ns14EJE8hG2J3FDg7/4eJf0f0PhPKtSu5fM
PFih9fRS6onUHo13gfXVbQvVSr4lCvdWqVAR4JG6E5VwjPdyuSljB3mefdRB+Dhl
TVFcdC+n1MLkCazHCM4uAkS0jHNeHgU8FYoxCJK/ARiUwzmds1y7YD9afVYZ8EHi
thV8Qml0/rgcONvyz/xxli4K4xjBTeeJ2CQKS5InwyG7RCcpS8+5UxhVaMZOkqu+
WMcfmjQZ2bnshh5T71W6J1nbvmcStMxr16YHGFxCha+iDUHtx8qETox8LvPFon+H
jXLxp4a4IanNaqfiZG4UQyJfy3A888gjUCi2mGbAOkP6Y+DoEufZIIs8BFYABPnZ
Rb2SwWaRFmi1RIKwNKENDwymx5850PxwTsQVYvYxjHTW2w+GVu5mWM3yJHx+0T/g
8op/YE0VH10unTKUqlMCzW8z5ksDSoxqVjwqSiJnLz7upj5syFUk/+dQeut4x2Kf
JiOgmXWi7Ih4PFOLRBMnv/XVsFhHAw3LzW6hCMh8Wc6TWloAdjKP6L43Nb1fycms
5asxwvIiJ2J2oHtl8IB0mEIef7Z2MLNoAvytiVyx+rC5vxdMQ2k/WasUAuSvKM/b
loB9p+YgTT8uKFPv5wZvaCintJrThsGifyanXZUGqWx6Q0lLjHh5adEke4ra1Yzn
fsLhyHXO06nMH9poqL3eVkahGICDJgZN3lHx/29g+6/zFhw6a0DtHK5alif+y3BM
zG+AyjkrDjTRMRSs7QDb4s/bLtu8jtj3Z61oH3ygCPeYxoo6QZcPMdtjuBrn1qLe
8V30NF11OuY5RLzp28Rj2okquI45upM/Nv5vtOWa3uxlqaGGCeWZZg//ovW/8Oro
2sZzPsAJindNDb42Kz5kGPeuNSHWEs8mIvYSAeU/CL/lh6oOSlQl+gKcerHSCi+n
nLnlNn/CsoDtraHsmGbS6xzx8r80Z7VWQl+RauV2t38C3NBtAgPRpjIwu9EDdNvy
cg+5L2rveCCr+nLbyKY52FwhLVZJJjbU65hiVt0zq1h0n8dPTW2KAMnyl3rxC823
9gGEZ7VGXOaGkhyHaFH6jTz3UvBRVk9B6f4k68yMTFoqSvZJ+FT7xwuOINV+eaBg
9xQ5G1znWpNyvjP3TtBakbTtTc57POUQtSAMaoxncRUcw7mrtwLWBbxLY/jhGaWk
ejWQ/TFPJJo0bqgSpgL+CV/8zMUP35JB+JJQlrVriIXJNmKdmYlk1EYArTkiuLqN
vQlHOprrOHmMOfZ1dr2vK5p4I1XZgqeWNcrAP22YwntMEhXGZa0Zbp+T/xDHxlwh
Y2tBuwK4njFvxqDwRRP6nLH5R+jkWeasZbKN6vGdqMcYZHugU2o3G481A+h0XigI
sKpIHXbK2NsS+bzcGBF7B0hAcWhO3g19cr54LGbW1F47+fIj6VHxefhIUCXGkxEf
R9ozttgD1tYsS5mPbNkggOcUGW+KwdlMq/GUYn1WxcarfD/YLgLA31as7GUGVVkW
9knsbVwgWKs55oWYxOnlOwbdU+MjNDEvDw+DWfy/0KWut7auAuvcB/j/nR+9HpJl
e2NxtROlHAaR9+atDCY1S0cnZnYBzjSM3IU/QmPlGiL4nli2B17HicCa6k+p7CEh
hfedR+/I/xE/lZ9e5bRCNYyBQ+oWeLABb0Gy9xpfd+1Ivo/34Bs0qXx05ED+Su8m
wauxCiActUO0v+pfcey7Gki9NOOYhXhg2cXHdM2Jg5u2WdJ4xGm2kw/3Ivutnplg
OGGU0I1sEPzXiJxgEycBuq4cj4x4Y/aZAEW5kcndP9kQ0EWXAH3l165OdfAw9Y8O
7/Tp4GaXUsQe4+V52D8DxwSvFCvqXXQM2Lp2J96WWcLczKN/ztykwU8D76shmsc2
/3BRy9rgPuVSWUm+1havZQKCVBuugWDfZhStpJnNL0adw1ld1pz7SLQPKO6shQnc
tTYdl2mu/d5nXtn+uXYr3vNMH/5iO2zalZeiJvqDQyEzmC7RiPDnAXlBCVGRtuu+
Suc3Q5mK9jmxYblWtuWhNJO9cFrBvLoESfWM1YSGhfpThWuf+Sf536UwtTpqInld
7eTZIi+sjEqSDkr8EuofAMkZVgKI8xmF524ompweSESJSzoS8l0QdA1A/3lIA6cd
53ASBJMUatUgS7fb1rUwzlmMWvGct2k9joUhFKrejZeOVLZzFYoIpbiImTdg9gQD
coPHgxtLeEsRR5Qro+9y4XVcr7N443D0TbytLxfAw2hUR2+039RYP4aavnuY63Sg
NgdRx7BbOO33sBfWfnYst5mKI71WTePL/cEEuDj18kEMueQgviGAh997w7w2MeV+
/2p/ihArphnHIG42eexYVVh4W1j3BioH5JJ+hxCRn+Oclg+3ht6EGonuwyvR/cv3
LJbqffNnHJGwvEWUMfH3w+bvwOwYnWmn7biGjXUGcHQ5BGwf/cyYbJyliPpYV2N4
eXaMa5WwuhZLK7jVsl0HT/zAvlQt1q1xWdCxCJXPD8ql3dYRciyh4ufWzJvMjCOL
binoloz6g4qu7cGl40mtuZQAM+5lDkrmG7HjCJoxMX4smr47iF6GaiMc/V75udIE
NupwtMH04tlFGfrB1/0Ujt7Dyr27Tjhk/BULuaZLcUaH5dWTxsTWU54XHS+oQuyC
+6SwdnzkUmbxll+rb+1WdbLBs3QbQulkNamnwnuSrsDbQ49p9FRrqlreKvhOvK4t
LH9pRLkzEIEyTvKbhzNzdh0k/Gu6HvK0WOtu7Ui5A7Y+cnF/IYPtFEpSX9FEZAxe
8WWo14/phQ0exT5MbvwB0OI9U4/taLFLyCKyUu8CFh3O5VOyj5omPHbf/WhNEA4I
h/n0hoKhehSC/Bmo62+zjhDReQ4S4WKTGMWaT6FG7UQMsjpuoY9ObJ/Den8jPetx
6ByQ1/K+lNWuljUmywNet4qltRgONvbNqAjzmXpgKJlqbP7prn/LFX4stVQSe8T9
mOmuGtrwDAqRMluOedCuRcSS7tuu6+skCtY5B0nTsF4s/o1nNY9bfFtMVMdTAHaV
tJtBkzrxtvZcq7Z0xxveHowzc9sBrqSayAXy5jBxYQJUqtPaR98zYXuW/hgM/7GU
3A38iGzSLc4QDjARvBgRu/Ncl3ShYWeC9l8Y2N4P7/gqUP0yJ/BKuL0QLwv3Fz+l
tJjjF71IzsqkwhKH/R+FyEAdioPUjeOFYeVb9n60JhGEhlQS6x5dfn2AL++4q+EE
e8RVPkvC/HyjBtBSI71gGgSIK43J2jOckU63maoP0xw/rwTjGSAFi4nOrK8/uRiY
KRvivq5Zs3y1CXiDhnwAzhIbyfNWUJTlEqZckXSgHA3Pf060FQ8/MkmvNj8G3nGp
2A8ks1o/x2RqfzrR3MGkNPHhyyeZYwzRaYEykEbphezVPizQ8RsHa5qmn9MvEVe/
DyDeQzjvh9hS1kj/COSbALDBkGpHjWFjtoTamqUrrWe87/PYzNZzRzltMK9u8wp9
2p9qrkZ4lQBm29BrVt0PSjRw6o82OgA8MpcspOFOt46CrOenb7hgPmB6IztN+x+K
zb6OG/L2R2WZxkwa3zzGm+szwCTmeyVzMmNUpJkCg/sLsjecTBvHIR8ezU8pcVBg
9heUeje2HxRt0s8rKsgvBRbTyCo6W0f3a76IgZmtS/JKNrHa2apuiAl7aJ9hv+33
dVk0y/Er3ewG7V7W7pJqTo6V+b+2otMcE6SzM019GdS/UGZX0GZI34I0u3mwFK56
PEz0RUJH+3Sz4ZTX7i2fxILBfgQCHdIIhNMph5peYBu6bXLCfvJllirZm4btLDlG
na9exYkIxmOt6PGzwPaeCRH1rp8Aa+N7+tvTPMIsFLBc4R62PDblvdoxvO50apen
6ifMSsPTKdwmlu5Xz92b2qPWhjXr/Dq79xjtXHK4MRj4KMalQvQt54MwxK05EP3c
k0U5N4PmP1jpo39xiZtV/hQCrEtwC/HAS9sgfMh2zsQmyDHIjkFRDQgVqSuYt8Zg
KaUAXqtLBJl0LrgRuJECjS2Ed4xvkaFplxU+NPMIWA6rMmNKvqKpaoiwwGcDdLzv
miGvck7PGDeQrZ7Cs5OEAq64BKjvhSxJrN2zdwOgmU2akRqvyDkEW2H7KFtsmZ56
1h98kzRFn5fNyJs+uU1SgSabrJOW5p83FgMAGvUoALjsdoTtdL8m0iW/NNVvUkLN
eZsYYWYahV/9KMr7q3EmgxplhmtvDDrBozYUqHwRtsBQekTmVY5LeU7pt6ysqgHI
xkNDvZKCunCXqkh6MTrRSDA4sf1L2hDNMebzU2+MxiTZnI+lDdzdmLdfHLBweoQr
3kIjXF5TyQo/NTWvgiA5bDqsOMxBex0EVJHUj02sN2p0wlu5oMdP8usx1nPZpBeW
h6eaENiTsNk9TvkV+wfuU/3ql1mq7z3zsq6R41mhB83fG8mV/ztY3/znNZK01VYl
r6WOpIcAzpd2oiao1MNps1HFFG16EuzIAiaEW5K3v1E3miWwtPsjSnPH8iims0Oh
2viv7k7EOVMSuj3hC2ttFkElAJaDe/sWrxMieAMgBCNKUrErBkdFuaGauslJGxNA
wcKbafYnN/OmgHZix3WJ/VMtY/agvOMcT7TccQ9Owkz6MPTsTq10ntUX+0K3CNBl
NcHD/03tZQqKUo4sHgv1WBJMwdHGz77TAMhomVaIkaQqRrJA/Fdbmnvqd2QJq1fM
H2wTVyd7u5nO7jOiKtz65g7WQWnikSfMJns1/B1wIu6A2b3p/1EvpDPJ+xSzkp2t
elqswWxfZga2HOxU9N+wuOb3Uob0y0n58ezGwNBXgkm5W+TK1BKzNnUIVvjuQX6p
hPJlbZXNXYXUlSptWC78V73F0ZtrqZ0lhSk0nLtgBT+2badKcN/H2gC9GF0Os3Ck
ZMPKkdXBu7IMF7BbFsp31SpKQv6w2xnw/9iK/1pHIsdHsVe+ZCqeQAN//dZVUVRN
AzGJijivFWlSr32ZS2V/lwr8Mq5VP5md6W8RaaQsbkQ6IJqgxOCU2ZqKmV6VKBn3
I1fKTrJWSnNry4lhRL9RbbQ13otsSyL07jvRHS/1AQrxDRmVh990xBOpGvdsv8Hk
+es3hjojvzaCHwdtaWD/A3mtHD9QPdd/QGO2qcxr4SxHoLICvN6QzgdfoE0lb2kQ
gv8vVr927qTcHHFM/mw13yTkP9Vp93wTu6yvXnWdMqGev4fuQPHB0/2IZmu3JfeY
MBBaKvMjWuSunRxfkl9h1oXegk5otDrNjTvSJU/wOhAW508PJkrAKe4x7COS4Ccd
ntudtzIbdGu8sLCx1UE+nyejMgNLYL4jMJxtyQE5xt/BCXwtS1dcpuU1FR1bEfq6
nZc+banh5TSrGH7Uz+nuk5g60+7TMrq5CiOQCKG99SxtSQwcDPzCcWwKFZ4IKIvH
Hf/jTvTFFCGJfQ+2aZ7zZ6+72YDfssxpwCajWvua5UNlhFBISoxvmKL/26+hunb+
ZO3i949MIphaN5A4iDZ9u4VZQcJbeCe0s50hfZ6Eh3EPV0NGcHgFRC6vkZELNQ2H
2Tt+xQpFUXU/zJy03I25zDh9kqW5fYn+ZQlllovGZNo9JHzYP4DhqmJDKyq3wfDx
bFhfqToKoBYyF2gvWkvS7YQ7+/BDQ7LWHCRQ3u16UEl/GCIELSjeAfJMt4VZLYdN
2UkV78svkHdsZVtL6OnK6yhCZKRB3r6v2ittcn7f2rUsSYMRxofoBQyjJLfcZqoE
2IWkdheoSXvqRRfYgTYokgNTCmkSmk86hHhP//j5qN447gVOhtyIecpRH5qm1E9y
8gB+mNF/V2t8+ehQcHP0SVDdDrC0v/tux5L884aTmzvXKIl3DMwlRUw6VkArGOiC
HlL7pwyzp0XLBns05WER2VS6UuCvXGjMHTYeVAnsnpEdR2+l/qYyOqDd457+zNxR
yJcwBoSKRybOCmX9Wx6GXRmGbp0hTJZ0g7YZjS/K8ffYvC4Xz5dzKhr4tMjy1qth
qcNFDMzyU6y6xolw2DGAl+J/cjfePcUDzRJiHD/el6tpZu5pxjVLZwRLtkQ9mfVo
kx7NcT+fhKTjBJJDPIl5Xoku3qU3gskw1YmdKzn36h2J2rsk38K+5UWDH87nkRfj
Tsr+RJGn2qXkDn2skxr8IERYekLlleUpwfPcFtef5JLKdwSv2fKXvjukB/c0CuKi
cbTsJUR5GcQf8OFzyH4vNv0xOBjPE5iIwrsDTB3SbWvmXDpSkxAsAy20fArUF5wr
JP5wSdCIVU+xHb3WJNJjPLGTiFWIZjVFE08fMKia4cVxStoiMz1bNF5pB8Ga/nPQ
WPKmwMSkOpCbj8QQdloO0Uf/bnGbxLNn9yBSEUDt5EgaQeFS1QV22auBtNPlKwoA
4lS4KSuoJUmG99oaNxQgVpiM+KutpdJt+oBjSlbl4iIAJCWELuYUI0uuc67SPqw9
GIazyzEcusAcdcvbx038LCWd3rgPUqknNZAKTQl9hMmXvVJKNyX54EcJJoJTtwxu
1RfpuqauB3Ag1A1XRSIufkoFBZFaqBbU2Ez3RQgWH620WcmTQhw/yRbUIfhtQCAe
3V1j5vZR5nyyABAuEUSsNgk1B4P3y2vtago4y260TYYIjro8B/Z6tDGFjWEYQaBj
94EcMLTBErXXdsw4Xb4ZPQviXSBlZbTMyQOR2SKUEKoIHewDpUmJ89Jjn53f3mKS
fUuZr3Wg9cckMCkgkuvVYs1+zeVlSD7F+yhXpJtn6J9TfeqbrRWfQ0Rp1gse5EQV
Do/Z/z6Ex42X4VvF1MtdlfghyO+8QZmiycQYCB5uP3rjCGvdRIlkMJrPOwme0fbr
AJcoAr2mPYdRrJMbAA47tdO2yaPsge2YpzXbnKazR1kAfDZoNv5efutlFVR0xrpq
e69snqq4/2TyF5Av9YDZGYCVfJKVnf39c6t4c+1XcB1fdikBLSBTskPskBUPnQMN
uEmMZHVZgxtPtjs6tsnQ7qA0zds+3wVuYc9tUnACEV3u//lMrk0ow76wpWlNn3SR
TSZznFDbS5J2ja2doT5/bj+Q0wvzU4282TvVrZ8juE2d+JfjjvW8sCU12MAaX0V+
9lg9eohtCmK9iqqJktF3rs5mDYEB4dtMkvWmKgEHEGh+fAX1OtmbV6ujuEstZubz
iC39PnClFlyZTMehSNvz3iot4D1neZM7XIqPO4cGBSfs92aEVkqj7SRtW+sWbf6r
E4HOjZm92nIdJOQQ3ujb3onyDIJ6+AyebwlXqD/mbrao5/OblfaDeq/eSIT//s3w
KBvpIVAV8ali6Wwm/y9CqSv6rXHDwA9MRDqTsot1GeqVCtwItAk6st/sVVN4ZBCJ
FFg5ffaXrsQK46h2GpdeBQoZqbRGf5HunBh2sm43aP7bB8uqwroRAXI32Ok1fllH
lDdMcn0N+FIEvhKZWmQJ0QRbIvt0cJJfvospWXgKn5IuCz6+MIfDHhg2njlqBBJc
Yln4NFtXtvKuV0BLBBbfOVowdYxwZAU9RWtCdr4P6Ot+0JYg8rZ3UMZkXBQB/cuu
ql2A4zmFN+1CwHh0VZxAKOl4qpV18nYR2IMou+JIK0V4N0PFOBUGmeidnxd7krDe
yYMpna+ChRyVKnIjQDOpJ1cvPGSRiG3C6y+nVLBXGilQb5dLK4j2nWEmxmirA/Sv
FRbbvVkktxp4d3MRAEFgFBCafuKEBL3KwH7qOZ0gNZJ28HPa7QipSVDmoFtBXj/L
GbMeAI22QROCzAHuOKBB+DE11Iz6P303gCHV3ADwqzSXeuFiBGzeF3jRW3LOj32f
AZoB4rQDozwbS0Yj2T/Ry3kPY/dT+OvjvufqzWgEdWtRwPZ4pjZLhFSHofd+MGAs
119y1WGYxpBHP5iDq/TgPVkyt7PQ+HSAACRQjYJKmkkQRHn8Lq9S5wnOtP1KR47J
FTwgahZXZ9+UaK34PII99/+k52ahihiLD9VyIIcjycLHkdh9zlokTJX8GiGGRNNi
47mgxjhWyVya4KE8b35od6SKH5u6nKiKf+6b/55mEASyveLtyuVwxsV1gL91ivaR
ICb7Gv/ARPEz+lTbifoqUtGrta+bfe8AIU8W8Qk+MgvEyRwXK7wR/p3vdOLlq6Y4
n4eFsfrGOZZHgrZ1g6f04bKuk+IzVG8FHLWlZC0B5IbYkKdEDVmPcP9wliYRgoyG
RH9yIGVCNJ4Jpueb0YaYFCdo5GsEY8Mq/lfYjGN2AeAw//gj4Jev/KlrB+uuDZC8
jl0QEwdyHzVoq8RwFhdWbnvO+nsFHVn23n8WhavosLxU42JzqKITSNf28yz0QzK4
C6yhuFa0jYmnCGq/93Lg/L+gsEvfv2FhjLIR4fQph7tqEAN0DsBPFNZ8nHch9wKN
TFrYsZ/u/dW4GI7lQacFotCDExTQCaM/rd58DMVLNwgiXIURwYX/LRnA8drtBuSH
fByUIEp6FUaLy2LVGKOyZ2bAShLYzkxcO/JD9Bh6VaEag09c5kNJcHy1N2SXfJ0u
IO2fZXaiFlZiBe0NFYDlMTqBzamGg0JA2v4uyXM/FoRXYFiFd6VkWMmCSgfDW1Nv
+fByHdA16/5sBce9S3OtiGz9YyKdwdw8SmDhDSiWbxwCFiOqBJaOAsT4+iAWDHPf
rjmlCmF/fqRUM158/h3M3DeRsHU4GicBUsdlXd/NdFrvvhymoNiJH5VuxdBmtCQC
dtmbXz/AHhNWeP/c775WFOtKqyY8AOQdGIMGlntUGVFPpF5ZUu3Ti4vxppQBDaOF
5PhsxK2uBOWD4kHAnr+nDftmdP7+g0rjzF0uGdPz9fUtKiR9tTjWTQZTy+9uSbgd
oxH7AdbQ/JJ08XdWk6SAAXe/1OXfvAJwsnhu63qiUqVjLTh0fhgsRTxQToD94WT8
fOd0uST5i3V/YXlBEyigPMGmJr9N1+E3qzbJc/7bTkgstvIwkjnvvjShwDDnYEx9
Lao6S+1AKkazBFn3mPic9wQ7QZgEH28hVQ6WcWYyDtMOd/jfj27SRJXLHTLRPQqe
W/ZA8/wjA29Eeio29OfP+JMyvmSc0JF5B7jX2fV3/bsRE1hz4ItHpT/OrGToRPsC
oXmcx79sRfAft0sRAATua9kMWKUW/Um975E1nHWM+ke3Z9ZpPMkHnCw3Njay+Brm
Afg1QUv+2WQnYU5H6wZCKXAvUJCamXerwAgD2GhmHjnjx32Sp5rtblJP907GLlTO
R5rhi0HfmUqkWZQCwiePYAt72OS43TgHFLG3n1f6RPUtHgRqpmJfjvr44dlrod+j
MPLD0jBlbiabW68tTcSO4ZGb+eKjpCSo4vKldjZ4KTuaxyiV0FsUuo4HPo6RE1Jt
XIY1j3mYjuh9tocBrJCNlyWAt5jEJ0XtT9YK1EiM10GcDfjLV97xDNLhf+BnjGSe
TmoKJtDJCI0M+jAWk5Fhwojj0+NoX218uQWcvqHSnqsD5bHTXXXaJJ16Rx+xxwys
bh7n6J6xVZIQbb4wX6CCQsK6qgouu1iFGpSS9JYLfhmhbQDF694kNzyzlM26HNth
JBBnD8OQkxjHTfgds9ZtKigTkIf96/JTnD1KxPLC/TZAtCA+wJqLaGOCIgInOcxc
2SLEf2M2yJlvBzQAHTSnJFrpIZl5uhzoHeLGY99nOq56ElFdUBbTXmAj3q+4I7Ku
kakdNr9WYmWfhk/Bo12sA+75vKZmNYF4NrmdH2xXUHQPKPsAVfEOGroBbZ+g1LI0
NPw4MRj6lkzT2NfKYvSByx1w72EYHQzG8IsgbW34KkyKq0erkqkuJrLNpEFjxTq6
8O3rVnGAU64pKEwSL5CeXVUXNJHt79P6WJX6D+Y4F1lGplT1DP3vSdHsQ5+jDBXy
G2Q/oLb3lxw0MnhFzMXITSlxz89O1ITzauhBB4X7Tytw9E06QZUjABmGgeQislAI
vTTv+IToKxz49bMAZtafG6BOaoSbz7NRpX/LAFykxGxpWreUVLFGAVH61xoNHttB
n9USNLE6ymF2mVHiAB70SWXnSkAmeXGmXYdr05j/XrztJ21HvMVdNgrT/5azV0Qd
JzeMZA8jIQCQaL2fHH51442tWRh3Pi8N2T8yKkpDNeZkV8rwBK9nJkCXKfk8ku+L
6K1A1bgDi9MC558O0w/grLs3atbXWKUDaQDnb03gW8rLO583Z9H1DLHIjEKAT+NI
8iJf+v5Gvrd5v/E+FYdqbygPoH0INKb4bZvp7E1U2WqD1lk3YxrY0xPPyDCvsYnz
58NQ+UVtPyd6Mk6xbAdbET+fhzTCNYD7E3twVjArXGtReEyVfuOrn8swIFh6nSyZ
u+61Z94CAnVmJXM9Jcsyr6lGYc7+cZbNEhWsUUAPkTXvPibs496A3tvVq/3R7dYp
6i9yXgm97DMfUp8IaP+Gob7plWRsH/UBMgSnznjH6A/g5/FE9kYbWrU/H4R6/0kk
AHzgrglHpMkX728BO90tYga+8eWdvv8yoVj1R45s/MrX4InZVR775xo6g/blcjev
WxfHNvrg+vlh/LSlodaOOlX04uXTlyWdwDK8XOvEZFZEe0N55uW3BS5IJK9wWyuw
5BCmB27mKjEpmqWNrY6Mhydb0sPW4BMB/xgAEEznzadVBOJnXmShhCP9xbcJxDGz
IMco16qikdTfqAiEmgDdZ5QYheksDCx6g3C0rwR6+teCOeQPnotvnKiCuT8iLTc/
cBItmrFiSm1YkoulWQ+JlKTBs1xqYRmh6eCUiuxmtqjMou5sLDaC27awNNrqkXYQ
q6ELeKE9lHAXmYsJ0ty5/mAUxiP3l5JevLUN7c3VotccNQ0hYIxWFlbGeQM36w6U
H/NHuTpZpDt2RkcPD8fcHirPhXdKfftnpY21dfZSoyGviCfSwF7JG4LMthpqWU0T
obEuEF7t2UqYg5ADVoC5pf1w0Kji8xeo5eTwbBpiZoGP80qEgAuv8k2ex//qyt6O
kVWZohLlCpoIeQHnST3KIpxh26tdm4d7bqgQQhe4We/NQVtEMxDvqoTkm8jbsKWx
6VXKYpvceREetrpNP6TtzAFaMlxUP4Af7X1TkS5ttLKQBOdF0uAtbqbn2RgFl145
2KRlPTHb+QiwBoBsiIrt/VW3YZYnPNHaDHWdpRUdEGTKZOkg0q18FKy6rctZ1Rsj
ONqeun9ju9FlrZRALMqRbx0kTjzNp29wtynJhYORzYyRgRE+wkkrgdicOFCDljnX
ryQourZ91lm4F2QnWd93RIE0ODNFETYvwEAtHvedtk+m/CrU1bmTti0mpUKgBbVd
FHF4IEuBBmIdbMjfHQnCXE4Z9yAUAOnE0G8b7aEVWlBv5rmu1A4JHcXPhGPfuD6G
/Pd6tNWXcJjqdxQwl3Fwoh0mwpucDaOALGANqi9S1De4/Va3bdyCoXW76HbroYQ8
StRqvjR/XwtqrYqxSmZ5rf4csc7+INYoo5XvRB4uK9+tdyYawNlIyO8Nf8OBGdmT
/3p0YAJgRllbKK7f5QALd/JMhLHZ1umjywShuGSikxSzV87hZTg/LBJepNlHMWHX
UN6ltViPrN6YDtHucK9FLLBB4mJ70rRz2RZwb5mKGXZCPL66n8SfDmXCd2yk0raY
jj4CASi9BQCsUHVX+cVoalP8XKxeQwD3xo8qvQ8MqKZdOlBVc5nNWCau5z32tKWm
WshtSs7g7ZR1bgMKrPbmnpcbSxruf0/4qznchBZ7+5j7AoDcIvB43gYaS4Ux5NTK
hIoUsN3IaqKHlILxpCPFQfvP3jtlVRQEUzKnnxZECk3If6R+Vl5e8hIBsGwvuso3
L5f6zpkHJkEEb+5RbxnDkj7kfp9fd5UlnxaOz3n65QHXqVYaR4LoMlWmtnM6uGG6
m37Z1uae0GVqiQ3jbSl99/Uz5S93W4vfv/B7eIVIeY4mv8fOBPPrTA1wdwwmCpyA
qPkg/+N7tMIvvT4xhZ1lX1aI1bWszLYrRdGzhAQ9PW+rTikmvuO+bqXaOyweEiLx
44Xby+RJVieQNOb/3J28Z6dLfohGkVPCzVjxAyzkaAJh/bWC+Nsz6nMPqIPt3bPC
om9i1sSnY64LTxFc+OiOPaQHvoi/1g0d0+BYw5an7sVcZUZiOWcMRGMz7IpGlgsh
KmgBnv/IdwKUPXo3emMZ53oqjLcTbwYSVT5YbsIyVnytwujORhnNNv2HSBLf5C93
M0WhOuy+QoNzFqiwnP5NEXdNTAxhm9RApoOy5v33hvI+TrMDhcfRiGkJG3d0Gr9b
mpwatp4I4za1BfkwrWTPOqyCxDOk24DxsPRQKRIswTHBvRs3t2gpnzz6uExGx2Hc
LGqTjdJA4EB0dDACCYCEI9AT3N+5cjyZ39lp8fGc2rG8wn8dobVy/RuQDaNkdcIo
+4sVyHtFuToMlSjRw2NB3Q8VCpV9PqlNsQnS0yJa6Zrru+eq13B7zSIDgBwwdRX4
5iHOYkeFsotz5Wb9s+G3l18BVYkIeObR+gmxCr+n4tNHpmwSt+v3IExu+24iSHoj
k6vbJI5y1TKwzQUx5j2jE/Is3VPOAWG29o7g+vSrLxBy4HI0sPApgI7QScRYn6qt
wkQjF9/S7mhn9kXA3vHjvnlyMd53M6jVqX2rNVsnh6q7CTqVOplrFlSIX98MW+qc
iYAk5xvtQGyLYToIpZrdwM81RJyYJGD7JxNG81u2IKc7ZKxIL4igFgLYrlFXRIIm
mt/OJoJdz1f03Y4N/YI58UzZzFEe+i5gQjZ++nx4ZsYmerXUfTTx0G7KgBeFob7v
zqJyc3UUYTVdUyJGVL+2ovihFHh6twQ3+jvlsoMwgPbKon4Z+VWcqyTsdFcVhrwg
yVAqtECPnZWsnwPEdJcvpuD3UwzSL7kOXvOjO0EApXlMuxKGhn9o29bNtkQwMB9r
lqgZsNjBVJn9Wc7Q5QCqGczT+uX35ykkQ9LWb9CFlT+FeSN9vCBKa4WqFD3hjRPR
iSESsxXWhOc9V+jyoIqGkUmNZcLs4E0hk5w517zsVq123ebUgCYApLFgNPfLdseq
VwNWvOBb69Yp/ZJXnDxEqQY7Qam+BwEC6PRvn0xPLfr2cLhY5xlvMAWfGhHLmMaj
thcnQIBtXU2UbAXThLQC7fz5MnQ4ONthLx+w2NeKYyQnJ+TNI6dEujOynEnBc9br
embkWTkXo6uXFWmlk7qxJz69F1Ic+A4Tb/IUkpgGXhtrIIePird78S4JjVQ6nMBP
r1QpwC0/MTv3d4tayKj45AXqccitKjWX4VVDa3k1ZkJMRo3O51RVjA8e44EE4Kgm
mTiu5HhgbqoPohL5h4de/lb2yUwQNsutmAUv3jkkQAYq+vSSJnEP5/Kzp8Xle3Qz
KX5B3Sdalq9svnztHFOOg2fEyzG+ICvrRX13B+WaPmvfqes2SQx5gKBGtB/5uI/P
xMjaDXiTfoOSCcjX/A7rH7nXVzkvnwsq6eK6lEM+XvxQZFWN6mlhClDmqsdbQP+h
xmWp2utpmclP+7ShPIEpAeUrl+gJCGNOwRNUriSEhHesve25taSCCL78akLoNvij
6IOWWYza4eCHxryGd6SCy6YSnAPvSaKfOYmgndPhjfBgs6f30keXfb+xVDHh4kF6
mwDRe5WzyCiyZ8nTaJSYTVC/jK+NtIgG8BHlr04QAm5khapx5KIhLNaNgnA9nz06
rfN+dp2VvEPcrDiQTVokdkA9I9AGVC51L0gWneF2ZJYcjnHhBmG7I47487tZ0r4o
XtaOiB83I7mEELdYvCQTPnTPOpxojcKEmDp94hYZ1/QWhvqZNhTO68XtzUFyMUmx
xBjU89jtbUgUdxlOCO/bHPhi0X+Zka0lgJOe2CN3mHUnfj/vCsVvmXEsqmfAf+pT
vMYccFt/mjWuGTmZdm4/Bs6Cbq/iCz4HMRiPMhqQW25ZTyK/QRve3xt1wwfgDiCb
46znFo4+JVwq1n1A2HEhEAA/6+dDaVnDfS9DVLJVfhAvWaxBLczZ45aAeQ6aMCoH
pbTPB5d7LWN8TGrtUQp4I7bHZoMZ2MzVYB7eN9Iv4snfQl089QvOaXQbo9bmphYZ
nj8WGt8Is1tI/kO7amwYHyR0V4EwbmhSg5Ny4fZEBsk9vyrtjXFPyyRlfcD/uiJ1
xVatG9bX5Zw4jMbZbroEYiMPeed06tHZtwRBWjbJoR99xjAH34bfBMj9+macwuj2
AJVjR38AYVJVDU0+Sv8W0LjaERHDW2prBuKnclgshRpxWSRLU+yR7K6vDL4R6pK2
mYahODjpp5vPkzFkyHSvgkox2dF53fz0pQoHDWABhrkofVRK7kBC1BbnRMNYdF63
cuZMNelEUTifXTpLoWt5Z/MK9YNCuPDM7QmvoMQTb39GQpxTMj8GTd9yAOb3qpZa
fR6LhwBStEg9eApKtqB4WE9JIqbEvwrk37Mw3kq8tpydmXXDnsXCvWUqU1hfkK48
CXp0Ey5rXvgkKY4dxInC+P/e6k4FCHWlRhwd5rqBab7huZhP1XFfuOZfRPJyLBva
QnFPuBcwoiGlsYaYz/uxKn8H439yJxNliQn8Td6sDblfuKQpH0mlrxlIKNYhUqH3
HE/HQbx0iBbt2LiriDEte60qsXWugEbRpddRHQ6qzUBgPdeHIL/lquFvMtLW1btB
nds1Y6LPh/GtYu4mDBJUd2A0gH9AH3q8XIUieWEutQNudXyFCzm9xboeV2CSZYsL
IKD99Oj9rMEQY4+n3f/dK2TV+kXgwb9zlWygTCYvvcdKMmRxnJAOQUcYiECWf6Xb
SztW1CKdrR2MYhddUBwcO3JEERlwuLlACMXTdDzoS5JunJeXsCK1EeWJf/O5JWTG
staFxCZa09sWkWyotk3Zw0Th4r/DBrLQiDGeeJ5pXFBAYSfl/nyk55SUpu+vXCpY
a5pKZzpBBarHpskcy5TYp79BFw2gL/bwE5OnsPhSyaYv4sGrQxwWp3jDKfiRaLdV
W592EfPjAKWS7ZpSAxARPwi68Qzbw/PfZ9LT+LSkstLbJ5gGvrTavKLRXwBOJ/NC
BlR6Pd9xUVm4Im01WEeETF8/ApVFQZzhPf8UwUhIuboMnQ9RZB4Lc5WtC4mj79Yw
BBGL64He7EuWUL9iwvgbDbcgPphE4ReR/lU2ZSXE3xMBIs7FY0k/CjTK6KSRK7n5
RlI865UwUdnNaMSWZXuuSmfRG7I4/PPzq6iMeLGVPcJX4zsbgWlJKW5pH9GJMJIH
TCnGMTpLu6AgpfVfgEJ06ArLPzPMmI/di3SNQK+92aNvdayWwiZMRguZcBzYbBWf
rwzw5H+AYrCpC9YMcnhaOKer7lMnarE3ZQ+nilVm3WhV5pesevY/evBHQBEJ221U
jb4+wc7RGM/pC1x3Pp1cSzwFyGrRJS9jkXSt2Lk2seWZRayH6Tc0sr0H6rCs6YV0
kyBfUQyUv6Bd040yTrn9TRU7rQXOZCDmMTtSsRtj1L1wKquDZKahq64/rZ22Wjb/
Pav8w6lDadUed0ANlgnpNjhkDdOvBvqAeRFL11/b7VbWjUOUWb9S71dwhltEeAis
ZKPb/Ravv+OhSi7lvDB2NG1/Uh08Vwjv8fUNRMoPCMV9k29LKIfUGF/V1FnTkIQe
+PwTtyE8QUVcseoa7YiDwRhoQvEyPmk05gLGcssWuzZRGou2R09F3f/IGODYkzHc
DADqetwluUdFCoZRx1B/nczVhnuvJSBcXV2nNv63wrHLtidPG0vW8lRH458RFNUB
qIhCRIupCPxVaZmzeW+9aNHqOiQUQiAiGrNwMXxSumzh6zVvd8uqJ4Z/dHh+JgGf
MNNDDwNTngF6mAIb7gZXMSswnkQ4TdGwfgJTbfCT0XsrehaPMO4iGHqVD70r5rdr
QWwQQ9v7eMhiLkiBrC6NLEgd678jToNDYxlgG8tgijgOLVyKpwKIH4gT1SSlGXpH
RDD65RMl0rdHrcof/k8MhoFPtvEJ59xwb9rvPZoR+Xi/Y1gs4D/ZF3YArz10cxgm
IB95L0VMrmtbeN4Gaftcn2d5Ke6mQy1xMjv8vJgQvQR9vXssTT7c8kvATH77Kxw0
7mHt4CDpqt6b3Gd34HuDMYs4fLaaaTOSDBjYsIk1pV5R1CqR+24CgHhr/nP7Q+uh
qa1u580WqAt6MbEkLVpbdeWPFyIv/7d5wuYZMbNuwrW3k5aQYFNEHgq9zALxpVC5
gJLOsHRQK9CVb8NzJ/mVi/wDHr3FdgprOSBREV3dnvDnWOVeT9YX6ALfz95Gu/b6
IBGdXLUGKFmQVTcc2dOyEDQTFY8KyZe5nzeZ/acvfzsQM8LT+jlGXBYvp6QRJD9/
ggZ9mty9sASrutSV2GFvdcuShYrV7ybDNyrrIk2wivDowdK3gIP7r5nbW7Bn4gME
QoN0ytvsxXLHSPAOCaRKAiR3Wl9KC+BN9/eHyDVPyNKF5ODftbkIsmAP5ZkyPn5i
a2iJ6cqSxIEASviShGAb4G0n0TZx6VbHsqPE1y9q+63FvIBa5F+pXjqllUaSRqIk
A6/Y3cR3GVXLP2Irt2fNRmtQy7kWJOJcD85JSv/c6rIa5bXw9Gdj8lbE3kYTzfII
tw9nPmGcP2j1Qb4PTshYtFvoyrRqZCci3MpswWT6uPcYJwC/YvgjcrXjZRwQ+axQ
fVtnFgquZeOM7bkeiajAwmYbinbUbrX/odT2Qx2Y2e5cua6fEyb/CC9BKYjjLBtq
1neFGGyDfp2s83tpoGUtnP7fXU5Akbab7qqZp7N9+eoK7F4nFLdfPZaJn6ugezHR
PEGV9OADhYtR8UQbVGZEq3PaT6mHCym4ZuIohNPrDQKmKnvstbH37+Gmn87zwmlQ
HqPhCG31hbpGec2NVWWx+yjIZquQVG1C0hFbqSlDSfEJZudYFll48kE32wHQSAbl
wdRzrc3NDMcGyDVcgDk5HLodP+PzNCU1RzbDPdKxZUYxNfnSz6GZhK0OGcXs+pPw
MSAo5ryFENy96q/lm8Pp5PrOk/q3bk6n9PPpGf4pKyF/qL7ESamT3LVQhI4etzAH
/3baFDB2YL5lpUGIbQAXNRiNE6bAm79GAod/hxRzvI02k3E6F3dbKlG0I8Gt2QpS
e75fTQIBzILSSN/XGi6eNLntveb3rGBoCA0omAhb6mfoMP0zH4E7TYjttXqFBj/5
Bh3YMY8PVcfNO7u3GzlUrXVhxHhByTviJjn2nACvb/DoSme/fCPSCgQM3D/m2GlX
8PrOvyX/VLVIyS/F0jhBvaOkqcW2YKrWiiEwyP/8TLOW2lefpZ8s4EPSpjFm7iA+
BHdqXLEELSgHEzoQG8U5vnYvZin7aHmtTk1xSRe/ilgmPplH9meBIcviKIC34xGe
Ym0/rUh2NrNbXCNJymtaMeplA6jI9NjhruWoPC0a3//wVoT+KHjA+wFTjcVtoH3P
zCeuGSrDZuz/8hMyYvjO+SE5tlQSNNq1eHIMPm7zwbravWJ86GqXDBFWgJc5GirC
8+2GHWryHoYs6eRcMiUZgreu1tk1l1JvqVFBVgb5n7yAdsSNVUwkHpMBwMOoGK4V
6ssrX0KS30Ngi21O46TJolbMDkVsjtLyU/wExmmdLz9Yiy/WEHxlJOsqRYne8059
Npwh7h+DFEF6SydZXXlPlFc2aZJADFqKo1vecTSozwwJ1DnS+4k0pLvfi0YW+qXS
g68TtPsxErCOoGNrsYHSrElwqcld9wxP16cQ4zYHj8L7RAsVTuNZc0E+EHo6pQ2t
FqcK1E3XgU/sAldF3qzzTSuS51vQyt2EZq9UDEa6t+H703XVFcmuwOfOXDouQ+mC
qjzCJrulLPTiMTXf5YxuCooEEVHJO/f9eaWu2qCTF5Ne7NrV2pGkcNLv7kR+rU0X
tpknaIEazCLbf8XXU8LVP/VCYwjo1Mjwf05YiPa72iNblzTac6jWihAGUr2sxQDt
HpX/dlrX2Xkp7Ad7Ld0ov6XHbvMfHLtfRkmYuqNs1LnhZWQ7a1MUBDyUBnKgcQbe
ZJdhdX3W5L7U96muH7QgU3ZH4Yhc4F17/7uk1+W0eas+h8zmU6IYO5xhypllrlUY
uM53qS3zS3KOzzrZw5wfwZ/XtB6U0TC+COYfjuiAf4UvnI5XK8TFeZyAGtGSdNGI
ptE6tyRwaIIRhLqiHACJPJtmABGFV2B7M3dTQaHJ1il1B1ah7RcNor9Kmnn3mL6j
bTSxYZxnlZfibXAt09LfJ0KgHBUjgxaMcmXXhtIynvGjh7DGrowDVwcODB3f3zJK
kRNhqP2GRBpECN3FHvFwewVb4dHQDrQS8btI4Lou7447obRVm3R2M6XVrHHZWbzC
YB6PBfvASV4idQU7Z5IArQwldquBwPsFb+zatq48rq83ReJNdBtaTDK7HxgxFekA
UxzeCQ55QpRsb7jl1xVVvfalx36wXPXscmlzXm4N5s0+v4b710pH9aSkA7few/nR
DouLca/qzlOlvaXfmPTCf5YtDWcSHP4jKUoJxftXWoL7rk4wTM5pwoQKWlcHn4Xg
OhmTShOcUdanASUm9TdmiCu/a5HK8GHxGzIzuIzIlNtqF6/2tHpAQB9mrGKOdp+H
fA04pSF7SL+ncRdxLsequmaBTvOWTwtYcZaR4Tjm3AJBy3B2OShMScT0ITkoK+iJ
xRg9Y5G14mo+jkLvNOSGj5r6b4Fmgta0mI1aIxYP/4mhQF8WqyhVlK3C9gLCxgaY
Uy5Y8obSBrI65joR9go9qcR5cksgzVB8h7cH7/JNlJFwx/4QyJmDH63BxAsmeGAF
sumnI9RpWCSHuJtjkQWMzynpborcpKAtrOh05mJsZIZUSTKaQBCDIknLaqcIipUM
+3eEfN/wz8CnR87YFeNFXpa1cLFN5/o9wYc3Kk+kkdaHAzc8mEa8RQJFsZfucT5S
GMwt2tZcrsNVQd74wLvFTozhv8F7ut53Icl/58npGo6wLNm9xuwekAigJEKi6VSe
kVA0b7dvXC2cHTOEU6a06+0pmCk1ZSAVMzYMUfmjIkqKUvUVjloQIAEtH29hS1HR
W8k9bJchObZ+a4WRY9b5POF3C8hD+6jMqjohEzRKd99Mh3WxESziIxH45YAVWBg2
UIbINnYFg4XLRu8bKgYy3v7y2Zec8onR/Y9TZ8+O6NC1fANskpRqA5rfMOLDL6h1
e1qynmGo+zi5A7zP1FmDsDtaPCn+JuHzHPoBpYe4ub5YOlgzIvh4BJ7W85nlaYgq
/S2jkpfuZSIm/to9jK8etwK7G6De020e+sOBUGvpLM03mkGb0WYusHLpJqWxqyS6
sIxxa059sb53kJXT2Icka6Koshz3IixX8V1Us6JWE9ZgbVwoyhG151o0H9JDhaK/
dz3nSDEnzRNMSLckfCtDEi/oSFiapFesra3/fRGAkLKRec9lHhUCR+dY5R7fv6i7
462VQqP/lEF1AWfbwr+tuDF3xVJnXuajQagxrUiGp5rBp0vP3jG7dYsJhYvNn12f
twiNL2rBJXyiOv2aU667t+nQ6Ux0l1tZIci81tFiV4b0P75nIBAy1e5LEeP/pzqD
KMkiJsvpyK+47hqVrvABemX0/yk+SyoAKSzUHshGfigkEK0Hj/ICjdELLurXK3gu
ApbrKF8ZLwM+Irs5+wdFvFplRrKhTd7hbyf/9mibdPPgH1JE2MVFbg09rJ9mCSpx
RfrzA2StxTcs+yFM37aW55aNbMXFbPNYNYppLt/IzZSJubm9OMk/rQXVRLD5tv3B
E12o3wzIT7EwC7DvzKEgDeOftnIct2xuQSAOR9OXBeOgUyx/rIVBPWzBDZQcG+YX
o3CW+706mG++/Y7DyWcdU2VW75po9zg53KF3cbXpDwmMRuIQi2DshzLOBuYmB3z9
zRxKkjQwKxrbDHuT5YaCfdAiKM5fAEeEjm8KNp9OZXmSRN5BdSfrBL1ElDBLk/j+
RCH4BWBvyhjbxPMBd7e8m4nNSqgRotBiZuZ0PM9iyvcv9isbs3FX/Sp1qOZRMp2b
F8hHtPSlWLQnkKXTO1AZPz/M10O8rTca6vDyPXzaJ7dapqAdVfnQQ10JCRHv1LRB
zYpnBOSCPNbImsmoVwJgw8k7Jetmv6Bk74H5Zao3AMXuHiAhG2HEqhxu5a3TGyMK
JCcj3XJlcEcuUTnPjtqmftGO0+jJubhmWw0gq7R7yFr5RPHzibjjTVKHT4hoMDjO
b6TuTMXq4MZI1g5RIXGgbPig3Da87tUaGK1NetkPRItmD/KOXHMslEcWnDGlwARd
jjlt5YRYDq5vxypQNDLVBCMhz1fzTDAFBHDl0mIvknXfGB3BOWOZ9XP6QPQJo/PQ
kjiw9w3zLrVgaYfAE+sh8pOWE0it7km49ks6mCMwyaVPZpFp4GRSi3L43CaAmv8X
WXbCLtrQKJPE48hcv2UoyduntQErPJwu3jIL1TxnyOX6fzkCeR1/HSgz4xCb4Trn
AHbXNAET2GwFyXGlChtER6Kfu+pe0nu+tvdkQjfuJ5yNEapkG3XGmGCtuz2OJ4nv
m2Hg82TnJNaqobHkDxcKnl3BoEcs1aY8/BUbg7cTY5oicsBGBhSC/3UyN4kRY+Gy
FDoRK6xKfgCVh2PAwJzONdcF6pLjmxQTn7XxfelHpSx01Hae2TvL+mGFa8zX7IlO
oQvNipgjKppBaw5Bh7PWUSvH1nWTafV122QbLEoKxjPCn4s4WyccpUb1ipQKmV+Z
FosYP7LTxaUPiqTyFKtMVpglijC3x/9JqrMnDOv3lBOJ5GDW6j1AkwP0r/qwOjU9
kcg+37PRlu2Rcs2izU4rymUlmcl3NmA2XZ0nj9JUCA419xLXzxovZpM30t8XWeCl
FLjMmiu/AK4JxtoNRpHX/+Ghkl6h6S6haH31cfvitykFDtjutNA5GDJLtR11S7Jn
C1YqZy/F630hfXG4ula63KYq4ZJhudmTUKqlfbGL06mD6Zzy+o1KJ14YG2h0KN6y
8QZcHfQmOtsv/jI0SjkD1we76UKSenLOWDMrunUsBDJnzWDaY/l2647NAufZBsZG
Sfc4Ho7qgpmgzZYF6dYUh9kaFMMpK5T0J0+tFpVUTUWbQxt7H4pvKfWrtFv/wEb1
E7h291ZKuBXVL5E9cW4E/GKToEAXlCfa5FhHoFnST5lOuR8+FwYoHcgPnJkNnUQB
gZvJnjuZRv2/TjVQ2u46DUj8FBruOn0zpYehJ+fWlS8aXeuMZdrIa1Ml0MZx+/cY
/UymgDEmNa9OzPreA/fLVidRL7ZU4RzDsU1uejRiEX/1kBp8NdO0/rRtwx9y2wfv
53QdESpc4TpNvKC5m6PELv202KiVGGD1DklAGjj08hMMxpfkAyrF+bvEYIMRfxQl
elh4ZOstFPymOlmtqlzqWkCLzcpEESE4i1EGYKVWpoBltP+sJNjfKB6vxVdMqEh3
udeMbsUoFyrTKq5o++dQcdUTAbnLq+VR+fpJPp/eN4cfbulJKdJ3L1w3eBpyb3CC
OpXkWpmQNXngZ7rgctThA1rMhnXep7BUl/rXUaMvddi5zn7f384bv4NiakvNr8Jr
zsuvYpg+sT9Ytp27HkkXmnIiTDtvXX1KxG7ra5JIHkuW+9VZxkWKTkGpZrjQIY/f
j7np/2oezFkwpsh6SO/dQ73aZ04BXTkFgvwX4atoM4iRbtKAsLFaKQSdUizjrFtV
j3ZUsUIxaX5IYaRh8Svhi6Q7BBS26gubtsTOmA9QLE6Ivhf68x6OtoKyjrDtpPDZ
TKZpWXJLEaskEOjymaiMr2E5Blkwso2Gy4vn765KYrWOdN3btQCi6wvHdklSEwBJ
hgKa7GIak/5j22sYXFylkp9R5B8ciSYDEt0dwnDMrGAKbqueWCzZsnpvFJX2U+MV
veGmc6+XgWUMWLwBID2hBqEhHoU8sslC+pQawKjrGtrFRo4oU768KfJT0BECzsl4
5t5oXXctmeWlsb//KDIjryPU1RUJ+LNN5xtQO/g+ietJYmA4tY0QY0mRpCKuFHJK
0l8JKQgd/DhZx9ZoMIarhfC6lRcdAkj5aKvCT8yI2DJgnVwG05pfKrq9uyCfNfTV
cZJmJpaijq9TFN5YAoJivCGdNI5XDq9oxJoXRO0C1nfJgO1S9YY46ZHhIJZnitJj
mZstl2EhmNhBsHOcv51bWsuWBCpzSZGABk7vvsGouvIfZnibGN8UafHxNQKIqjHC
e7H/Aw5Mht2ztJYdxPM+AqbnacLyUhxwJULi/FEWpsjTX4zRg+9By4raRGVLRMVK
7zXgdbvvEAldL5GDFww5C5NBA0ejMho/gWtWv2UQBtuYJGqK4jH/fEIZNL0bjsGp
gp9IaLQjAs8SSFk36xMoSevok1vUCVZPdbtxCHcRYUBYhgA5V4jveu5eA/uYsSJB
hMsM7/tXUNqPxCrLzIEbCHjO3ax2gxAYPF7UKBfIl/JIpd4o0Qts+XxVxN6gvnW8
cHNYm74CwHf9B4fu6Wnj2w+wx1KI6c8lsrS+OQZQ8vbUHuKW/EUEpDGC1WvVUZ1T
k5FMEFfraQUgUPRiKployMKJiPc6W9fiEALt3DxSCurq2uh6kJYlPVV59F1LU8lO
w+YSjJd3GarvZlsHgnfavU4TLTRxNf7z+B8XVx4OBNEVDbc3X1ZahFeRti6HJcdf
r9+F43ZymPqDxXDdO9+ir1Wkp8rSdYeKz6xBxywpEXszBvvbdG3PgkZfxhPeuwP2
5a1Qh6sOrkSQKkf+hAgDKTfUyvga6L80WB+DOfsbV9bBG6dfKwYClMADxq5Niz3o
CWrBIwizQAkNBbMUdCI1Bgc40Idq4CSbFYu2TGcwHx0sYf1sIoZbSSHgiuLS+wJ2
11PcVgH2JDEzlW0cnMtZP0hzpfVEP1VoJuHfdOQXqR1HvACCeyLcIoVp+0h5zcio
wGpa7ei2AxhZS5lO6MostDDMFWRa0oR61ExUzN6Dt4KO69fkZpN9f7VJyXIX7le4
FevDN/vIFvuAVKolcSrI/DXRI7cXPfxLpBMhmsqxof2PDLAfmaGs1utgEHjhbLlX
5sN+rD7r8TD0Gcqg1OJHny7uUZeHK3eLbFnJ5eFlZWGA4eml93lRXuYZr69N5hW7
qoU2JJYiGTEevUW2UJThX9hWNiv+eSRfIhY6xtTh+rWhOHiCKaa86vMQQeamoSSF
YtRFm1uU3IDaZRy/sw+ViVDcaLTI1qfHuttgPE/7x4a6dNupQenCl56WXMza88cW
bzGSQiwBIS1N1u3IFCrivs8fRBvERy47eIkzMjx9Xs0rjrLWFLwjaK289+PivyzW
NicUSzbty8N5pkKjYajGlL+X/HCpCl0O0cnh3MOsLjQnnLxfmR2HhShJc0mDwOXB
AVex4VNhtUrAscYe0Bo+S7w0S4I+WY0CsCkuiihI4uKru/h6aLrwD3/SFvzTSjaz
lUdEmjm2ShFLKAw4RCW2/6UjC3yN33qKzy7bZ1oYSfFNLmkiKrV+kWoRG+4nuR1W
oQmGAosSleQwrb3/mZH3XyyUEucCJ89mmIs3qnrLfLdbrYjAjMIfHaebu9lCCA30
tavSSAGHLzs4XveqkZrAT4FfNZD7Cn0mH6/0M0k4vcrtgsbPd3qnByBO/n1k0s82
IxWrErnz/qknqd5sJQMoLwonkSk9MxKtFbtXIM0ogpSbyiAwMnEOGVIcgsg8riDJ
4Knr6LBT068sThB+oE3rvjA2lOdH95kPJA5zGwkshr/eqV/KcaBQGpoiVpnREDAY
pfMhv/kplhM4p0wmuBPeb0HE228eh26wM1o7Z1UBtjZLvQA/6QyoEsilh7xLnx1i
6Fj8BgNTVBmrueQCsPFCC+nuHLoPTrGVthilXObPI9+0NgBbMjTMv8tBREHFnm/f
Wf9Jfc9PwoPkNUX4pyQKjB8tGbkfRL1uIG1Ml9VmpURdnzDVKnNoAcM6k4DCb2wJ
OJAXycDTS+Cj6BqxV3e5i0aQHXhQyzuUwS7bnfpm9qlFpa5iuaeVv+ZRHF3udmUH
aap5TWPGoGpXqAaIMeTQ06tA1sqVJx2D8OVObbTKrDx7cswTWXG6ZhgZr0kDP9NX
9etl7Ujiqh2sHacu7G/PquSKUPF27qnr5xqYUzIRPaTMpTv4TqvednCtJ8wdKLTg
qpTxoKfW3N5vCLoHPoCPCSlOn0ZWzzSBuOQuEIizQfaEXDbDznhY+M8VL5mSilBJ
wfPSRr31JfNxRpJKOSLWFB8vcSlE8hi7bKd/38gcIvVAP9oYla9+WIh2FOsdvrNI
EbyG1CDx1dUXZw1aWnume0808dQLzV/cPDXkAUNiOvocot4ELxQIvkLEGeL7baXD
w3y1hTc1vUEbtAjMhnlqoQDFyFhlc+CdJ0ii1Q3PYGvT1Cc//UB+DMn7KMefoFkQ
DULY/jJZQ17cW/T+Nc2Fv927Znea5VDZqpX0t/SuAzljZ1bbF+W1P8MkXgopFyNQ
Lm+X3bHzDkBsJ7rrHmOZ5i2b8oeBkz+SHerKcCgFaCKiZODUFITg5sKxZQDQJzwj
3kkqmbNPRH9qD+kNHWh+MF+pfmgLRux6zJ6xcwnQ1oc6PnWnCMlKamA2UA5ghzed
Ck9cn0pvu7TkKaMINMbWv66HyJOzMFK2pR3NWgmUDz5aU+E7bAZe+bMuFx0oCzup
Q17zaidSPQC8zA16IBbUFz6A5BlUp+2WEgwPRQvFBEEf8dJ98Y7hGhtdAAntqS86
pex7++DZTaPsTXt1Pp5oL7HL5SppRokWaO2QuAoxymKPg3t+fBmvSh4xgrQFO8xS
8wrMIzKSplPmZs62XrlnLKrMim2eCzKKFPMSVmPFxRD424SrRq9X9v4Py8AaekB4
ZRzRQnxuiwN8NFYZI8zoF+lGuZCtIjgJeeaF9OA+H90fbWKZ4v8Cof0ZV9weJgcn
aC5nR0ToO1ugYgpyXI18KAdUP0+CKZtFEfVK2F477qaVtSAFizHBAV4rxowTEKI2
5o2O022zd8SbiNgl8AkRh+IlPlqF2y+XbAQoLkHTyUaWExZ0nyZJTzclbftTWqyZ
7Tp9U8ubNipor8bnRD+KXykb72qL+AfeLJkODfp0h2bEFHOdBao95WLvUwhJYfEE
RFYRBTu+DvDkKiHg77Mma0jhPGqi0NUmz/XdG9NRI/v+CcfeTzg4e6G0h+2GN+Kb
+mcbji4XY/AKKlWyPVV0LETIsEGZGfGbiJAityxpNhKqNdrDZBFZ9YKKQQmc33Tl
y5QvBclPGTJYwUY9cp2VKQXXEJ5vo4eEHHZ1vVv7lEfDlH7z16fM0Wp2B49M8W7z
wowMnaled2vWke93wU+z8Ove8tVUhZtNXFTPreOgPt0Ss2Nau0GzdqySbxble4Tf
FisBNNk74Sg9LEQMJBUI4AMbL/3asFepzg2oODX1rjVkA1eZrAgc1w09ideQ6qkr
QqY0XSz6oSi3v00C13DA6NVN6aYir6dTWppzeyMVQJoOAFBkijZfZAdHIchktODS
y6e3Pv0rDToe1GRSv/+8sHKeeJavqrnqi1KA1U2Vv0ovaa0y8sjTwq3Vax4kF38g
KGzqVxAio08PZkQ6+jbL3oG1ADjBwpOcADbM2b8ZB4hRZlozkBL8OkW0PpPvL0dg
4xe0FrTewb2/GTWZ8Y4gj9zjxmCniBROnTosUxzHBHuMJ2VbgrQYPtbTXXE6Pc63
5p1MRW4AxlISnze5WsYUlcPSJxtR8djD3lZgeAY/CKXvFbNpiGXhFeHBvyESbvoK
uaWV2sWT1bwunc+Dcpg9+pQqw5wCpY+4dQkMceDkuqMqXRxnLXXZBITQuRRpDZAE
jzNn720zIqudfgnrAXNANjepLoO984EmYz8w1aHgPU+j7V2SjYokb58R/DbhxS8q
xmOTvwK6tgOsJo350P3OeVymXM0j1ZAphUkWqUpuPuRXWSTMZG59r7+KiT/UUx5q
89NUgxrhprv6DijAtmSZQrPxahH+7QdXoWH7SPR2oaKIINjHpyJGcLB/AwBU6S78
2Zqi1uU/7c+ziMx0N6CBJ0NBCgBJpXHrrv4zNn2QgjYqTBbL0CNjDn6Sz3u83+k+
Z8tmKPQMyNbAegrdBj2JcEHG707mANJmLi2qeiMfqi2og43eXicHyIKS8UPFaywb
G1yp+KQJngnOPApkdtNCEDTLGpPfw7TFxIkuSbzvkspQSHEzE2UUyRcHdpx8T+EQ
t1ASb6v5RJWhYLqLbd6+xlMJvybE+gmfnsuWRXC3Rlz/hWjVT2lJPpuOJZYrelXY
uolFiE9Ziok4ilBWalhVZVFG9SypbVN6VhD0YG1xZxe5SNZvDuVQXLeypUGn6xPd
HOaGabV/alcFacEZfwKSwoQ/6h2Pl9Wc2yyXuzqWUKCGckK1wE1Jegbx28vj+P7y
41LGUFY9eWrwEucOIGhw/0+o46Z1X4ztaqBhUCWJ5m7n8tVPvSy2ln/n5zjbAcPe
jEZSBgOnrMLK8BfMdebp3QhsCLSYjGhLg1S35iaJ/+qgSoSdv2YeB+ZflZQMWN4z
X8tRTN3e0PR8fA5m/Y+xOjxeVS8IE37hS1a6j2Nbb711dc13u9WxoYIsz84Tu0an
SazIcPD4Yd3kYee/m0M0hcgkOtJw6Gm0MNcudL3TT2iqTFQR5z825oif96gFdEwv
JAsjMABqySZt8KF6oRYiA7Ja6J9zoKr7fpSHkZIbJVvTVMldCiW22RmMvtn9Q//z
c1ziZTdOnrH5hRY/h8tttuX+zrE4TjWhJ+NCtXttMH3XCSWBcb2l5ffu3Urz+cn8
qIe+4KI1YwQ8nQvUjildKiCpr0z0EnSYbYzcHYnwGh70A6Elfz4jCcxi2wdtJGon
ZM4IUTrO7/EZpf9zQQcDSsP4C4VKUjWmWj89GBToFLco6bfqxhEPaIU4jV5iuvlE
GKt4cElabM/XP3/qfPMzOClQk85NUhSXUIgnBQJSnG4a644i/uyGi8G3/BuSp4rg
NfcEHF3seNDrrNgqZvL1OBr6HHpuckOdFZ4azl06GiYIIDABF7IYhUc9aKSA0yP5
5G9T1ZpyOpyyOG8NS+qAwL4Ip6HfGI8X3NOgWQ8a62aIHb100bZ0PRhOFXtmMyb4
qquEPh2GBqAATFWrjWfS0B8QvDWNMyTD2JHbQc98nO3q1Ur/KVSbiUSNHFLbAiRt
sr+z2wdLpRNr/4JWe1LiE1Np0pTGaQoDxEEtsebnLoouyPPUoOjcIKqqQzDpgnrI
vIDol8VUK0mk+ADhFYiLNwihEObBX2KAaZReDBLLDmhuO56EyUyH37eaK1YjXsb7
bkqC32HXLhArwSwrx8y8g4P/d/Dc6+TWKH1AJxJ4DrM3pScrxXk57sb+lHFHuVrs
KHExNipWiO/Wtx3kdWXIbwXbbKtjrr2ALmD+Tt2KkeAdCGwZ3/D8LzLwH1lsuXUy
4nyxyLvZtuUJGRuLxl96wwlIF2hTYWjEvf8xiv1uU2vqEJq7YoDeQECdsIrj2tjT
i7JCTVEPO9Azo0xcGOHuA6umM996XQzFqAEz/IdAKLEvK9+F4zB7zTjWgwKL+rwf
woHhsHcUV25R8mSqtegnxM9MwJvi7C8fz4aTw8KYN5kvzAyICNNHRcnkPx5mEWoQ
ymugrnIlhg/RbEUBkt6zQ8ouFm32l7m2uzlE18Nk/CCXQV72xDoIkPvWDiOJuCGM
/GeqJsTh5khuH3ZX730JZ4mseCjPciXI58DiIL2wD3Sv++XXohLs4tdGwF9d26QV
BYHF7lFNjkHOnsbCXAlrmAZqhJEznMUNMeRDTe/iVQRUjqSG6rF+kTUsBpxskdSB
8pcnLnn8Bn2daPIXaTB+hA2R0VN2Ky5AyQy5RS0GAvuA+DPG5gXXB0BdGuPsQ5S+
gIqywH4ZXfIqkAQWlb5dr01xIOS6I6pPFqlzHw8ufG97pbhDJcA4p98J2bXiZXjE
LfQonXdX0vR+lYwCtW/zObTo0sNqNdog9+Ljba5LA9y/0SssjUVjySzq6IRnJJtW
3++HLPtVQ4gfEmn3IsXRX3wdXBfusJkbiqqubxo6K17OQ1okaAq+uNA4AtdO8o62
x6MO13tTeIY/NtaNNPamD7Lk9WzTZf5Oz/kZd1A/rT5I2b6ztfwLY+Mg9kSs2q7p
6njNl4uOAgeq+sWWYOOXKJOWuUPDGAg3ZdL+oI7e803KQL9Lz7U47dmoqf+IgpnX
S8mXT/Z1M7vea8KPZsxKsX9DfBRHHwDsMidAv9pYfFK4pRJBLRp3dHHDqLCAwihC
3KOIbG9IJ6sB/YZLDlX9tC8rmDM6wAYbv4t+D0anXvHTEpCC0/dITFzSvA99XRVe
kBVh778l/5e2jqRyEVBxKWJEF1ty1nRi/5sfOqKFK9wNoy5Fn8HMorqF3kqLRpzA
aKhzIAZfycJFeefOlCV6RMsQXKBeXYsudHCSXPhshVarOLc0G/YPBTgc0Q1OXYFf
1dM3OdpIg3R0KLA0OvHdaU4n6SDt4PgIStc1RYCd8pcQYkeTgIlSg1BMlNskZIYW
kJPaQ5iIkdzYZ0+L+LyJB/ZD7WUHholADbmTkplTFErlOccxutmPD6fS2ZFFt2da
XcdY0lQHO3ESnpqAgr1uejWBUzlfSkv8FfdayTLlAAOLCmkY0+3Oto/AU7fVs/8z
cBIoqGBDrwmAxjTb81tVW42ixaWLxRL7mH1FbC3EHtx+yNDi2q7Ab+0a166KRWE+
1MIWDQ8ggP6PJc0pzuQI6jGZeQJ+hamBGOsQtcwqJAXtAMxM34YmShjo+1blw0Ts
fvnawy+qdhFrSxboAfrCEJHF2QWqBZle3inlXC/ncpJ8KFk0fUi8JqlsN9HXwvwq
lumyu6aVVsUD5aItgfv1jWxWYoeymRPSNgvbQL/SrWUfZnYlkcNgKkoqRdHrtVJG
ttx+PiSXv6xbw6VUR6TVCKWpxXU3l9lmE0IMUdMu5CNlWTsWw6Hl/IDaaLoYRDcf
rCP7uwueTXHw4aiF95Mo9v+j+MrQcZGShy6oZvHH2K1g0poYHPstAA7aMwg/smwh
PvoGspWju0+9uv6ZkkOnZ7WrXNNj0dscbzBtSdHkE2OgH9HtC57heVe5veJ4CnIf
SDyEwyWmBvLQNZ0Ki3fiHuC1M3c/foi279OHHR5XSV7X5TiOZicuySwAN/RIdF8u
rGRXSHdw9htWNpVGO7vcFCJtm4vMplfMQoM4lGvTKl6P16yVGBtEI4epnNz9hOjr
I9rE+n/wGLm4U12ErhMSZkI/7XLU3qimtxOlcn7j8U4KOOodr7zxiB7TcD0HpI6q
dyXnQeZXQkREEw86x82NRYBRmZ4vmmqALHq/1W+uAib9Wdr2v5hhYHPPLr+y5TsN
QxyRENrhvKN08h1nlcsMWMaQogKYwdjVyE+GUCrP62YABNmgk5ITIaNsf1CH7tGK
QE2jObRR0hsDuwMQkgkJ1bilk5UvZVwI3rqSgMYMCIXt3zQ1pttPzZ5gr5oGENh0
59RcLKHBJlezqwZMv970jtP7fnAZN7X3YERdw5nzQiQKFQ3QWVBmJ/qA3JhkfNgi
S2U2MoNE9TAc93hJ+M/zXXcHg+HfwA0ENxdId7LUGBnMz1sVlbFh0WZ1BoAbRzEi
WNvhKaoXcpFVXmaR0e1i3HLDm7My+Z15LyFUe7Vw3W/6eXHMiVc9E4wqcoAeIPyS
LPmbRFLgNJ/e2KRJqlW2i3H3VWY1ag+p4/+ojV5zJ3uiFzBhJI1DBQ8vXxKTOlRf
fpSGPUP2A7CNoWMjVoQWc5tCn+sbs5K2rfjIxM+Cl3KhvXv6G3MBjLnN/FegKNBo
STdQKO/sRPfeeC4Q5tBtEIEwIVvRVMns5BdocUNqOfTxqjVWW9VG+49sQnGzo/RL
HSOaRassUS8DNuu8QDy3Hd4ZsPAFRuW1u5eKSrnH38zq8yENwR072a1u7fNIyP+l
pbtMrpuxl5u9MSd5cC1X9N+U5s6Rq0aJxodookt4uZqi9rph/IFA287hrpwXp8J4
BRuQGKsKU7vSGEUE+peeobdMcCO82mQRGJGLTRPgUOmskEpRoBhyusu+F8EAUSAp
khaDPSQvLoU8Q/jhCE/4+bzSz8IuoyTArlJQeoMB2otogpBIP1SHIYLrBaWVExgn
RAkJERxjzWe3ToMZRJvyx3fTACnT5VjE2Dcx4DXIP99cturwRrCQDTFMQJpWngKW
3NShkBM+iGNq/XU4egu9NAE4GQrceogxr5zkTz8ZvCgsVSPrOtFv0o05Yd/bCQ3T
k2Axzs3Bkuzu0SDN25m0d8SFlhmh1a60DdKQBW7lGZ43e4nWIzD3fsHDuwCrkXfx
+Am2ZITIbl213uVb4/KeiExtD/Guf7Xje7KjSkUf1q5Bcpy2jO5CVanFYS9mGNKK
/SN82/fQf8QBpessVKKmK+Abw781IjX/kGrxIr69NfNIam7uvzc3pCnmN3BwFhm4
Ha58nmOjTR8dsrRYT6sdzdUPqTR0ik4DtkvhME22sq1igv+DdqD552OELoeVJZe8
ZDSXmfn5Jk20aR0usKWmx3XLqFNL41W8t4eFqjTMIYMp2APxBNr8YrTFWgKoUGCn
RNicc8hGxtAHT4p5v76gO91Jtrsrmm+u515UNLRqI9xW+qyjSr2sIfoED3V4KK+f
upocvZPdGXbFhAutHqlduBnIVwzb/RTblqG+AgyNUhXWjIeK1oOjRhzlxPhAJITH
eNoWoKffCtA8iydO8pJ/kVXQk8VnGmKyvlX6SRX1mmo9Pcf6VdWl1FDNw+0u6K4I
W75+MIH/2sZqs1mjCe2bfpAqlaKVcct5nypf3+aSfRsb/QzQWP1IolvctRFMpYy6
xkpLVPREqAdsWE36rGUB6DQTSwfF9zti8mLq8Hh49Vu8DXJdXk9zZE1ahbGUbvH0
92Piv+3GvBGx32X4HMH1IvxULlCms4AbhJdWgCnCxY1n/8uKOWfH07ZdkAc4i8oM
ucMOirZmlaY1y7e4T0gkUXW7uEuhDSiW+Mfn0SVUr+5nMl4gHsYs29IRi78d10wE
Jx2H/6Uv4PaSpc7bAy20plRJNCtRf0Ezrpr6MYaomjZ8Zpyg/Mk1qi/ToxwZy/Gv
09L5aNDo2V63Mc2tJymmFZG0AhyY/GD/MwutVe7lzOifNEahnVBvyx95S913gTmX
V2g3DPi/ekN1N1/DiS8b+wGrBJ76czJyam+OXhgCXGEQ1p3VN9zXWEbFpLrFNIhe
nA0/BNaF/1vce4d058/FDVGg0BcR+LVprfVHdJQNP6VfMowa1aLjSpBDVHc3XoAW
HZtg/RLjrdYGyUbldjRPhs535/i+DN7F19xHEeS26mqxQ09uO2zqtVVPQVVBQD4f
VXH0YxhdjFodejUC+ZpgGz13+OuawFpMtNH4RDsihA7b1EitxWepNczJy56v/8Q0
1ORpT7QdDrdYg9yksMbnDo7zFiEsZTd2RLirENCkvwGcvYZyd9Q0E0l5YN+VyV9n
ckyvEQ/bK8Ij6Kjflo8rNvslFeWFfzdCKiatuDFu6toO0/nvby+zAs6TpTi4FUOZ
Faw/60gVmRKtfx3UBTezG3rsKB+R4unDLePEW9qqwfIqMAl+mt9iphosEmJRFWxz
lss4kHgkChBS2ACbM7TH5KhommeIg7bPlRoyd/w5EpnjH5chiIcLhoaMkcW5GdLX
ZMSnjyLhu6dMjVYSnbY9EqPWUPNNtKn2QJRvReFDh+ouIqDv+1yGxyDcxlN/NMdR
FHPEpqZBwrlWlMY4jq8W6xnI+x5CZDY5HZG48qXdzgL+r/Ab1msj9/2+68LN9NNE
vKNb/CLnU/oZAbu5SDNWQVPwPP1n1nuu6/bxNl9Y6vkFcwu8p5K5M3kkEZ2zhoOo
kkUZfkSM9JxE6Qv9FeENf76yeYo6LkL+v2hW8sDcrQGdH200Y3JW82Nx+/DjpVdX
TdpUFkIzsULo8WkgaFC9xODw8kvHfdZluZ4f04t0GMsBRUtfkyofcXbSxjsmssG3
vHwf/M/bD6P4h3s9o4DXwloW3ZUOmtReFa0IMmranXB9fCUMSLtaf77KUy3t16zr
ugmh3HsewAH40pfDIN9xCTpCRwYW5iz9p2Mqi1zL+ijQoRCh/7aCHGw/9sHX8pqu
hxA8ymk0okoZXMsu6mPItiXQ9LltSYadQq0jhwLH/Hk863bxf9rh4nL4OZzP3Iam
G297V0zMuZkETHVUWuYx1EyIYgmorTZYBLVMGpE0xd2ADIHATehfl0PET14u6fLO
bLcDtGePcB/j2zwqgE/QwFoEIg1dV4Cdoh9ZNu8B5S5tsgw01I2YlWn2OJF9YBPa
RrFrTmGBD5NYu2SCRkeoMRLJT7lmPJltoWgMoIFsuJ0ONEhw6iBFH9sR3qZvUOU7
nRBxqYaSRIJExiyEvg5w5JA+7yfQ9+OclmXk0KVR5UoTZzmEIkPb8cCGdlpGdG3G
tdFCGypTD5OHh/i+GcDeJG0mxy/iHiq3MFfRVnhXOI3m6nojIiw1QyGt4V+iHl0/
mx2Umn4YfxN+oyTBwipKBtMrkGIRe7rLt6rZhd1U8ue5b+bP/T2J63snvz8SyUno
KzzU1hZ6/j0OgUd2KYVa20zdVk8+A/dLwt9kRE6XrRGR6Vp6TxhyiFoxLkzGk4pG
V/pwqDgTrJ0sSOywhUb5Ea/naoRt0Hj6Py27Uobpvzgz4WV5zv5xoYmsCy5jP++o
IRg2prKI99MUXq9pPiA39BKTJqfV4wWB9TGFduy2NPnev5HfWB4qSPgVsMNSqw34
CAFVw+0IQ4PoHnj1GAPdxVSZQGM+Lx0PURX7DCXYLpeA1T67SHK849Ms/GKWrMvK
NHJ4IwK+dMCPjnuXenAzYPK426nwiFKtl46fH9Rat4JGVGnmdp9UwiK54ieR5U3V
BIPZ4ixfxOTzXq/eukP8cA2GfB2QxqGORmCnQjfgEq2qSI+/4kGgCeS8IdEXHUfw
lYyyvX3NU87wNCjvj4MR3LbvksN1awnKeCqu2MKTv8s9sLIUjbOURnghSEAznMhA
f9yFLX3zZE6sjkoAv97TvYBc3soeRowj6SnzPMKqfl4wfB661/S6LejeipoDkbC6
1Lyt2uRRraLh7Zabeo9UWCP4Es3FHqJ/UY0/2fKIecheBx9PbydBD4JIOctZF04O
LLL4Q9o47Nx9MDJ4+i//igGpJoR+LNPnq3jZCIVK1mxsD7zqofrvl/BWB7Q+PbBP
ibl70VLHUwswYerb2Y0ws2ni+4q9QzzgGa0vzsKYkTjIfq9Wxj7bDeVJz5pnu/J2
PeoNcThl1/LF4ASQ++UxSY+B5WKpKttpqs7xzFHvLtlADO0z6SwsRnbr0VO+HkSa
1d8lKdO36qhDHiNCqHs7lsY8ZTfB/ap74zM2Nf6SEzXhjnuJlbi9/WI5UXnDbn5U
CuVBMxQM93k1LGjcGxlIbkL46rbjNEdQAApUJlWDcE5xrch3CvdD5Ft3VcKKwzVR
EJcElyeMJyMVNhLRoNk202GO7Lp7vxOrSlH53AvoGs8Jw6SHm5BeMfetd/kM/RMX
qCx9rtks0jUhLOGyvpzUbM9HU4BxTSveOFELb2C9zPgI+jGSl+lh9AWPQYL4Yipd
AV9FaOjORg9Xpd2CNKMWkkR20n2yCyuaVeCMvduo8o1DyCYd0b4UVH92Wp4Md7wp
C0eZJ/AcNVxCupbVOli7XKa2V972gv5YEOqcm2wDAjlciuL/Gy4fW2DMUoZQec/D
REoEpDFRrCjyJUSwerREzDlYxjV5+v7WRho9hhvT1URnNGafZnvd35lRUiL1Yame
3WdvilXEdxqLajNNPVngrsGBK+ni55Em5IJk69Qv45I/Jjs2g8BiEX7Nrdy8nPMW
FhTuA42HhtAfFbGJH7SB8NC4y0m+tytSQfJyeMacE2q64uGY4JbiFlcSdBuKNUtt
X4NICg7McImQI5R56jgX1SzUtT7sDc6g37iJRbzBsYpKil0eIMrrFqyleGImwXjz
rdU+X6Du2aqzcxB5sBkonpc+pfFMr7hlLhs/Kp2KDWx7Qooz8FzKO1g8QfaYQTf2
m0kt/6HGoEKOHz+fPDRcXkPJiGVLhb/g8wl2kAruu46tu5zcUvjhVISr6KQ7S36+
1Ii42o3ytKb6x08A21R9G97+/98Jck9ScivIlZlfMbGnjFQ3uXA91y4WB8WapXBS
J1x459XOCX2XQUAs0F1quDGjDeR1MSHNdTZGXRIlSdcVAwpR+8o/O2yjU+7ODXsP
QzzUMiUZNS6Su2z8cxjPZ895YVYfGIzEgV/NEOA0H28Nu9gziM+tg6OqFS6FwAYv
U6TOKQFGRdM3PG7N1rLQV5+EZBmrJefPg3ILphsV88LJ8hrv2ZnOjUMX6DAAvZbS
MSiAx4sXsxhzFuim8qIvZrjbLHht49Cy5rJmmVe5qCazL+TeaQvz59dw3tL1a3Zg
KuFY8RbK6KLmOkbMjZpIerz6WuzZ66FAWUmqDeyBmAcf+AvtiqkGlKyLWkAlx0V1
RdCniRwMxKslT58i0hSF4J/lr0ci7XlUeDua+tSZNdppSFyOJL672MvVOiVzAJi3
X/GfC7lcMFbVCYYkb0/ZTLIaUy1eUBlGWVZkjdn1Uq4DDXRHa37os9lLyyqHqU7b
8whSeTKhQImXVY29XhEnMrzjysWBZOaSed4mF/7/cWsMvvGjEGNOPLQZhDWwzak1
IYjmvYUdU3lyrjwNGQmQefnazAHNGYIl75Tbt6Ci9EZgI41LlNNiJq0+obL4Fpye
1GRRSXES+YplLNl06G11+nkPQ9cLHHhf6uDl67QwVzRIM8LJ96WMcH9ThDPkA3GO
c99pcS9f2VsAyg+KLqCHjRjg6yGdOpWctVy8h3ryh+NgElS13ocARRZ5ZqDjyQhe
NR7mxnBXvRyVDSaqiAn9DbgGzyxO/F30cR806dFxm49RVOCuwnuQQbbbvDHd//I6
w8gmCykoRaRmOpCIaFyuMiB21M86gV1L+BWwbsQtw2nlXX7nu0Y7MDJP9QI0vNyv
er4mPDEN9C8oPoRvj6olqdOxC7nCcWTPCs3FC0Gj3w6WB4Y2MOUAUbgic0J68TDX
0frzirIkDMANuJ977TKes2GyWbfZCKyX52mRYXTomcJZlP3sUTpqSMMywMVxiCJv
HW4Qc8XsQRjGJsmLaOgRs0zB+Y+Lt4C46sEYDTftmcAFgK74T1lH9uhRQyY3yDSQ
sKTbCHbL66ByQ/Y0DIgm7pH5Aw5zgMSYIQv5lNUrQ9WqG/V4pgGih/m0h60mP1gj
S8FqCgWzuNQZgjUJ6D3NgsujfM5IquhsDU28or+aIrtmeTHEtdZQPhp6OyJMjH57
6l+pNJzkbQpKv+3kMZ/UkJ6vUp0A/wWyqoKR2iq5zk8lrOTkGdsK4M2itDvME/va
gKCFls9q1oWsxc5ivrHEk8gbDrPTtCKzhOWScVa6rqAIFO9ScgEywo1kv6IlVUnE
wU2x2yJ+lXZs120/3FHH11J4u8br7bV+xqxXPM2O1oAV6UbbgqLnjrtqxNkzosRD
gJs9gYQQjyCrnU6w+C5cHkNb1quEpHwKrV8X1BJGhT4V45PUbCiTI1Eaz5ApwpE0
Tq9okhw9ioF7k6r7WYgVOPvfBIsR7A35264f5KawKfSfKB1HlT6hpxSOa2KVCX9T
DNgOYOLZP361VmqIyDu5pWsBVHhwcwm4+RfmeEinsRZVA4MM93qSk96bLTjEroYs
on6QSt3g51Ki+oVdz83Po/zEVLFiutqTysvYYkm7NxS6ZQjgHLC/n47HA8LdiPeJ
Qd9l3/Ya3RTGBhAu+i9+5E75A8qmZL3GhF/dNrNu6IYfRVZufyhxxR3+deLunmP8
tXcvPCVY5QlLKyMG0CQb74pXcVACnrp5Pe3hORn0zrrAWMqY3Qgz24L3r0I2e2Lu
2zMVY3DTVNc4St1I1yeuf6p065pj9t4ZbCJuUKOwZm4ENNa0RIuwuGVFwiAJzpa5
1DybwWYWyKQlxS/F9cUdxD8F/peez6lZ1KBw9FRgqN8eVCgVjoR9HTw35NmpD12N
25MnjzshpVkbpU0i5uGf7J9DMjmshi5I6r5wuVPUesuLTNwLJUpFnQodVF4QAvFs
o+nxYTU98zINA4NlNiJs7z8Q16YoqHUgmxdFG9Ji6XmB7DTgMmVtnUM3UW+HUzi6
aqLY550upDuVnmijigXfVmHmO59idrW5eN5ALepsPxTTd8OWa2Hv9kbLNPO05jPz
NRagwSfbzkzp3GSiEs/dildMKCrEAX/WLKbGem9hiFFxIBqWYuj2NaTTJNUlnk1L
4ZpWkjA7MqCg42/8SMwpgpg5HLvYyEhZlWvI5/pQ7bKBDxCoEp5euTonG7EwXTTs
wqPeIZjSrm7t9mvBekR2g9mV4/dLi9K7KuhAOYYuaxfMva1OAgXaskDgD0X1JbVh
WMM//XrubuK1CMboSaa3Mar8zcPt2Oo3WxFASwxbOwTj0aKBjKZTPhcHG/MriMrt
ULqg6hygUjy6FkMGU9onAlHU3K5BQvWXI2Q3qRTxt2Jr750ff8q052KYoyx7DPiH
6ehqpFaSfJUbqSjfLnjD2WwlfCW6Z6JOaDydcKVVMGd8NGcvhzC2pWRm9FN6zOKg
vd6WoIzgVp726AzTVtxQWoAP5fliaxOTJsEBgeICEj0Y7MH0Yto3BoZfUnUl3mWv
rqbzP0g9flgcPsM4k4das4acpRIIorj4TQTvVdyLOKexxMObCVC6ECxhwMuS9510
zVYF2ETpLJqWiSTT86i2+JAOx2+jCBGTcAWg36INgSIPQX+g8L73XB7iMClLkhLu
HaRWGHILrqqmSbOiKyo4NJCQUsMgetfT2PliexOHyFkgwiz2jKSKJ74nvD1c2ns5
dZBlktJiU1tl4ETp0CF+mYyg9J4EA2EMmdlzuW5SpEHaoccAElZzvmiDq2Lazlxg
e/C+9iMxreguaV62n7qc6MD+YvsliFTUkojh4zERBDoKc4ezPS4tEz1dJW8YZWO3
EINg42yf6Rdqy3tu2HbhuFkts6XJI7/BAQsx/vm8CizBAK15X1uFI38/tb8G/54m
SJcoUEWRtv5yqUyTKGmd1aOZ1X6oDMyuVoAnGvVXDtTj18MSwY79MUFu3/kznwQn
3kzXPhjPrMUkCEA/t1doiO7hif8xg8G1bVgIl3iuYLt6lzc42Y9esqWRGhYd3XOw
RangoTXgHXqBRHxyou9dSSCfy5WVnWvwzmogQpekTEFcarKXnqUPohKmi41DD9bK
1T1RDF6u3zfR5n9Qr8OnUF05kQeRuH3nFy5ne6siWzSGSyBvQ8Y/mmOxWgwOTQEP
ufanc0vly4yiKc6goYNLs9uM/CYlvkcccfygnmxwiMixEmKHF/3fm2Rx2rGJDAMm
CRpY15212xv9DIcqEdSD9nCvCf0CbjHiSl65sPfpBBi01L0napELyKzpTEIVzOlk
RfMr3LcZs935674uHb8nTk0mxa7AN9sj5GWDJXhC7+CWO1Tjwgvhi/gpUHKJQAsI
KMbif4TCGaWUTsDw5y0lyEu//NP93t4n+YVeAIS8IpGZg6tRdSpm7RkFoAT7b/Ap
zPsGfk0lmtKyyU8lmBrZYlPJi0EI76xozVpm9dUEJbUIjUp0NB48f2bvSMBeLuW5
lw/1V/tmabPW0KNmTAxfQzZRCrKnaGsMOLeIhINAGa4KGwbjrQURCM1tZ4kuP6e4
Cu/b8Uo1KyiyzN3ZK1w5wIYewVdMxDdleuWlzHCdM1ioE938qA54URm/IxBvCKc0
ea6/NJtN51AkHTPuzTOGu04D+hUQUXYJ7yH0gFvYYAgusO9Ax69qAMuiP8o6Pais
z7GALXaBIrgSeX89OnFY9jBlNBxddM2lf9NV514rBwl4j6nPw5f/eeCLR7fj0/FZ
SDRW+5eOAatLGnXp3Iubc8jnS1AB5OmfI6J6eHHScRT7NSxP283BO+6s9BxM+a+2
1M3GaZrJNHLK3Gn+UMQCfwE3EAehDron7d9lO7/hswCqhB0rRJDkzIUmviXolEkw
tHPJMFkKnhQ/SbuL9wJwtTF/5qlrl5PDT64aqZAygnTp9U2uAl4gLbDOc7KYQYYu
PdgPNZU2WZEUMczgNcpxHewe9716pkfcYQN9/d1/iKnumY6UzjJnouS4NG5v5OZy
p0QcTJ9sUhyAJTARok3mQUs2F8A2fDzNZmAwNk0aAnlQ4128ivGW6PSpyU4fMnj1
4nQeEgC3vrWRf3RIsBPHvf8Ji93v86CQ0indqjAJOQv585i0a5XchPiUa9bY2oNn
b6ujU+SX2g5EeSK1Jh9nJF5kHXGetBWcEnK6C2AFuCftl776GKga11agVUpR656v
3k3ZtFzdDlLq8/W8V92++xlRz5DQxEi72U9DMATacaO0lM5+jN5z43qJaS9JHtaI
OnCrd2C7j5HkMmGId0PBo6zaLMOfgHilgRjz7WHK5fIkON7R42RfeNi2sQgrHf/I
pWPrqvPrSQKcoXQKIqvrCr/Z12lUKicHvCT8V1SCCjHvoQERkj/OlvJgE4jOwXGE
TvMyBVKfIfdikG8YGdLUI3Y9KoecM2x6wc9TDh35vNVYJHTZioPhDo3x7zakROBu
8sW2MKjaA+Szb4mzhSCZJFR5fRy7mUIo+kCBVLVpmHDVrPVJcL1s1xosf3ZIHref
fPr3I0aLm8zg4YEmdzy1WC372Rku8/7Vtb3juqGD3WRXV9T9oawU3izyLR/E9ku6
7APtQWhR/Q7tBS+mog2/epdpn7W6U0ftBGwnFaLc1M/J67bKm7Bt9yAAmWW6nz+9
enhOAjRTtzcrbnU2763g8OtwB9DQ6yUoLib75wuz+bkK328ZipY3+v46ltPeYrGU
pWAdbREZvY83Jq8A3rUp456qnedoBcPiaMeK97ySEKcEuLrNeJaG4aSEi9Z5KRtl
t2wqwEAIvfDNyPUYOCZ6mYp8EGpZqAZObhsiz5wxKJ3T9jGHYM8OdFXpBb/c9n7b
qJnOGFJMTtYzdKDiv7skiX2tIBUDFjWSNu75g/hMZjlfzDc4OQFAtc1mpbCjZjvx
QvY1mIzF8NS48fKvP41Cz3jrAif+HYGzN+l8zE4YYKWTmlLmfY6JMahK8fZEp2nD
WK+rAMwLM+sTfKPqiEJg2I2xipoXmebbSnx3Igemk5RInZAbXgfSAuzb+MLFeJtP
br3AASCCobqygrBGMYHFLehx6aA6+wJBiskVbsNiuKc68CFEUMmMPH5Z6t5L6240
4KxLx8ptWjTjD+tEXUzNvzopIm9i5utlS9Qd96fAmzOzdFOg9DEFDErc5ne4Dph2
3UkyRPLlqlFWuX6wt4aI5aW0h4sJmShBLttfUln0A5yl0cCGl38zsOgKjDbhjTxD
zkni+BK0jSIo97EJwbc2tUxrJfWLA3rUESfd3acf3+Z+87qvPSTSja8iPM2LJtl6
aB4XIn3snyge9hhdGRlaLh+vJ30T+CqBW2KNusWWN6R33vXXdcqCeBM5TSxostSa
Be67K7AySDrdxGkAFrRvsWqtQWHcW7IMwEr46UfK0VW8/6kFfMheYl9ni137GqFi
JPxscFb14PY2SzWtbDwFbIxqtJjHkMWXJ/x8/lo7dTProyrjg20GuZ+CqTcqYwi1
5vxcJVyoF4j3yXV9f5zGHzVS+MUcC9SiBCIW+D6xPsCGbXPM3Dgr+HQIAMffnqZV
F7botqaw+xLOeQ4f1p0/j/nrtp37w0egP7b8Nps2jPy1UyR8XYw3Hl09G82Kzbng
DvtBw5MwOODffVlWI+MY8hW+CzS5TQ5F7film6dMe570McxPBPCc7pfWEpCmX46N
ngd1sGMTottw+0dnz4CnZrnkHOJHx9fdkj5XcN4bD8ots4esgxJ61XXqxVHXEgiT
H8IfGSzoPv4Ft7g1F2iYRJH3C2Ehdsh9yNVI7AP2+yiwLt0bUybM7EgWsHJ+K5KL
VCAGX3uSfZl+U1bvEDOOvJHNUNB3XGW1Kx7TSC4DIBmVW9UlQb23lWqZk/ftUufH
dbXUNOmlH4IvwymsPy9rOog2g9k5x5jcT1GRXVz0i3f4UFS99r4RVFdfRtc1l6OH
4SzE7R11E7wY8DsR8XKcFpiUuAyFGUu7kM6haClwoABNvIjMx+GKnqxNTj1YlYTN
2HPsHzzuN7nf9Dn7lD9qa5E0tWq4LrmzItGJsU2OgLPeIz2iU5M+kvaIkVH5G297
TfiD+ED4kFe6XNQnfCKKd+WmMFH8qPQsFu00NXRJW3EhMOfsimsgY4FRLI+4R5/h
4YeI8KJGnPyhNk7q0DG+3YAXQ8MTHuYVKQePe99lfoX62payCyxRP2vlvRMGzP6q
c9x5fdWIijOYevouAh/bz3fFAu0EfDU61aQ1VLrg+l67tqIkB3O88+VFV93070qH
gXCkqFdWRIUPbQOAO/lS1qWmf6olZpluj/40IoH1aNQjkB0BrQd9TPMEx+Fbewvp
15kg1ZIYTzUNphwZMNyvKLqRpPGq1qSw4wwfb0kjr++6ARdL4IcnuKAcVknVkO2r
mYytkh15yGOfVb7QnoOc+AuK3wWtTnfZSfX0PKT5CTVnw/JmRbPnwL4MHvvbCa/T
4Z6qyS3ypF2cKWQoUuSNmi1UBRRA6zvWirRHbl9h48RsGKEnIgd80sdKvkVdXou6
eRBUMBBXeuxTxIgiY0E88W6hYlvLd3NKqBUKK3xFvpKhGxNsTJWVtO7Zgc/6oyM4
FZxGqXvGwcH5Y7pI92RcjfBqUW/MAE9xC3l/B43cf/t55is9Ql65qB+vBT0kZqPS
jDGw5z65lievNHZ6r6kLJwwIqoAkcq1PLS39TW02n+5+THee9YLq7aKVezMtPhZw
xBz+zJRn8ZTcQ+FiPuhb3iXkSbaxxjk37PZQH5OJnJH+QidHxrNMyEuKA6GT12PQ
GQpKLxy6YfcCjzVUl2UeKzu9IwsSsJbLOzlraiXEHr6MEGLpUPdjh7baLvi/feHR
Ed9L/NCRmqDp4R+fQ+AJtCiP/d+yb43FzbhMvS3hNP4/WhkrH0f2UEo5XVsbCApy
WkXmDOr5cqWLjdwmphYuzBNVU4iAWSmFuPSf/Wbvha13VmQ+AiCgeQwodmbfGLSo
yrAO1ygT6xZ8vHRera2xHZgAbMkYcPsmhUimLgukovHOm+IAfTC2Kp7UNdmXDa3y
6ZVa7C9kyy+2yYR1fnTDWjlO4zIRYq3nKmVTTNDV/VaDBiUvkedsa/wPue9sCv3v
vAbWQQgVegXoOzgEMC8vz9sD4noTirZ81HhPmttpVCP0sXbdkoAlGYvzbLJpdgNQ
oY6wrxOS9RguagVqw+zO3wioSSnTyse1UT3YBQhgrd9KLKZKUnOmNaG6srr0XbYb
S5xDFt3RA5fdhVCiuGqYVz+K3+nH6rbyAG/8MYKXv7M5pCEPcZzjRXcOziHpaGZx
flValET8CrtSiA80skAjXDEsGI+jJW4wM9G0nHrSz3c7x7S/0qfhIImdjwor6QBr
HEATETxvJCH3qM+vYwbyjaKNW3IJp623yFc3du2ahf6xPRHMeaWjHdd4QGeH2g8N
WLnwJZv3fnICINBpwsS1gyqBJ1+34P1O5otWjDdNxSrEwuWR4WU/YkO7mPIxKiLa
E+zL/UWmKerAkqgjF8yPqbHepfS/SVojlGctGKpprqh+z3BJpGxaC/KLZqwM20op
JSHdedvg49M6x618/BXxiIjM8lucTs1vaSafiIf9Ivl9mYl3ti4Au1AQsyTi1TgS
e2UXY28DuP5HKhA8D8c91UPvE4HY4c9IYeNsMwr6ohMgvjAEkjyRHtPXdFCOHOj+
BMuYcjM0cNSOGelJFxKPKk6OzlioxAgrObOyzMDzFom43ORXPZuSDt23nGfvKT+g
SR64iSQbsVyFB+gD9b9b6BjjkZ4L5r2LBq0qbW8oGioFsFercpkGGnmW/fwBzPzk
AWW0dz7OO+d1fCUTSN30IecYKjshAcUM7xhXIhbg7ugTp+KQ70fA2iv7riRnwxhP
QozQcZECUUXoK7Smw3ghMD7+pO8C7HuG4jpdIIAOMjegcwpGKM6Bx8JqSctervjm
xTfIBdSNTCNaJ5h7oqbgqyZ6KDVMiO7ZeHdp5bnt95BJNyM0YHR2pCAaES7vUnos
8m+pY6eJva09eVRD09i41wIeEQD017iT4+4bXCKeovT0RhCfCoUHByiI0ayaWaB6
HuHeIZHo85c2B1uk1mexGW/xJZ0XwSQSiDcihbA70SEvEu0ZQQAFHZ+jyXkaCaO9
Vhd6YeXZtGt1IRuTNtsz0xQvr2N4uBXQ3KWhDMnOExt02OCECU4U/LraN1b5pAfs
cHfsSWVuXGZBAJv54/32oGcoUv/fplivSnuSMB5ZR5itBiQsJOrY2GkxdGscAbX7
VolTVF/6JEyws8QGITTXavROq+dOKR/q2iiH+GxqgfXX4sBa+vR/ufRyShGQC1mW
4Qo9usfVWXxENZbwo+dOUqe5wBSPPd/O/tFmqpP5pG59OZdyOHwQaeiAqUjUa4+4
FLmajr0vB7ZhEE86KtattXfoBpMH6SHNSKIgnVphk+lHbWb3y+gvF2U78KtKePZv
+n//Kupr/ep3r0IoJVTqCvtzktvyosygTi4fFFYZOgZ2uUxBNse1IL0Ut1mbTcMc
0317iPWHdCLYmtQD8m9RlXBZtBI4EV+YZurG433rzsXdyrCzTvzril1EF7lI8V+R
L+rxMR6iiQWRpPcJxLETDwaZbS7vTVZwj7iY4gctZACHvZBYFHoOCYQWktQckNeQ
oD/ihM98QC+hBGu3OgJaJkaPKExt9FOqhkRsIZ7WiqBviOQDBwV6uxtNZsTOb823
UG7XQ3tyy9jCkiI8IOIAGLWspFw4lL03yxsFPfPzMWUb5Gs1gmr4xdA7tz7wZrn8
7tQBwGAsCREkubTcl5z+lXzIjANthyu8YzxR9ScfH8oeVt/NH2M5jqQIKvApsead
cN3LXbaxqaoGNvp/EtnPcZuJL36ZaF9P3E13yHyMcuK/ngye/5JzAuct6WOgyZ7g
LIxt0uu5muYGU6VGfcl8NM/zn/fgF6EH6QTP56zxI2vnaXJiOxHtvMVmDdQCKkx5
Gm0JBgvRz/IxX7r9untYASJOrl7XYM5ve+04ZzV4cyWhg2tcIHMsHtlbeoduT3Kl
84HzKPM1O9t/NSyJxsBsyzEAsI+bsjMcvOdQLvbIhzcIB+DUpdMxFo+b2DtwH1vi
dWLEdgIsSg37wNS9/OyLfEIeaMhEACMyGZT4eF5q87XGG0NOC1UCh8EAyJjgv4xp
Oc8KuFD0KxizKRSFYwg32tplEc/GJIm4UhHPqMBLuQMk10orUhLSq36CiasUl7E4
IwcvCS4f7yCdxz6Q2rsXMNXlJLJTbuNuzcen0mgtzKBHDNaPbrF7XYbgryIPpM4y
onreHa21CjgBtacX8rgYXX5c6wh3sgb1O3ME2am4KOXSr0Is+vj8QowtaMSDZ5Hr
KJbDBuSpH7rACvLcEF1neRj9N9XPVXj/a0Z2YJceHwn7MlwwHtAtcL586Q+e//b2
XNgdGYt2QOar4GE2WK7Vg+dHkQh/xkJDFnE5/DpCDwIIws2YG+/ou8FE/tsS0H/O
RnaImsL9JJj8bkQheWqgGvrSoDNcxr4Nex3BnLM5MtCGfftLdbK9bF59dhi0QVmw
3HD0TL9l5zYyKRFEjsIKvCpfko+W6kx547VSQ4cGE8zX8vTQuSPYmKgIWbVK8Yk6
tO8eOUfxFE54BWV8BJb2xWIN7MBc1l0d3wqsmDEWJn6/zv2faeqKwKAUtnkvJu8/
6nHkd6E+VEKS8OJrPktnu9wjRJu7UbYNxSu5NvaRJ2a/DiC4FoVjwCaNyYgeh6gn
ALojY02dN2tua/72/W1qZXODzZEYGG/RZ0SavuMAExaO/NDOYv9EQAnLXsmj0Ylr
IpvH8Rjr4mt3bZ3aC1EH0yEUX6yyvih6BthZ/XlD5Cvj9fMwM1G1+hHEPdApJxky
uLyAgohFCwFQ1XnSXQsllfRmJMXsfpQFdMpLzoEHzJemvFmcMgomq3gnzhKy1al+
Wy6WDqSJYoDTp0URL/WBM7PhXsoNbJRob734xbK/SchJyXpgX6FeUnUnB3w9UpGK
ibcobzAo1nmPQSSMuEF+J6wbwEr5uL29FhyfD/1K3/H49Ok1hRajcrdtSmgxI5yh
DprThm052OY4Vl53HXpP2U/uYLesM7o9/89Nf/OZo3ZAiWzoQ/PtcIlge5Wz2lW4
bwGo+9v0e+PbfCRlD38psKOaA49l/Imgi8HsWj//MWgQxTq86bmJg7Bs8yC4SFvA
LL3fHJmAxecsN56fOVYSZnP6Ea36DkHhhZ9enXdw+Jr4giOWY6VK/iHEhTtLJyDj
Q2oqZGCkB8JA02d5F8J1/ajrY+5lgeeWjbVmDK3XxGcZKmhgFE6lBl7+TXPXD+m5
j9coGCrL6ajogWoI3+zK/Vsxlo2vxQFUKlquLsit5irlZ9UMaPYnR4LZINwjnQW8
U2OUZfB/COgJnWigTNF9sKqhrJnAYOoEHCg+AAgvYxxIzfOhBolFwn6gC08pT+RA
U26EpHgQtBzyyqBnFT1K00RZN5mO8smoc1FHRk3LP8sZnHbiUL6kJhBpxJj0mjce
IZWOn3j4Ar2bGY6WusmVOj8sfGYZuKU77/N4XhbJ1wPFPP4Bd3MIkiDXUP7HW3s4
v16lvh18QIYtwvgj12zZ9FXjRs9QpAmmXHUtLhSbB4OL+gcm7Jb6339/Viqbb2To
/o/HFGXTiFMR9en+43LAyK36FNO6dnrUt/BErwcapcNEcjM75FSEa7gMZVmX+3JV
pg636LzzgggR/sQvyntgtZVRzh9z/gA4OLXv7/uEzHVgpBZK4rFAt2QVZoNfSZl6
USEbUJjs8Le2SnaLhJE35yiMoYOg2qJTBjpONwC6RTX9qm1nYCKf/JIEvvFYFdxR
qzapsoowiK9cwthNm6U4RgeynGx50q4FfaHPSr80m8LX+mikMSDcDuzpxYO0ZqS1
KYGfJLyGR8bXUEv9wusS5GWX4ZV9XQLH2LUlKJGsaVH+lKCIiPJvv9Rm147UmJnn
U/qaLWXekmFObC3ygXURTNj0b7amhkoNIAM56t9rfF1tV98S2SV7N6fwxfkze0sa
tc1kWA8YXiaaWYkMhmatT6qyHGHGPJhfJhceL9uql6ITVMB5TDcNvqg1kOhG6skw
FS3/IQicDSXyIL95tsuCgIARWfDtZ13kKpB8BSMaw+WidnMFfyF0dZl0tLJiRY4b
++bnKGXV0/6KCYQvvEKI7ZB1lZVb3KM0iPwWdzDyKmiuJY4kfWTIpJ/8wDQjsJzU
Qf7vBlqKCnWjajt+MeW8QeoYdg/WIn8EQz/zd1w/bUGx3GpKRNsV8qtCLihVfuGb
Nf02f/l5a6igQ0e4oXi482Pbzzi5DxD1kV9sJg7qPrBHkFP74/JkLM3K+RgoP5wW
CIRSgzBvQFhyraPit4nXjVwA/ZM1UfqSgzbLQfGaukViXchdLXb8QzopRiW3VL3u
DacqBlZ59DsRWDo35c2AoCBF0UUOi3FkU0WhWjL2uPgtv7DXwsRdzmwMb+Uv3Odb
sFp+JxlQ+8loE9nHOyryOAjP3sCI3dJXyKkema+uFSZ58G1TkzDkw4lTGoFjKM5J
Jt4wdG1R45jpf8deJ1JhILsehzKRIMg1BKTG1ZQILyigCbI/wgWochUkqcSIxkgZ
9dTAnHRY9XsrW3JhzaSHh8IZmK5cta+EglMM1xjtuiZp7wXMf+do4fcqZ7g9JnZA
/TA0huh2YWWDx5dwApKwIaq6V1JZaLbFElcYU+PBQ9iYnRL2GqM8y3FLIWk02y2I
OwdWom9pxQEQrmmEimIjHDJ+PDNfMkIO6X/DZBm1ERTsCqA8CZY2rIf2GJf7TTQw
+nL/wReZTYHutvOKqUyrIzjzkVx3UmB7pPX89gL/j8WlMBjjQRuDaTt0TCIiWFQA
AwcE9QpVIALN4+HFReg3JcK21EKbfCXZQ8nfWWTTDaSgGmUY1weYeDFhom9hKpFD
sMyUAmPpkGj7yII2lVazmakIQr6kV5eGwwiffNZJI5WoY6rXAoxPEQdnyBxM9Jdu
FmqXkOSPCX+VGvG1AByEccWlQPk9n06WQhqvE1bBgH+Hm7yyRAsTAL+hGPO+95SE
T+i8o2dEKLDhL56oBMcsmr2CeIwzyl+iC+xq+luQyMEyEHymAcuairCdnGRzgb2u
i7JB9eDWmgr2o5GWOmfP9zD/8t9KgGi+FroQ+MZpBWO+nGb4YgIBiRlo87ABM/Az
sM7n/HayHwVPEhaf/KI1f4SWctbskdbwNAOOBGVtTMtu2YP1soBUeeWsshpqdwBu
xHdE/FuArsnlSdySAMX/ex/N+opE4nKsexRC2EYVqZ5Q9WoGmEGdeyvwtv4HrDue
kMybwl9EfmdbcnzfhHrE6LGJ43EXi0CqYka72I6SXxZmnG6LuTrv2vMgs/nG5MqD
vN2ubtIylHJe0XuZTqSgW8Yo6sSJBkl6ogU+RnDtRyrBbfU6pQz9GWuSfZjQE1aT
oVL9Vab5enhhRrT41zVIj7NmzJA5DrijNJ8lIBnkExHwCZRZC+kFj+Dpnr5lpxng
a+j110DTbaUVphP7Mi43NPlQNpcfYQcUZNUly0dIQV94M5MlKlE6NFEMlbX7k+64
DvutbbsE/WiaoljUzFBPzwkG5GdARWSw6nnccLViMt9gma4NIM/Ilkolx06UWEn3
RejxTkzlIBXoaKTBF4T35O7IwT0QaiyR18f7joeNfQG3wkY0mf/cMh1ATE42hWmD
yL6/1KUlC4+X7oOHzrCi/NClFAmmlkj0W5n+WFCt2e5QP7BudQCPhNwfrS3dD5Jw
`pragma protect end_protected

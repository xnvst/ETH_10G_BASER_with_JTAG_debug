// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:32 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KEc1nnPQ6x6Mv2wsMjrjGWEVgi3bkeKkfZYK9gyqgM3DGiAOfAXjf0dioqM8FFnX
LBgxfG3umjT/5rYn8OQ3M3lxCxz2IxmgvAjThKYz4sI1Cs3enxN9OZ253QyQuDta
KEF4raLMIWmOWdjkdKEkgaw6ND3xilKPzn7F7+7xZyo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10400)
l8dRJXt6vwxc3kMiodaP5IhY3ZrxAfzuEdVV6Qu+Fu5kvYLJGDjd894E8BNDbgkT
cK1Y/kqW/xW/VsqtnpO5qeYmC3bsXnOTpilV2splkoaeawrWRIYnHTqHCWVhkv10
xhgVgrMk3ySZwKfymHQCf/y/qK1RlShfhSx1wj2cng5xkJrfV7/u6VM+xz23wjMp
AcJtzelt4X05VoGXA6CX/0UwLlJtBhWi4gV+HJM9r87wKI0tn8rvIGVeBdSPecWv
W7kX7zvBjwHHj3iMngZriwmJI44pE40f1C0bQbrWfYjkUrcR4oBiZHdEfmX2TZaa
0Ov/RQrmaj/0YGkRl0ys9qlf8zbkCQr/uf3+MeOH25H8Txw2nLpvwUTcpM9DZtit
/iioNpCIbXDlKX+0C8qIgDVK66Oela8iLFFtcv9ZCVrCzKb0mXzOXYrKj6qOjTtt
6Z33aA3FjUdajn0C95V2XiDxEDwhcRghPzi41LMZjmatO6zDDFDM0IybKUzUSxtE
VS1ZHCpFjPlTfvjAKR7v2DrYFYFhTa/5tet5oEl66ePRd2uICn3+pDVjwGIup3XY
SiN2JXIOBBwpkmXINheKjPDIwE0Up3FYT30DA6C4ZL4O8JqQU8R4IddKGoWhEGDn
8eWkBN8e7M1YYDG0m/rHdBgQXKuxOvrsXtDHguIcy90Gts5lV5pdNGTB9R4+0WXi
gpDmHdkZD/0qJFe63tyR6iVKTu9E+/Sn4C8Rl3f7Bgk37o7DDjNCKMKHw0oOH93r
zkMsNmFco5alxoOaSEWx8Dw7OD9758Y/mknX/UOoomF+ILbPcIa4IKnOt5OPd0Bl
wup3/vNP9nQFnKur2N310EPmkx5hHCNpYuKVG4eTQUoYU3tF5iORV8ziCKVHzzsp
ZXJGRdSeeBcGd7YbqpThcrlAR2hb+2lps98e4m40dZ7xAvycjbvw/yjgdn/49+6H
UsEMxkj9RHZ3+ANIi3ZvS1xoy1LbLH5aYAM3f0/uyZoKiTr0wPvnwijXhmkBMuUe
vaG0qLvO7X4ux7WwOwC16xjqVZlXTSbc1QSWTvJgbsIO0O1FUkP5cBMa9HSnNKdA
f0YaJpmHpyqYoNjnwhPcJWWqHjhI/0KM2g8j4kSOG+gAPz4b7lG/joO4+TGWb86s
f8gbjSf0q1kMSdeu/nhb8U9CuDI6TAnRxmCJkMziPwPgR/fK/GIWvdIPqZ4MG32h
HZfPT6Oy6H14CTPLcP5FLlqBM1of3MrAFZ1g5GtI/iCYbFTIiVpUkFKtRtfTxu1t
YE4mMuS4jonbK8MIXrQftgSdVUGyxvviq/JCM2Lwk3tHB1z4830IhDOnSEAHOVSq
8R+vLqvTz7oKL3/AeEjEUaA0GURO/vV4z7NUWBPc1dT6ETyEVr2w6C0pK69Oa3R/
GPsxo4f+mmTxSi8WEMieZzZWeiWA0HNdWouK1nGEyd4XkFFH9QXfwjPCTHXmQsyP
ZGi94izH8+nH3LY8P6qRoPNFI/3Bp5iXsA9BB648J8sq4JYkVLQNl0k+lVhxkCGq
cvFiZmB1FDS9NEl28cHndswBaX1cuGx6zmH2hQiz3ID2D3JjB7omItunTroXlddk
FsxzsKFPT63vD324gayNe+NT1WM9qYZ4peVAaoHjGsBzKQ/rTHuirUH1DQFumYie
BkD9JHVUj5RMQpFhxJEFQJqn/ThIjJQDqOz2fuVrhlA2y/E4uW/Ux5nR3f4tAcB3
552s2Afw4UUtTSIEgMwfZ0Gb6zm13PO6I7wi/NrAAHbmfjfCOZ3k42PBaT1Ns3qz
uUCpyJ+sKObH0D39uBFaBzYsSN2hyIGSVByvuZO98pz2gU9PyAekdleooFF8AO9O
vvKeSZ6XxLSUCAGvymezbbnHk/pQSG1X+Bcnrr4KwkmK86VQQptAK2SHCcZUv2Br
miZkH+d8l/LF+fqcGRLnRXPIfpnCGmoo2vUG5yPTpzjI/aksyg2+6nFgJi1Q2tvC
egbzBIO7rSMI4tyToaFCmije+Dxp+ERnhmqic7KfAqxGR32IGr+W2fzEFm1RSN0C
8kQ7zjC502yTAnDq13zeX/lyX4TsMBGT/D7kZfM3fxCo1vxpKY8Az3T5qS8TkNC/
0jhod1u/eFiDkwGD257wN7p/8AA8J9lYEzwrkHgCn3kwreCX6698KxNMEr8V91w5
EFJ0MAc2RloSrf+50IVobzfRWtsXAAa5MTOIqmaW74v8aPO2o4ZAj5RrX9eryeUA
0HE0hRAXK7XJeFCWYbr2ZRo+SBTl5pCS8x2djIbk2M8VdIhYxroqj52PPDpURjNO
V49G/vIl1RiHJeH9brgZj9Bhy0fUkTAazwd80o318UdLvETfRm23YXwJfh1xd9vc
43cF0d9DLHJJRnFWShWTpsLEL7v4yL/6Ww6wlyUKDoYlGPUqatW/C6HZWfzcIqAj
UbZXk/5hd6wfNTUSJQd5SrR3Vnray+mK11ApaXfGCrteKsACphK5NZpXf69QSghW
pkTkti6lXF3jAKv9oqNDZ/n481fhQV7aABhLikM/mcxpQFXKoTiAC+JO0DTUrwP2
ZRv7jLuvKpqnSNUiHNYfvZ+zLzdoUGbBziIklCKMd1XdOPL5JGCSgblnnxiVqr7y
plNjWjxRkwI82xrAx/uWAbSKZSfZIMZr2kKcQWts4tdEYm7D6h0UGyHA4w2rDH2F
aSrA0F2vDndHC4JrAMkVCv6qn39MkxahKXTqimoa40e/V4sWAKG9tdvg16s9hcdR
D+YC/p9MQW7+r1SM6cGQnzTbePIzlP1OqTGErTmCLgyT8AP3Pg1K+Xp05HyFdama
UdrmM0P02xvQWWORWz1k1y5SqRsNs+x5RKH6JLx/cu9kgyA4UEQxryehHjEiWcQu
cPMOIOIZCSEE3+jCwZUUH42fg93vGzr3PnyoupLroFXIeBfty4Uhd19vHr3hYGb5
K2P8bM2wi6wY0E4e/ZIoNfcCJYcMNAnxMNIVNI5l4nAW1F+ZrVdadCOUZV2wHpwu
PwIpP6wsQzTjHT0vQEUDd1zZt+3mylGGOmLDCViXlJkV+WJasCvTcSs6Gve0CejA
Fec5Lq8K6GJP7G1Cn02QzEFUYQW4ujYms2eoDyMky6Eu9W64CpFACgaQE1A4kY7C
5qRD5ssuPcoBybtIDXPiNg7VAYCyA/gy/AF3msmgDBNtwSKNcbBHJjO8XpNbMprD
dlbt1Oj83S9R5eFx5tbTAwFCdxKFr0igDZRRbHdXtHRFVBF8a2EP/A5oAy8T01op
kYxLMGXVMkNrvx7iKKg/0TrlrOnp+P9zxeZ+trBSeUNWyRp0krcn4B5ItyTsqDXK
4mbNedWwflLKhFAQcLs9pCY6oxHiF+EqyJwAbsOrlHP/J2gSloMGhX28bsHJSW4t
KysIE6qs34WwHgo0Fd4t17fIDQ9IH/Rbzlxr92Vtx/XHXDsGvbdMezuMxgCShM/T
IDzjjf96z1lL+GzPDe6tGmj8RjG9KD5i8ZgxvwGP56D48jSsgZ7bVK6AQTDdBoQY
xE7MKXlmtuIjJoi7DN2ZU3+s28bGkRbJfKumril6C7pFFCZJBAkKwVHZvm3wNgic
jfjnHBMAGlI28agZvKTjBIOGoaUr1MWQmaxO6xyxux30E46lpgJbMtCmJxFfQvml
SepuBNXGvfCJRLpzFQAd6WgAj9YadevPf+N4Jf2YpTwZWjb7tAaaKBvKvOKwsVSj
lYBMGYI4sZw0eaVmEvPLNVP8bf1AXSLUCyqq8p/UskMAXrW8BIuW7n4Od3wyWN8p
goQHqiid5DHnLrH5Yzywxjv744Ia9fKwp0C9hB5JHr0qSpwrBdva6TgDhwpOd0C5
yXKg3S94mlFnqHL6kigOkJmhcJ6fgXmtWyDLBBTNZQ3jKu1KSNJHOlkDXl8N3SkS
fWQthtCbo6zsHRaFECja2ZuU/FITgEFtfoMHpa1X7usyawoaNfiTfP3c7SmmXiNc
Y8nkSK/tzMQE2Ddz4zUhDPKbnnQP+xyqXc520vkm53pEtRcH9rmQ3nIQublkSbHE
Vk+IkprxX7mYVa6SzsmaSDcWio6wtjLAy5NsiTk/aKexQJPtTD7mm8jsfTukqY4X
KZVjqYagx+8HYKv7EKa3hYp5j/MWRJqTIcEseJNF2zBL3L+sP0+l30Sh1+LRS/0/
/5asE6MNGrIOikoIib5lP7W7Rt1IA29nxlPHKbPGXGW96JS4ZjObqU0+hbqplL3b
j/PzLWwsxqPgbqyodmpSoe5EbIQs4IKVwPax/O+ONzDpMINUjnV32RTEhxFFQTar
zu/edrULXl/JYC/VgSnc6UOfmSq0OzzQDLhAA2Mlj0MMGAc+AwRiJ8JryZB1yvTA
b0ciLzUtfiEgCOo+HjeLlxByGMVA3oLDcpjx33jOkKlw/mU9hrlL7czmttmQtjJs
j5SaHHuB42Y0DDSBKgM+8fmtysgSWuvK9FwCklxAou5pzf7gjZVedSlUbt44eyBT
7mDXc6RLkyjC1g8LODYT/eLA/iwg1XkFgTJtEoDoKV3+EdZg0Oa5uRi38ADPnNw2
Pi0XcAK0RHARbUgAhO1M2uMWH1XafkbzKkHowj9pI5VXGFjmzh3rCDHqfOFEEP9F
s7glOVoTQ64D4t1HPYtrMnA8Cn4uBu29+lNyLXLyvP8ISnpnynpwB+RypOhEiBBq
4cbtVAPi4i53//vbos12fu0y2VoF83LpF2m92cVH/7/sN47ZXsHvcO70KLuMfLeP
b/PPVRYCd0TAXFXuKIOYafXY7gv+tbafKkKb+x15gqoNJYzL9yLtBjI+4unQy9eg
2rGoeeTGsBN1aZLQfMXUr9YQUn6pvL5wyyXq+j95eQxC+TJInKiejiGEHx4l+wS4
FldG7324pXvxufH5MeKDOHE8UsWYB1T+MXRB9/FX6AugbSAGSCT8+9/xH+HIV/vs
p84+rQxhh7w7SSrrH1AOYlm9uAgazzUmovtnz6Gx7ggzHEvDpTZXOUpxwIJslP+/
pvNNzlXTL9taC6Ni2Dns7cwWHnDVVrkHiq5YLoYCclFadMOn6dycNgsDjXKCyWWk
KdpIJsbhlLYYxU3MMScm6PZCxXrK2jDa+6CEz2LRIKHpkdF8205C0rLN4S3HXM9i
grbA6qp1L718NnUc2WZ+9mOO6t9HkcO+O2dwNOW87zldNHNqZrEAp+znHjfd/517
YLu1RvNdPQcpAdEfMw80eOGH5JNvTz3Qcaxpc9EtMcTuJ7ndeZ88afDB29qKod86
T914PsN7jxQ4o0J6SAhsEOxDTkhmy+P4vUmMmZl1nCHMZyjUi030DDUwpC9joVd5
ziAd7g0mUcj8ks5A78KntckX/XOLpCO2K3R2w17W0xqE6euekBiypxLkz5lsVhbl
WKyS9Impw68nvuYmsE2ttbdJj6oSHsUdvi3BWHDE2/rBUmtvncwNEsFSQc6BixXi
JknIyyfHh2lGIdSfZ9TANUUDWBT9mFus3mdZ3+Vnp4AI7X9HIqkfM93AGqFPSnqN
Nta+2SBtmq8EbSKm5d20Pbi9lghhIEluUCj9zPbap/mkLmms2rqguRxgYcVEUijM
1zKi/moupD/4y1MUyKT86DBMkxb5Y/1Gf0C1jiPfmzUyEv6Kl0ur13HK4QzMuLQc
XuIohIiI1Se1kqHDycZAvQy+AF2vVp2bhCJMh8908keHlKcZazoNhJ5i30fdOEsx
BetbM8oRjItAUQ6NvZnADb+Waxe4ZY2mqVs6rDQ45ji/wNf9J89vo7BHDKemow8B
ZrQU3r6UV1ybCT+FKAp7EvxemX0u7kkhhB9ytAI93Dpe+AbCN7jZkX1p6BCbXqol
bNzX6XtbliAW4JJ0VEk4Kb5WYUbTQ3u7OW6YFWiKLIh39qWPJXPqFiiOZlS95Iwe
ApNq0DxW0kcwL7x5/IryMbQoVGaY5bxhqZzuHctQ4FS9nr9G/6Wc5QvXUtsXP/17
hfC9pUdmAz9aRvnrWKdsAjzJcvvUl9tVNJDnLTEHUtu2CgtiTETyuJsVMDpUXkWX
kBNunDP3rqBeT5xtVlKNJ2wbVAyrOYlZsDGCeCdnlpbj60k0Qtgi+lfut8E+SZaV
lBoVS6ULgoTGExcF6egMfl+rUJGjwXxK4GJkJzMh1/Enr+iSZwJDCMAtZOL4hdTh
AWXcfnkGLi74C6ZHDzMcKtYEOzD7n6Of5fhCntkd2Hc7zU6LcJKuoa/gBnaCMnSw
i0JN+p2gDcBw/Gv0cM3lJDuh/0qCE1OwiMO1ehvDoEXexceBikdkJ1DjMXlckzae
GAQtE8VGofxT30oMwFpHdUYR1xUW9PsGEa2VBnQvhizdLvEbNBx/47PkVnV0VddR
9TibFrKT5gSVEODmnvoVPUp4Ns3s3B0UMYRDu1SXGfLhV0YZtkGvNks2+EU0sA7F
Qw1LCYAqhd0v73R2lncl97xZcEz3AKifcNx188SpdmdcEhYPlidy5Jkp6tlEaQek
KGbxL8+jPC78TgP2mrlw7jQqH8rzc59GWH7VtaGSjyyYVkquqGIJpCIeWtxGX7aX
tsimxqNztPj3Q9CQRDB+OSS9I+5Wg2FAHrxUnOXMLnSdaYZwbuPZmW+jgA5CcR3M
5tZpCcpOYH0I/a/are+kWU0q7dWpgo3zprxYzOdQ2nRkuUZh/fv4VvRsQKESBFNI
Z7lqmiE2qD8xp9m89e5xDr3uUkKFuV5qypT1fV7HGQpI5uu3QF4FarrHW3ZxpU+6
F42jAdyFvfzV6i1HrzF8VwPuuAn6i1cxNJ5mhVCcE7MemhsFkxPJMA7Rxt4HiuHB
935HIbK7YOiZacerT+EBAUxez65mx/kFSY2AghZ6Lom+Mh4FKtbquT3xE09Ma99v
XXmpTjCKJtKxtPtrzuNf9Czc5oZ+WQr1MX0FeVMPGLNAarGi0FxqYggzUSLBuBYM
+k1KDeop81fc24U79bdHr3+BAK3j7xOYFj8RrZu5zJbR5U5/E8RMD0V0wxXR1mux
jeUYGnZM2D6KxTQhxds7ipgW7BfTdDH19XDGZyhb1Sdx7340qqmdiuAwcNqrLEwC
tJLQnW3qjBFWrwXZbB9kAcMFE2egPM8++Fe/nQ55l+Xp/4wBDLrikPw6HUT/pSn6
fINM7BveAM3o4F4stLTdrgliWxYLcAKAsTCT/4/0HgsaoX1qnLhKg6Azxplbu65K
FkViDCMRdwb61gMb7ymUAsm9J+S29bWOZ/Qi7Tw1M0h631XxePlrcOE/3aM9q620
IW53w6SJ7Ln5/7vKfvGPydLOZ6jqUQnpF9bpIk6+PTY7SdrShhXmLvzz4kVj+bBH
jPawXpH2SpTGs8FkNbr4FbAX4f4GSWLu8WwSd6sCzVUIS1ivFIoDUUaMG8GWBDDt
J1jaNYhV6zxeQNHqjYVPgG6weZTQgZQMDnyWhoUrXhr3y3Zqr2VeZXix0jSt5HtA
DA0U5SmjdqQ+9np6UWtnrU/F4ZMvxeXz0trHjnl+briC/o54Y+fx5JNuorfMt+GI
VSc3x0rBiy/BF5ZHdJO8LH0JYQ7QARNi9Lwrq84rv+wfEIStFwtCtLhg5YAngMjz
AwWMIryl5/1eM8D0XK7bgIebPAb3p+V0HW6JnfEA1qrJjxkBwmhZ2w6a1yuYHT0i
CdA44NfXGF3OxpNbMWxrQK+BKvB76t7B4ADY8nvARgbE4bzSviEZohuRHqFLB/7x
4fSduzAQ7muis4e2+GgfKNXFWkwcUDTSbIpnlrRge+d6sSopXxDlwux8YcctgnSo
OKBxHCHNgngCLI1DkEbUOqFjhqZfEDHOr2wxZqi15nQcdP1d8LBRNbP0FlL/H8bS
NToBUdX72vX6eFqTa+NIBRFhbmFw6esuzNil8h046AbV7KPfyMwVYEyrzyVXzLhE
o+3ACyp+zTrt5t2PD2oj2YFIXdf+WmjB7smZ3M2ngr/wm+CEhjiLuay86/2S+qmm
Ab1INZdd3FacFKFjHc3+MDy8YHlovxoGw1/N8j/B3I/n8Yr9rx50GV3ug5VisOv2
BD0tbGUkxmRZZePX7cObPeH0ooLftaETuKs892mRSBoYQlhFP+pxJIPqKn+KN74A
eRNfDzgxRuDCY946TTH8vdiWs4cvD3s4QiOlsg4kkdvC5A2wBZwFiqNMWTGjKLhL
ILF3n34yEWOXVTU5couIBYphRn35aayAcBRHLCZ4EMFOdkAQ0B11GHpSIvFeNlWx
cF24oVXPcKNXnrdJUdU5o6JSqEZNM9l7ClnEeI/tK6Q7ge76BwlQCfojChcWi5of
Q7191PJSBd017zd8l0/CFy2zXNDINLsjxzgREETb+LKOqMhxaYhDvR4J887bp9Iw
giPeY6l6YpeFowPfneV8fDJWVIGkRZ/37AQ4THsFZEmxXNuyWKIZVA2oomMaXFfw
hd17b2eGeHGXaWRTrbI0OXAb3gmTULLsMym2Gmzgb6/oE/GVncX4M7mNgBLIiU44
Id3M/N3vPPNi6pgKq77ZAU1f5PA0q5IF1WFFqzux/MSzT4UDRsSXqVQNiy1y9p6b
p7p4vos2hXY9dqH3R2WRWbhEzqCx0vJRuOwYpPCvrkhG/Adcq5Bj5YztwpreY5Sy
6T2XCziNDoyefNYAVC6SRPqs/+gvWwCMynQE/AKKiH5COoGJQb5qUfhn5eJPKCv7
0f09wvBSFIPUEL9Immq2K5sSK1r6V7ttwPCs7aM8Pxt00HSzw2DecVxaE4VebLPq
DuUwguHRpHONgZFR8xR7aa3/WZ1JzlSsVZQgUXWR3j6nMqe7WQcblNO3zPYOkf92
By4b9IzDBI54yXKmr7j41PAP4ASaPPQX+MpDqLCTmInBIEege29TtyX31RNrOkvP
EXqWKfQNmc/mMzcyKEuoHTwyqzuaDWdP/wd4PAIOlD2+JqvmZYT116yN1Gvfr4gN
//vFKCJOSSPPYl1wOzoHBii0SnypQ90f6/Zn1MrOMuNfZG7PXSvpOyY6ayH4DaGu
wyVdoly9UwP5MIVJiVO7jLe0sV/Q+FaRaZWr2YXSjIS+qgAQr/leoDlG3krMS3ru
1BrjKcGkTeqjLDxyBzUHhTrEanN2BWFg6/VH/ejeQTI5qvKEdyUb/YopZOLzbWwg
+ZIb6/IbyZMspE4YutU5QNYwQPjAVKMpLj5MoE8lyNxgGmsPnwdMdYyKUUOnqQYw
w4qSrrdi9IrCiwO5idrtTnTTF9a7VhESzpSgAHrjHFUlcNB5C2JcBE5RtHYrhIEq
VGGkca5QrfUIOBhQ6Gs4H91n/BCc2zNEm4B4g57wuY8DUaBQ44q3ThCg+rFEEIkn
RrzKq6A+51/aflN4nlwYlbj64awH2fIdRkbEW5JVYFQW5mXjUyQ2SyVOVRSqM6jc
AsZUTgS0b/nTY4+MNIuXeDjynchWF5SKzfOiBsdppF+0CutAD2oVEr6N2l1ApMWV
rj3OXxuFHUHE9lyydF4M2SGoDPngHO+iscgoFZT0eToujUyR+ODyw1F8UQCPq30C
aIBsFvNtGvgyDQfDo8jmrsDXkyJLmhXzXUWUxwA/VI1Gv2q3NhZOfAKKjRUxWA3q
ZkPlEML71b8SBj6+skCs1g9AGBtowgcUufa+94r5T+E9PNeBStNaKE17+PpLVTNC
Bu++zgVGEpbJRImG/bCL6p79i7XjWJSaB93qoDDM+cftGI+N/ZSlYsGNmTzJxte8
xJtnDJQjEh5OQHJ4drs6g2dV/boWUzHtvTrLETOww92bsQXI5dBNI/BW7GAh3/bP
1MZOmHPbAG5mCwzwaDTxp+Y2tXhqiT76qujjKhvwaaD+tCsDZ/jMeVid6eCkM55U
r04zP0ZoMLfMZ3ns9JptvxFnBvLh1CTU/JkKkRJIxeVD8F9fGC1uafpBovusoQSK
T54++paYBsNQAhjG3LkJ9d9ex8U3dkhk75Kw+02D2qnv9cHebynnYOpKpA6HZl2+
uGTo7xiHJc1IUdFKEdjG2Td56mq7q1OV+TZeRfA6lPvxXQFWuDwfmM5uct0kL506
18z+zXVS/vrLhMCb0drSe/EjQMkZUm78NUdrz4lNLGpF5jv5T/GRt4q/wq3obZty
2olBT9UhihH1Fmn2eko9s6zAtK+CgzOGdTCakTdRzAujaFey8UlPVRcJ4q2jkFgm
/i6AikMSFEU+Oeiiwqva2KRC82hGANftVt06RO4P4QL29FYmyBa9c+Y/nyfmEG1S
zEyUnHnqzRfj2QESnMFfe+cEZtjLR+C4L2N3uTHBABIMMz4nRjYMgy011g1FIkfA
y7oIM9CR2VagQQJcwvnbFGReeKDwxu/CtMAc61CsvPnfxrjrmK7WVdw6EyvbDb/I
xNKQC0s4vYINkR5+OwGQJRoh0Vjau75QkjOmhMCJs6vDCzUtvFQJhqYMP6OKSUfd
yot+XiLTRULLDo/q81ozYa2d6OLByZWbG3zboXf4y8/leeo9gexxWQkOYp2gZ4D3
f6BjxF7ahcaXJ4xQIjxEQY6j+Crd4JPHmLW4dFM6GvoGzLK/pk8O/8MmlFXHDAGs
UVTCoXbTXUjEWjC6sD027M7DqZ5ujJ3NsQHEpzvRXTDN9uUM1eEanSLXKzRpPLeP
MhB4V6qL8zDIVeWlnCLPnCFU1OkPcIlBt+5sZrzU29326edA0i6v/gEdzO3joJwt
N687syGgT1xzbNUDUU0OtJwcRqLKvUvwOoPN26RJLGeADt/lnTZJKJtLX5SdVM1b
Kw45YKnM5DYHdQFlDSborm+kiAVTlaUM+D+C2k2k24/eCEDNoOnjJC2GXdsoES/R
Fco3N3lDITeAr3edPZIhyafjX+PORaRRAmJ74LaupP7NqjnVnpQlWHWDaWHrCrQq
cbpVc+VK5SkBqUJm09g/p8EmOZ2rypD1+TxmtZi4Vq6kMnPT3FgsRQI38U87VCVJ
gBCy4U0meZZCjWn+k3bsR+9slnq1q6OhbUEDI625lfWvk1ivBsgtU/lxuHuH4Csz
2cPlUHw0i7GvsXyz7bRjHIy/LLiQdP6X2tIKgQkPfCUarYGt2/FvwqQcyNaazVxB
WzSnAGttlyTkfeGvYQSPCB4Miz6/z9Hif8GRD1hfgEW10eKRfUgpqaRMU4qeYbA5
a0tqMtQJNqDpziqZYsO9wJ7M0HYQdT2OSciH2D/pggX8a2ydyn0LSqiWkRFc3VTs
NQ1aYwVqDIFGGWoGWTDke0qK4etcckcJhePWyQVA918P8P2VI7ssG9q/Xly5zqY0
tVH4FSGbHvva1AaRfjqx6OTJCfuDMBgwr/Ey+DBL1dcIenBKfyaZVphs6KArLcmU
ojp3twDsrqy91gIBjOINDm9XPl5ITRMCygb5l9VZ82oYcBVwDoYUjYbKa/f8va6X
fzDIeyP4SDmGZHFEit2va0Dq7CTQ8f6Wnsw56JnEOt0VtsjsqYHlq9RWuV1CvWYi
dH0QsNwOSVripntVzCEUxXb2WoiTo2lLMb/PfRwjUed92cz57ORzlQ0jlEnNAGoH
6+1Qqn3WB5TkqoPMj372l0A2pRZwyx1AnYTgyz1sfhSMY5FAFnr5i9QE7jDzXTgi
o9qwqNxlig+4zp7qKVJ6xhbwOsZOBlYbpJkA7XPGswMVsqVECxtD9QYcg9kASjae
Bvmo974GSxfmOqNB0gKMwj6KQCBZmt1LCMvH0GfC0b4hN9XUQNRo2Jk04JfmeeoR
f/XL4e+SG/IZyeRLlRSmo0maNivtMuvTnzqeT6WuyARGB2mBMQ4NOWoL4Okw42MJ
JmtWVWhdQtbXTGiRBtONcEbvWfdhC9Ss4B1Ia3qnhaQdIU3HZwaIHNex+PHfEKIe
6FTYKX7JpfCyw9nLq/PPuSH6MG+91ARsXO6cvIl1SqxxGE7dB8wf/e3fBKXXlF+C
R4U6PfdRFhIJTiNmtUizK8fKysYaaM4OavNKGK6Y6Hs+BHMGIHMoIOiQFR8d96hj
hQn7DN2ZKOGC4NxKchpc+RF8evsdglHDp5Z0qAKQpFlmM/b33qnSRBYdwmi1qjYS
eu7KXH6EJdzcNMBEY4g3WA63+ksMKS0D0klWORIaJxZt7jeXbu3oGOkg8vPfmVXC
gDgJcBxzYRQRZj5khJqWBvfNhS4Ic5DjE7adsOabJoPPv44+CtzSrKEWE+N9qLdG
d+I45LA2PoSXIkAmslganvRt1jhKektdtcooOx2qUZSO/xKrW6l473gxv3yBOvuK
s/7Cdym0bqeV490sOEaISDCB0sxRj0kPFeeuWoydxIE8n6YvMa8Jtz5yE7TRAatb
iAMm64Recr6wbHRSgmNlb+jJrhznc51HB77n+w1AIxEJg/R0J7t6A0kCezQqXvsw
wjfT7fFeNjMCUjglze9G3mPGNLvZvdQudm0KqJfcxdtpMqpkWmTHRW10tbbL90QZ
SraotCWe/8pPczCcTZllt3jJts61891JWTYbq2GpEpfe0Wmfu/GDdu8uvvqg6YCC
wg3B1+Y4tYlDK+bnkQ2wZ08hMcQF57xbkeuG4yfjQYPLuuSkFNs+PUs86FIWk/3U
IsATUwLWo8Ahj+ToP89CiDc7DfYQF5EA4ZbZtgSyyB5weDtKEXStDjZHTtuB/K/Y
r4tXzTmZfrBMv44DqIKcnvyPTVeqsrQVHQ7Wn/axT6y1PxEE6yfJDJ7J94EKL1sO
+IP+Yq3HYoDWpdUxoggMRCyJtCJ5ZWOGk5vg3IJl464WPBLcXo2vAm2nteejoVgj
7u8wR7SJB8cFV/dBv5ZOC6HboLzeDP3sP8qCFlkztoNIoUYkTPPyv0/EaLZGBT1B
2gyOUrKz4kdiZRnnCW19bP2sST164J4I5boN2vje19rLCAOeN0ov9l641XV47IeS
6dsrSLChXm8RnEKplVd99YI2dEIy3ojRkAYp62K8MO6H8KJNrvdi6a6epfa5Yl47
u+YJ6O9amrAN3bsi7kp5xxFld+Mgt//Nb1PqFE95V7/4mrFmIYfFJ2Ud+m58M1G3
4O7lPXazLWbL2XAUDzTgVcshbrTWevavDmt/aZJ6vkzdrD9wRPxkaE0di1XfgmUc
VirmDNAFPc8+pKC9USL9HeN1GZrFEjI79qpebU67ukNDUAfh/CMRmwwYOu3RWXcX
5UtSSn1eJh03V8rHWLeI6jr8F+rRR9VdC9QPkJauOXjq7bJXYMc11CgWNCdT04+J
IixjiN4rAJfnjOGT2X6tMQLoZ4z/DH9zAnzemetE9QydLjFfMLe93IrqgznoLBey
ZqOH+Xkq/wCq9ibgrKGb1T2rlJgzX8s8bS8rXjqV6Y1vZyjbUS8vE5vFEW+FqXqk
pOG03Sps+vqN0ApXsZduZ/6zBvhDq/joqN+CPfUYibNCT6OPCm6lH2LRSfWcQ6BO
XkxzxN/NpFV2pGroYWhIPYP98BwmqP1q7uLIdKMg2x55W1G6QKJsoq+OjsSXvYi/
+q8K2ogMvpwX0U1xfLM/471uQcMsCV1szjGx7mJRDD30CzqFTTS8Bf4l1tWhEFBG
zsZxuxi29zJQN6CRlnk5gYsyIRx8iI4lLIczvU8RYwuXL29lDSikqAtREJDORiQn
Reo3IugZFOk2NTmGpzPh9P5UBAnMiPkr9cnhueznEGc91OcxxvnSre757m2Ju+3N
jsLsFozFqqsnlT+vdfp8q+ClPG0++9lUBpTW1P2hoi3oWCYFyc9MMqHTPA3wvzUi
othJLePK7c7kaj9YmtRsarJ1tsliTlP8/yzdoGQaXfrVnkTN1nl7h+qyaW/IN3a2
4fvYeRm5l0FT8YuSJYnRzZrGqPKGiOL6jdnH0KCvGH6iPOGLw46P7cSlIFwFB1ED
Zbg02RJE4asqjzYEzoVo9xgB+gTsHTxIyo0or15JFDb2GUNak3MXjl1UKyNxrPz8
rQYkKeEhZxIN+SCDsD8QS2UWz346WKnr7K8zmF9e6Ac=
`pragma protect end_protected

// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Tyn2DcdAhs8owG0rxuCx0rDutYMG8ic8KfhewnKK2FqFmFrS9yPdzhiyvDji2dLbyr0JynZ1zIl0
OicHmrbzKoSXkspJSjhNjJ6V7IFFgoZoxVobuhGpmvT6tbBkjpZPwqb5+GrK+nMn2QYT2rf+Ful7
/iBBZp/wIjwN8d6EBtu/+mBdfKk/HIg6I37gOtd+yRRaZB8nxDRwP2Hle8tC47Y+ZLR2L07qwJZ3
esnN36KxDfwjd7OBq7eZ86uSTP6yw0MeLwelWMFcSBR7fDjFxBKL38RzyhLU5NDWtOIpC1Y+3+lT
bwy7P0bPVHTo/nuwjMySuSySxrzaTPC1RFDLEw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6mdoA2eSFNl86wDzXgMvAJUU8qdZFQLzGJw5133HQ1WTJjgcT23SpOVE2GcryVGxZwT9lgjptkFd
fDuZ47a92m2xb4epfqw5pve26fYmS2yQsrQqAK5VvWL4zHeX8VfCWRgXKc7k8QxXJUfEFW81NuFm
gM0DBu5ZlaseLeCQNQQeRv3km19jg0KE1BxBGBjfN5d1QQs8N04r4E4vaQZ4IA3smQwmw4rsg8fV
fVBjLZebGRJyjIyyr/F1Dn4BIQJDYHV5snmB1hTdP9iixZmOs8I2NxxkJhbeyhqwI8lkdBa4tJIg
SGm1SngrTKbsM/h3yvaiKZJmVI3T9MfNthkZmACyN1A5crgRyCnjvSn1m5t3u+1MUaVTO6W+akA5
+jU1HBWHDXW0ZgIyKs6VOZSl90WRpfrbHYSqPxBqrrUrKI/ARZtByc96rFU1/ZH59tcCxU07cupQ
YaVWm/vjNhIE+6P3M3aFVohFjHG4LjqQIW0N2/mGqliAZ/c3var9SW26wXGZtLcgbja48o3NzKCP
CrtSWE6o6QukD5HWhGkWY/ZrwLrZDQ87BFRb8UPQxbMUTg9CyOW3xYLU8dqcHLqn9R/KyVIfQOwH
D0QabYR3222xrJ1aSRL2XWcTLW5jnFZj+sCMNsKM6ZReHkAm4Va7DizqFeEeTWSrbGbv+DJQkn4t
nozy4QhAtfKTvYz0i38QBMizr+4vrfufUoghj9ffBVP4meGexnwHUTV9CXd5UXtyUrH/uhg8KlnG
fBfv0fo6YJ8PnXuSj2FkesWvi/nV51lc8ganKlPh54eLD7kjPoFhX3nCOEdMk/9dsiSVBE0cuU6B
yg8pGwkSqpOIgEqQGSrHo2OnE0IWsG/8jQaRS5wBzNUOwyWYSYO/g19G324xSHugAWja8d9/JRJ7
Qgwt58To6oz8Zyz4Tfgm6kiQfPfT76axRPV8FC3KXKxwsx9Hn763uEDvxKcs2QoYKJzLG9oIDIu9
9tQPyhZfjtDjpyezGMzJ0XLh2Df7/yjh7IgH8gaNUxsqng4UANnX6qOY0AzS/KQJiaPh7/gl4Nib
b8TybNUms8GYHFZWHmzl/RE9ZFxluGjdSnVFXUpNuh4XhncFnW8P3EGAdp0VXEF3V0SC7BHJp8xb
EMvDCNh4AzSAKyb7HlvKcrGI74Y68xcA/Vn0Jl7Ru04tEXNwdaTHJ0SirshGJIylan8Ntp+C9Fpq
jdkhc+NlfLdDQBeHlHTgeeD6PLAXa4fk6NeWeLtsT3risMKmp0SHMo/c9A/7vDyc61tlDYl/8c6W
gkGhIh027SDOR93+qA0izBRw93XguWGU15/Y+JjLVCNba5KfjKekA9BubM1ROo5wuVoxRB9YftqP
l/5438H+eRL2GzptAMOyR1Qd0I1rW65aVc2Qfok7NLNiwXFKVsq54UygOzXTAp03DxtFAQmDTSnI
7jWEZPZEsubX6vLNtrKRW8XvNzG7F/28FuK7JAPpQcG1wF1xzKCeJ3/331cKzssISXbFuv9oDNYb
orF+JUKbAsB66B+oi6pMdakx1c9VhKzSXVmkhZfkMEDDT1oKBOcR+MEWV1SVI/sn5wUkXDHfAUkb
jtGsedq400L/Cs9CvbZS6lqp1fAZZUJsNGXy9AVZE06PvagWlnjo3/lejlNmrBs+dcDkbCfmNeyr
7HJOt4SN2TzWESGZLV/52+wt3cNyZY6VWedttJZpZAYlk3pjAb9pxabEkZIdjQ4Z8/4GfKjcHOBF
rKG/De1g0pcecFgT1an4vBYx6SrxHDsgHuyaoUt3SToIn6KW4183IO7jLfMLdaEXmVMV+bIIdT9v
VZsalfCA5v7X6WkUzQE2sTFIUt6DHr/WtmwIVZEQMEdL99iEU5fhctWxID2cPAeQopXccJgXiU3X
AOg37aY8MlA2ox4ShjZQy+H6Uy0Ukwxci9blfaYWoIwkKvdr6V1W5ZejYUr9Kjbgz1uQg6Yj4sbh
VYzOGr5Ung7RFkiXxUIPkQiTpbxFobkKfUBr1LwtvnnLw1sNSrPeUJ1OVE4QfEvzgmjs9UQMhCHc
h5ZSjglESFKpcwGIrLQD5dU2owluxmiXvs0XBnejoqRBSBm3E17watp5y/LORM9QdPIPswURYRLK
Vvt4zIvEE+AqHEZHUwYItmLCEcSumFtNVyKHrxisnHa+l4Bk+gERA7ap0SSUpEhGsADwETajHIRQ
ozZfreFW/TrspjCyLNwET7rxNht08VQlT1En/sibFdxPeS9mPEVIjRxpRD3rDqdPVMcvr5xPBhF3
y/g4uLN661kzhUJdEujZLbJBpHzlPq1hHgkDGFOVrCvEeD000Tg8O3fmNCZuW5oZU+2Z50g34vPt
gXYhNMaUmoNHxhn0eETXNbp0r2UVaCXdPjNuVjpuglTPCcaqeBGh76blRMIxyGFnX8/kFLbvKdKO
Pmpoq3kamzAfWgF8A2ufj9W+8PdrMKNqGhwKOXfU+Nc/0K+afuaB0sV5GUX/N2KvoGc6S7i00hD9
LGde3zUds3L1xLXOYcMpyDBAQFTXDn2qfNcra9IUR+4yjimgBcX4GhhSjtM2MHK7MjNCpBbQ9JX6
2WluIqcaOmhrFgzN++1a6aA7/oJNHGVPkSqQJIN22nacIBi/oUrETFa5f3XF6wuh674Um2b9XgVq
rlDyP0RtHINT6Vy1xTi1DCHhqHs8PzgaTtimmFI5M0Pvd25XAs70bzWc3Qs5eu0ds08ZWJDTAebq
vctJFxq/w6QrLdwgryks9bKI5Rrwrvw6RFHicYYyV2YYLyVqbq4bsNVj4VH2UfNe5wXSnHdcEeVO
SepJCgA+a5hZvH22SX07mxO6o/Uxkbazl2MCul9TC/sE9TTutXa1XJp+ccemAHC9UgG+J0X5rpK4
fSxR9wzbXtBolrW+5wg1qK6UUFJVpTZ7L22j5KiCXSRFGYeHiv0juTj4w5SS3Np4doF67JwqAibO
+1VRDkCZDUVMjLfMmxgQSCe60ZzZloHxj2gp/CRAbBy1Tr7OQzR+oZqzSUNV7wklHdHotl54wrMi
dDvgtGPpYhkpo7n6kXyT96IaawmmTvKfjzmbM6iQI9zJ6YN6Xh/uPoRVqcl30J7VdA/1S7iK01PP
8/RsoxHi8Gu//0IjvUAh6gqxw2uaT6/xxVJ1QmaRXIB2sqYc1zQh5eYw7fftyDu3aigwUMsQ3pQn
k7QNRHTGF/7zdt45b29ufuIewj4NcxU64y5sUIjhaiQpxuv9jPq5UZSRnRAjGE0/kI7s6twJ4GWk
KSDpZlJA0GhsKn/D3FNckbL0dS9nvfGCUNlvUgPNKDDl8pUqa2OvuxMyQboJ1pqYpbRF+ivc3zF1
YGIz4BREU1m8REEScuamNVPeU1o2cBdq+8kmIjzBPa9iOFoK5qIlQwibcYvIlpjafoyTr7Mk3AF2
KiXUSJKFg/6HK4TDxOx1Mv/Dx8167+lbK8FFYi+st9CCZ9JpzcjboBfryVUK3lK0fWK8xR1gadPT
iaW913X4gs/qYJXeCwADFDUqtPXm57ZDhvkTmXTvMKayPgHqrAF+KmOEhNsHLFa/a19/IIzgri/r
0x4MuPxRWvNag/heAxoTf7POW9KjjHBTRylfEHZ7S4vGRgwpx0seL2HTid3v3ORmx5//pKtVeO29
mkGrdIpzHqaxHD6pHz1lHGJUqNmOma0dQ55n1HcC95DTWM8wNg+hv17qAHnhMUqJZoAl4QnmHOoV
FeKYAakyHxZBv8e8skZQzJuDxUy3WZdC9k5XoNAoaeQH+FJtX79wVSvycUcAj/xyUs/X8BkRNO/p
PkvG1FooOL59nCVv9/b8PeajLjcDt2AdRAfAim5S3WF7RI64EIaZvMtT5VrMu+I+n6079OVfrkKX
Iq6F5VIZaSJ1gwvLAj4hhlGiFwP4voJbLGPOXVdp+6nkRUFh+uP3GEAS8+/3nHpXArvGoa4+SeQr
jhZTssWr+sLSntVmg9p27ftjPj8IE0rUajY0K+I+LY7QywALRR0FqpP20Fn7CBudU19NF6w4aXeH
JVVzX0SAFcVpasHdQub3dNaNnKvzxQs4+JbJ2q1n2Qcii3qWTvqE8pSy8qtbNPqF/zkPZHdi+8wj
pyUYxccCwUP2+FzFOVF3OHNbBX6HUA2NF7v7mxWLVd36/tEUpueWpqspklynMWZi2pOSPucCxb7R
HqBd7T7E0x3YrfvBRKbset9uGB+sK30TLLxW/89NjVBLE3j5tr5my8Ej41szGsOqwNXDjQoH7xtz
i8EB6yNSznVEdC2qNOTTzmU6qDmXyn5SlBmL8iIx/3P0bNXOVXLBoJHgyqpEtB8OC4Amoq6Lx4Fr
gp1kmUxteabbgChxbNnCiZMqoq2fDBScSh4ruhvjqN3xl7JZ7Pez8KE+kGd4YxMoLMECSBX5m/eK
MB8BDKfJUI5vlgnCmn0Ni4aXrA8+/BHxkxNvC29lkxN/d9Py3OboKSBhqe7+EDIwNN7q9kSo3E0k
NsMaLoM6R6/AdPhqoalco8AL9/hNg9E9ewh7I1IZpPijN0i0M0pxo3FncpNaWW8+eXm0cxbc8M4B
es0O3EKHHz+9PFA+7dOAqyItATuisAEUuqlIGGeFqTpwNBPYYX6JPUuMGRnQOQ3lTr0F83vWhCBg
RfwFCLv+gnjAxCBFncLD1GlfC6ofw7P3U7TAQKPX+4EstoWC2xBXidtTG3CnMJ938/viRzUqGkov
7xah0F0DpuRdevNnCTr0QZjYps7tBmuJfHKvO5osNehrCAXR5PdyYEtTUrZFdwQjvjXQ3lC1k2+2
TNj/Wdol7gPUoALOfDyhmz0vwsjDxcQUjcp5Q9YXFqOBBG876ljj1/tq0EtVQNX0xdQiZawouYPY
2vuI/w224Xnl62NvsXCq7ZKJ1ru9qWJisLPQpqJSKL6PoGTRPXeFZUGFdxAtTCbb9ox73Hbgzf6W
8dDPABkMb8L/S+mAVLqlbZsqYJ0sgg/mY0wF2+pVqgWIfpudmPsA7BpeRJc/OBl6WArtA0Y3SFkv
v1OqdGMBXH/3hfj9GMSFJlxPA7SWIWSlWFgJhVsC0Wt1DnGYd76iqZoxYfxn1NxkrOipFOyw1Lar
P3SR7avm00w55aDqLpSQLg3uYY6mDmNPUFkdldV1OrFVtTtIkGErD2/p2SE3LJ6EvZaMnHBu3koX
NOCFJeWR8BbQhUma1+YHFOvlJXEGTpIsggOWzlukAIt+2dMTEbFkNK1LSed7qCMqYFaKNAUrTolc
P2KI80yXOwj2L+m05lAVIjn2Jsx7AugmRFI4MuYOXCy2IotHQuuwzlrPQOdcn3Gcb9sCNH0qTSm8
LtNEFQrah8FqKi+nbD21od/UQtbwlye5s3A1L99bHPLS1DW7F9qt2tOUo5ohzETXAIHViqLGbeVc
fb0zDX73Uwm6NNdXoK/86s3ZRnEgYGz5Kc1HdZnomBV/Fj+li1AWW2W/FQhKp3D1GRsBB9Pk/msy
eK26VFhCFwpTG7/uz5aY27NR02lhFwV2Gykd1M2STFvZyOlEm/bviKLacZVRycKoYh5JJTCnWhSK
AU09g4foJtkNlfHHZXGuICQq6N3Ax6rEaA89aXBjxVm0UqQv3xrUJFRz0ekpN61JBV1UQKcxPuSG
oM+WCIVflAAg7P00YE+ZVL6TDQ5gKMWJxsvfcCLq/nGLKQ1IwUGdiCTZisbb/DTQIlUuEQde/du2
2Nqh2gkguJolCoCoRuEHpAn/rAVKBl4WiXqmzGyC92VXQHBIhFSNQxRBIaXhdrHuwUjOIyzdMKdu
e0NSuAvr7NGBWpIwXuGVqZokQEsXWoXwKk+tNxEB3F/TIC//Ja2DDv/LhzAf7p/79dOKoRoBERH2
mTD4/L2JlOqA1mZkls3pfDzYUjlO52S7SzjWffOwGEoOwxC5XJVNfF9FHa4NMBmQY0mceYsLZY9D
fe+Z4JLoVx6raotszDupIIEbAtKsYsyjaRxwc0YMQCbDrfIMNtITWojZFwd/CzoV0MXBBxSQifLa
5na9ymp3R2ZGU/phED+xtEjgZVBksaFn0RirD2ZLMiuWQnH6gjDmQJP3ly9We2mMRiN/2GV3vVXr
PQOcint+jU1JyCci2Xe0JHb9m9GhpyCQP0nfs2/gWtpiEZO6PauoIHOYrOEkBLRt6Z6xFTiLPBgD
UjOCf/reXCzaI0REHzChTo/ao1h00ns+XOPGLpPfiAM4M3vUdR3J2yeqQn7ZDqMXaek8wn7mFmiz
2knQGjBwIVnI8FUxAxZcKmTBCF4IesuqrCoXIBYW+Wpr2wpbOazy9GJdpP0G4tx7zY8NJObydE4k
oxVh0fXKuV1ZcmKUpVovEznr66j9Prp4esBevTzCpTTYZ2vtgzT1Igo38Jc1+yS8w8lcKr+cQnVd
GcJCf0sxS9qC9OFm294tPtifRgrS9pGHrDAzOpVx8F9sZg9UTtSOXcZFV59OA4P049tTPCGKE57N
SzD0NUZMio/xqZI7HYdbWOEJ6M7WLyg7t7awQFLd3KKetUO+Nu7xRfJluJAO30sXl+auJ6toh8uX
gR3S510wf4L2t7OQq3pmBzdSrQh6UKoZ9KS/1okupElG0DgCe0a0pwzJcKM7yyERPIJQ48urGjQO
WmPqDS0Oh/mx1RHlRG9OrfDk2oloDxKj1hubzzy5et3ueoHtMZFO+/c0L6uZH31lBv6UOrS3FkEP
oHv9m1d1LISxT+dUBXgAM5HXKp6bFpcDwZj1+nG7V9xW2F3gi6nsLoX//pUyc8X/cM5CyAxtOcvQ
646iyXR/fO6BUKKnmujwRggF2LSePerJsVoAk973wphV4k48fg833RXibdjy4E96BKXG0ZBYZ8Cc
fU8CuN08+l9fEr8jCIlLx88GDD9yCn/hXlnyi04l1Ev6LUXLCWxJLnl6YK0H0f9sP4WOxGhoYeou
xfC99QmBFE+nRDXA620vLrXwxaty0+4dKxXqfub7Fraz1VDofXvj1Ix4RsikUDYeqwSK/cAPFoDO
czWy2yUwPTwDAa0PWj840KT7Jaqdc9PSaIvEoNuhGw8ejrSNVFQOMSNSG9TdLbb3ZmDw8DCntfz9
J//v3pS2O5BzuzmVHJ50kB+j9RdZ9RlAZr0yS/9lf1P8JsT1iAX/15ypVken/sCwmnSHSEbD9d1T
zAW0CLu5q1KN+o/a7jGupqDznXfmdneXO7dY40UvDB3fhwmXLZkBNwcJWcxIhbpmn4eQlrY/bh0N
d234NYB/ZOc98WGke3YxOcdK2cAVLifhB30raIzpzy1ci24pz1kLnqx3uh7fZYN3hR3o4VvnkYF7
jnz3g1WDajvD4TyV+o7ZEZHhsnA5T4APG5yVeiDJ4MPXkV8rhoicesF4xW5NcaeooTlILGl5IjAx
wtXwTdPmMhABIgxS4p/djVlhfszR4eDlxc84M8+OIdzZT93fN1PjZCz5ujoPuRoi97Z02vAms4fQ
3H6q7FAYQ/pbqQAVUhAuxVRw2mqdc1ql6uH/bicgABzqKIRDte/1IajMNe6NU1YKNzGv37MRyXvK
ejtmYTE6xEEFTdp3ircLzvYZUasSlVx2ZZYQ+BFF4FSLApcVi9aTpONOqPX+wnu3+PB4FLTtWc7D
btfz69T44XTBX014Fq89hGvoMfOvllitYhGvpZz3SJypLfb/Fpj7ObsimNYbjNUBGc7nLbQfL3rJ
o7k7nPF/8q7QXXdRAoqK1LBD264UVJfAoSJsYg7BBFgY/ACQhlXRpSN9E6bEL+TXUPl3uk9H0mzA
xnEHYrohDozfFzQzQHFWTHerlARgernwU/HqNmH1A4nf3ljzRFxONac+Mofvo91EnivHmd5nLlWf
4IclCYoNxYuxtUpFLzxMQioYDJIczBxUaP+AwdWCDMpLSp2um++nGj0EfMk9HBF79/jRbcc46bB6
+rTQS+K+DMplkFOEXRAC/8QGomxurt2QN2AL+hcX1X8WdKfc3WVjOVQonVMFoaiUQ2N7EvmV+lxb
KXBIM3vw4qBKiWjwcjq8PuWkb9Y9yCa1wHqiXIMlmIb54x8CkmmtHtzgDLWr6YwfAnf1BLYZq7El
lFWZvUhfgfrbyi/y+txaNO+kFLQZIPXx86hyN11W+T1WU3KcNlmPijlujLXkLaObBG88qrd51TQ6
HASDYgo9zaC0OY6GZzxTvoqlW3ysAPFjDKkMen+gLga8SFfc2qDCmTv3wwU2soTZqArkGVWkw5/s
StI3dcB/kf1EKHYSi+SYDWV9P7Nl+fkmjRuRunQxg1jkPTZewO2E+b7L29fXFSCQ3FtNp7xuN1+d
/8+0afOjilTk6KlHUQ4zkKze5tgfsMV2qdmp1Uo2HEYqEBmgItSi/RTws0wPyBq23ZnXSTXZ8rMe
t+xXWg8LjeOHGcQd6jKp98GCjuCSLNYN9HaSHcNXt1sM/ik6PUMM9R4MsXnH1PwTHx9179UlmRLj
u711PApQ+WA5cJpf7jGHI/PhVUmAnbLu1iUAW45Ug+HmQTz+VANdxLNXLmb6rAKXiaF8NBjdR+d0
6luuQnVmAG72lI1Ty1oSf22PNsk2jD62nU1KSzcrazLBJ6OnsZWsDBrhy5/JKsHxtIUZNJdhH36I
4fC5IlIeYdHwGFR55FqasuFCRxfPd/JIzTPpsOjXu4KY0HXxM30i0T+kzIJ3bkG6dgJE14PTPGbQ
+GpyhA7P33Q/2Wg8hucT78/NqYV2k2trg6kn4z2e78+c1TBVpjsBnTEUnW3UP9b5xUV2fUUn1XIR
rRkFLcjlEYv1RtAaIl0K1LzvYBd/9TnNwAb/WPTSykH9F3TwVsVB+cnh5qdj8a2V6c9FIMwpguNm
NnRdjhSJyT/lpd+yOcC9rfqUXrh920gL1l/NGmpTYS6r8fw7JAoQP7SEJBkGJdr5h0qpMtb//kmd
cZSguQG0yudJMojDcHlucjJOKEa/P3tyROM29VLXsPeiB92RqEEbZIwEwpidjPhxKTdlqoG/9pcK
FpNg26DlD7yrch3xKrp3ITQWZEPWZBZlnn6DlFb5wb9JAn5BFC2ADs8hnaADFZDL9X8AB0brwC8A
7w+9zcSKNUYwId8cUqvHli9vLRvVf9UfXetCcsGUnHmALIxSyli/Zs5SEzwtHV1phW10kKzqrHQd
B16CqmYvuoH647oOP78PHPpEYAREPYx6kbx9/D9FWk0+L4h7Sw7q53e7lt7ZDITRWLx0ec5CE+XP
HVXaFDeXKt+Jfk60kNdnjHcAJnqqIdxbU7kmnLHF8O7DN1uTQ0BSPIzfBhxXe6W6bJmc7GU5aTA0
DglmUHKOmnxFp3yorR52llr5xgdPwqohIiFA2BlG44Jb9F2Y13LWFjl1gJ67TYFeOE/Ylaa6Ii2h
ms/Ksl8EpqBpijo49eF7DvCZKGhBZNsGjb8RUY8qNgC1nV+evUhzcWz+eH+N/8Ifdx+/BV/UayUt
xexYDT4OCx5EAxF3jP0hQxhzBpl1FcAzmYhUg0LGTr2sbgZh7nZtgn+bKTGMznj4KEg1gugSoeNN
aRSbUZ/4VKRLfd+b6ITlEsPHNzORT0Iw45BL25aqiy+ybw0yT+jtNCRa35+JnDLkjtdREdZ8UGNl
CnQCatfsTdJC5sDi0DwwW+bNENOKWvkwsv2GBw+DQXI2f4vh4Ub/BDW17fCTitVmIvrG8y3/vmQ1
eS7x3ZeJkJE6S269Op2L0AJ2715wuIvbjmjHpMS8SuTYSvR1u0S23fHUXQglKkxo84/ExipvDQIU
GdtF5y1KjjrqG1hVz4yAmR7YTJBHxBxVY/xILTckjiWivxMOfIq/EU5PgfSGZ0ovjmu/QeLs8mJV
OEAcbM80wX/+7is6qlYAy2pH2dc9N2giu9GNLbw4TgQIREFNWDkv+sQCbnz+IDMYC+xL4GlaFUdF
TnYw9SoBj9c7YEXejv63UHuxzQ+Au0mEqXa+/CdM4AoRB56UmvCTrub9IDWGpVtyJPU2xR9lLkMs
FjvijlVAEQThWY/CxtBDKQ3oVPL04gXLVh97fV/40zuAZKv4ZAc20jszI19RzC5AQY0TOBgj7XSM
9Tf8xDFiiAtiY250uebuKUgJP3hdwGt/+MZeuNrkTOMnyhSnqV3DCCMo5cpn6RsEGEhxKJOePQdT
PpoS5gwRq4ht6GsF12NWav7vciSwfhs2kSWJsf9ukpnBKHusc6QzT0zEw7Px0klTkZcjCkz9rZoq
yxcJJ9yiWHxYSSuutc4zQM1NQ4GnR0ndpJs4VDu59kJf2vx3vHrXhADRB55r3j/AH+VRjSnehQll
CQaOZqpimaYA2/j/YsLzyEsJLxRHGGmNtEnVxe2ZxSKSSCkHA+DlOgB3uqzm06IcmDp/NB4oU0Dt
Ai44tSgu2djRVZNC1oYVz5dWjDoRPfGUe/EwDU9Xij2mNvPwy+x67yGxyXxfY7ZKV20oEL7/IuhU
P4nunehaMaGa3QpTf+faY/BD09iFD7E1KwStW1zpiQQcnpYhpzcLu5w5MFcQfFwnZb9cuP3ymJt3
d0zqVpFCQEvHXG+Q8orru40MukbYk3vSLS6kFDawi+OOrxI6ZJrnket7FRthWkdi119Q0RYk6GiA
eFmB5RKW4flD977MSMLYVuU0PXawKMM5k3eOsbysnsEHdwOB7JK4hwz7JQm8FZZdOr2R63AyJqdt
So0H6BaXhiqpEdGfMPKnQxkJBYfMLffcurUmkqanUGwQW9gFnCpATSeKp/sgBtyp4y9XBPq6vyCe
Ou6wlhll/sScBRqpED/pccKDdACbeqCcAPaJtxjsO+w9biP3ysC91R7ojthd8wQcPlwspnUTVrpg
vog+iQGf6iHZ3AJA10nxMJtnCLERPM2HUVh80NrZSoHV+pdkUSZUBHsbkIKoLXHKzeaGBYCvi1Vh
UXR4tQwQBoQBaNBc7sNzC6lBKXkQ4TQyc7I6gMoIbU5mk0t1SBwS70m0S/6Pr7PzQO+x1NeT7J1B
9sGVhMzmdHovbD1vaNDYLGBPtDUEmDBQtLkG6K4VipFPJ/0NY26vLLtZKM+Pf2JxSEsRUDMIbYth
BQd3TWlKJOt/qLDM78UWNuOUsszhZ/oxZ0RdWr+r+NalDhvj55Zy0dVMAtrUqVC529G8paaaWU3n
r6bXaUnnCngX3wldCDiEZTdPhk0z0srvms0wZdCq8jIcUo2k//pJNO204YeyExNvvvHZY+RaGMRI
UCf09v6cczZ+W6jhUis62xVZg7D/+9azrnRDbezuI9oUWMDUACQ8aDp1NM5VbC2x8Q6k0VoVnCJl
MUypuRXnesxse8lK/+6+kR64uUnj/vnKd1Qn21GXzohBYh8OlxTOxS9CBG1/S4UlV1FxnkOUG7Kq
33IGNadOSaNmsy8hO6dX98r/r6rZFpLc8dFShGRifiSdhBenVwkPKA6wxJB9c4ULpNStvUATXeB0
UHiuOObn2zz3ysiN+8POQcN1OAMDNT1mVEI6z2rhdIf70LOyTn/P3A8aEfm6mmiNtd+cODczemy9
8PWnLvpoAcobn7vCStVqifuAcJg++ACZn5XhDdnzT/EhCuSsRvc9aSdjleJXy7vGvztr2nwIdMBZ
w4qt1dK8RuzzKzP+taa2k52TEcLHRwRrU99E2axYrkzyKQnRfzcMEMteld5oHA6C0sFBp5JBy8Hq
cWD9+ueqg5tZKAZjs3vakv/hP3ZR7PPQOsPoHsMRHX/dKVoFvfIHLoz/DMvMwUcGLV2bVtQuJmU8
9dQfXf5yS0XwCbautI4paOQavquypT6eqjAHdNr618YuZJkZvFAQnb2h7KVO4zNx5Dch44ZqkzE/
zwYTJuqgaREkA0BnEY/JgxYj7GvC3spVR3QVwn4XeRscLev29soAXeNXQhnDHiFLHYwEjkxLxLlG
qppPPN+0f8wWLUBKML4YuXEurD3qYua6YlSS4gL4uIe7Kl1YFQ2P3nTmBWHLOnJSpLf8R0Clhikj
B5t1VS8JUCQG5+OI13K/mX3vuF1j7WJmqwyv9WKetpIHaGMW4Q2eTcrwf7V28ZwViKX+wBxJsI4D
jJeTBBk0OiN3+T+fU+3eI0VET3ApEsprOmQX6BI8WLMG4oJCIiZkimbaF9g1F8ENhMaK9CAYxdZY
1R4nHcwO17yB9uvcUNl1FRleXULwF7iT9DBAzbjgV0IFlLyPMp//SK+9Bki5anlx0d/KX0CK9bLb
XhWNvdd9iD1Rni18WoMOnBZR2FnNhdVjGxHw/gzTxZ/af+ijVlFvYoh3U35NIzNgsv2qAZPUcLZA
S6OBrm2e5upzXCebxddjcgrfwSJD+4bGdSzCDIVETuVcxOiCFFn90NQAvECY1EzotWnRoZalD9/Y
gqMGc6mbz71RYD7iurSFss47JNaM0ir7cBHNIAp3L4ynu+NmU+noT+TeDGp/JEXdT2yFIsGoLo+5
lEhWZ3BlYdm7eoq7HmYVzYp2KaHnSgqx2+qTH20y76+bSugSlI7OiCu+KD7/0WQBsKg4Rm7zwq6q
Ju81aH0JV1eZATsiI+srOXM4CJgzb0teLw7MCuXnFsHO+as6uh5q26eM52EIwFb9icp8+a7o6j5R
E5OdR/DFOnO9aor8a5e/YdFcqg+mmnsaCZMiM37DEMkRHryPiC9AogXCQMxrMs4xIj5lgIX8EpIl
05hxfekc0K7q6kmgAtCtijn8xYmguSS5w9R/nYPB4X7aGBsXgOxdckue7NhI2whYLv2SCn0rgL0U
e+fs7fLXO6lHZIJMvzZ3ZhMnVx3G2U8XkVOQUN4AQT3Vo8LAPtvw02a7T/aFFklOB3WcaSod3lmM
T4G4yhGiXhvgLDz+MfYo/CKWQVEZhrNJ1B74rhyeoX3r59fFglzzF/O6gC+VXl0JBxbNjrKrA909
bU1xbR85qZUHhoC5H2AmpHr3l/8FebEoEnDEsKEUsEOFkf9R3Zf+laRw/QLhXOW6+FHdOTcnqMK/
RijccxqopPqibxLjg0qnIwiDbxaovDIWIk5Kdx45dVlV2iF9zNbZQQHDi8En5l/hsiPDwSDRyd9f
gCRnciTUekpiRr35jkNRjfIfzGJ5t9fEb9vlwMqMPLbqfcfPNliiohMSR1TF7LbnuxNu7d4F3lJK
DyZhfd9wzRRChQiMCW2aHCUBqIcP45LQMbCKA2Oa+4TcAolL1z26Z/Za4SER4Jp6CVW5z7EwHHvD
mfTZIIjaFO1pjCp7g+nY7w9dhXeyFGsLYYU5wNy3BMwFrjrwBgwk+toN0+iP0kgfFFvT8BVXGA9L
kXSGJJiyJJhMEodl0lI107Ax/redzZjEMTYbAw0oQMZ+E+NDZb6EkPbxF3cF36qU9b8iu68vmbGa
b4yTh1JxMEC7bMqK7Y/T1/GdkucWNsmbgQNkp3NZwTKay9R/OL4DJJ/Ehen4SfB52xwnzKEVr5Or
F5Ei/s7CQ5HYAVFTtF/1WlQviYHSv7tKa5k60tIEJgd5qEr5gijJGZO7C/B0Va/3qUJh6QOisF+q
izC66JXXueAYrtJl9SNs/Ms+8E+R3zB6XhptQHmWZiBspdIOP7aI2IJD9492JimJtkMLtOq+7GaJ
sLyRH9ef4KighXYLLMb3KQzBPZgo0OtKqCRBxRAzAvSpC8z8if4v7K2/66VuRke+AKn+43xDZbO/
oc5gN9gDQLi8ra98R5ScxT05+y14wf0n3WyTG+gRUvQBw7CQfkyyYR+OpzujOE4ieBwuhdZHNc0I
YM3y407YWs0h3gDkAnYC5JxvSBsAq5BM/IWDnCTXKH98EkJwbqq5Zuo+omBCDzMjLHwSkWGxS3Y8
YsHPpP1i4AUXau5TwtG+JYTE8owKolTisrNr2mDldFrCKyS/sBcFAsC4/rC+qRwFwnpaOhShmjRG
a4gu+lk4P/I5LuaytlLiJaPtaG+wEePfhhAZ4kvl4nkp7RZJ/APdRfeqxfxxlovmVP1JbIfpvMUT
5au3HjNckDmRo4ac7Tpliv995ln7ljyrcWCaEKyCrCc1eAvlYzkSjjKEjqcxNQnxXyUcXHgcKBHz
a7BzAnsoXo6rIAwANnUaKiMuXXZkQGg1M0CSOqkBgV2snHf5oil3ItacWd/kZKiJ0Fr+l31V158H
wQ8lIAt6PK5m40mElFm8OPHSiz+V1ZQMdFQAr0gGeDWZgvxIgPPy6hosYnGGlcC9JRYRgB7Ku/sR
VlSxKXymFheF3xPfnnYabf0K4aoHlnQ5uaYV88ZuDwLdunET/99R1voLfaYg/zaEkcAr6bWrJnWh
H+Et+noJ2IlcHbn5I88k86wh2tgO9boiP2eBR7VThRkuDJyCDyaBuDezWQ+FVQiqL0APw+0V72/p
acr9+IzZU9CmolCm1HOLUGEqIHB82mHs5Om4Og5Sjoc6Koc+eDqv1OIRJxQ8Aq+Rc5U082IH5U1Y
Mh+ld4s1ln58KcI/o3i7V4RpsBe+L/ZHpJAs6ILFvSM4Ut8/X/GtKEeMY0FOoPvjKwJw75AwShyb
lWxqKqPbuD2IGSIFPW4m/K5FSpJwTMjDWVJ+zuANEqQlAZm5mi6FxlWEH99ILv1J5GDP6ljC1ia4
1eaW3Hh6dCC/CMJxmRJoBQI0WUTENv9G4DMpoaU7xL+8bHWtq4FhN40Fy27ZPS3vVSqgu19Cm72b
LgbTjsUsmHHCVZJHjV5TnTQfvFuL+QIVEJfVD+kyleflJc0M70FEGJeNo2qsAMfRdvF71xE9Wk71
xdB2GpGFzJISDEG86O21IH/+k54FnbR2EQYo0IyyI8QUSQoF1efnZfrPMt2UCXlpgc/DoOE8B/dk
uN/FbNC56uvwsQXq2WmYQXoAT9g7Eerj8RaA3wZa+SlgF3iO5Fq0jhgfCypxBEYDW7lAdqYG8Hdr
s7HEx7Wbc26pPul6mhnmoybtRrdIvDQ24f8s/uRLHxRQcybheAv8aEzgqS5q9UqX5VBOm6qX3Z5Z
4GPJGOtJaSDd/dDua80yen6pg/V/zXrgTL73ee1VoBkrTntx1+qDrKO1dbdd0RVVf3Jop3Xvp4WS
+9QHqVCQ+WrqmIWiLmjTVXmuNMLk0e1j7eHpi3MpXfIEgNHgh1m1zl3gueHYFXvv9skn1r1LtPXz
0Uqdu+FUonOrg+KKU8Gu/KbPBIen0woU67fNxv9o0L4uev/qTVxL9I5R9W9EfV5mRV88eRNp4Ny7
pys5Na3eu7eWAlOMDGBbGH6uRpDK1qGL3LFWfHqFw4T+EGFiA7QPuH97tUogwirQVldBEPVPa0YV
LRaV3DS61aoxcoyLypzvERzxmhui1cm1TfjZoOC7SXPQza81HGjrJir3BI3NJpjwA+LIwP/OYPZ5
YJDdj4AeZT3ORFouimxw42vJtosd1DVZh+yzXp6x27vye533Tfyi6lk5wEeKaLwyiCq4HKhLwEXD
vQWFN+6+1QsFLAqo+dz1gfoG/yCtAPupIwoGBus99ZwAz2laHOJPOkTYd3fq+vGF/BNh1bpcLFxn
6uyvoqBbkg5EWu3vLG8M7ZCu/lrl5URQoWPB5MY9GlIKx3irO4R8Cm2Qn+gskOfRhduiYDaKWgxC
muDGMFr3IZg6QWIYFbSskxl8EOcjiyzjb8LhuRCQmGK2Ogg01bYkh7r1RG2vm92HNjUxOpmkmoWs
mt7dsnCQ84zPwKAwX4FVMy6cqm/RIXA2CGRIvbs0JRZ5GxMDNRQYy6R7kliu1GOJQ7kM+3uRJ5j9
Wkz/ID4g8FkHWdqljeSIyzgaDEK8GYDCnFDz10p1B5UXwGO5myFnt/ZzwJWEBbewHaOdu7hYI/7A
pbsIueQZzUsdugyuYwUJSyqhXYAbK3hkMItkUf96DgRbYa2l//1uH0tPBI27pMsc3B03Pbl7Pvyg
VeF8zyDxwscpZO0e/bYrEXMyHf4ClufqzHoPGtoLjbU40fEBdoR+LA1ej3HrEWO3J8Wnk5DyM0tv
ZMAO0CKooHua+0/KhYqhgPzVJ2f9l10y2QPCDzVdsa3re5fKErQBbsACRzSA7yQ2wVHbX5L9oTN7
Wb6IAQYvJX8r3/DOWpHNcI9bkRpkB0iO9ceOGA2MatmTYpz+mWO0EklBVpG1E8Isko3oC4SYBANf
L/XGKhbcqZuNKlWzI0z6DjX38QZYiktjPDAk2+s7rsUXg66mKSy9CrhBVlteWd8cK/ERRikswnxH
Aknaaze/OSrTCMKDVQmUGUDPAIX+PH37UShJ3MSUUfudLYewrY4DwuUbJcea3WoPOkzRLxfXbQMx
5nC+IJuFMRt0GjLt96Rel5VzT7aIe5MJjRBiHjSoli0CGYkdaD6CApEMzcBe+dLruoX/HTLasHHu
eqkxbEZUzDNmKcDB3nKQgkdfNzh6E54Rbcer7SLnIVyEXl3ma3ZkX7de6o1KcSgXAYkOlnWLvRWs
BOjALAglIqGcXs5BacQ4aClolLntdukz0lFdNZsJ54EZJQZu6Avves51ANifWsfY9raJg19hNHDO
i0ZOp9hLZaU0/uDriYDs5bO7I/4kbpjx4faCXXQP9W+sss3g9KjixxII0GWjpXSJCaPajFatAPtJ
7wwW40hmgknjlIQsnQlFloTqf4amn3m9HN+yELR6rkv+Hok/Tsw66nkTRKsvvp07REq5PlalQFX6
7yALoL0LmyKVNWRzftQBH+4GRzP5Y7DmSku04tLqX8SXn1nckVjiP+WdH2JlkSaSpXqDDtVIOJLn
rBx/K8BkH3NcflW2nwiNLdo5tR6PPUNQW+b3eCitPBCvI9lcqMHpB1aJA/zOKd/stR+O+JQE1DU8
w3j8zdGXhI0OmO9rh5RwoKH0q8DInB0W6nuBXj9urJJ924B3cxQks2LKW9oXvXtNO0Do7Q+1d4Hw
jt5UxwekMMo0Gng3nheS37IcbE9WRgRb7x38F0UA6bQnvXa/B7wvHO3oS8iybsMS2BjkHidnTTzt
kWCATW0CbTkcPZwRH14ac97rzy0yJ31tYt2qqKqEU3yQcclo+u9U6DLqd16Uzo62IarMDa/pmqJG
7bEWJW9BfXaTst6ev65P2FCY2wl/4IZapv1Q6kvvz7m7HnpodAjLmp+UqXI3icUD1RoBZA/6komE
/5n1imNoR8BEMgjF7AGaXPL4c7MgHgoX7qPzYpDLT6vM+KlkwpdQidoEqC7F5fmhv197Gh4/e+gu
CS2Uk3HnStxCkEigjMLmEBDX6qDdK/vqcQsuKMaXxQCF24pRoU4d8fI2qFmNbaX+x7G7CzX89yXd
K6zWy4wIqCL2OkoSabPNVoUuByNr29pf295x4/sAU8OT33C/tFsYYq/jiyp3+omZ3uKGO0vL8BZm
mQlWTIS6FXXlRNCIi3N/fOnvVEOP6/d7ycWs4Hqs0P0LoKFwMbG4lfKz3ts46OPQzhnbopRVXEu5
QIjbR8drQY5ofFohW4JlrD1OWKwQw7DquMmpZQiRlFGBZWIdWKxo9fT0HWTtLGuqt1XRmiLnWpia
h0EnPAu9tLBzWeUl6Vuu/vGeyDQ60lhlNTASvRaQZDTgrdTXIhuoA2BEP+tIYuZDSkdJs1nNCQ/q
XxN/yVaWcV5fX6RAnChVnUbeWUIv3mHUl/AVPw7MpVzthrT4bBb8cy7/MR7Nc+NU0W2a/E2cotFU
2gkyPgZ4CDehUJiAGZe8UJ/tak8lG2nPLGuNeB+8z6VWdTrWpkFwcCmrY68CCzI/g5yVYzOL8+Fa
6n2AZUs80oNbJMc+bLaOIxMWoAeUWoW52RB68LGPtiAkx6i/H+Z1MEd1SOV65MBhBp8gk9G1RYVr
2DKMG5xo6Rfd8lsEI1z7MpVLm/7Pqa98A7NSAjc3yREFmNmRJegECFmXGNvdBaUL/TSun/npERc/
kAhL+1pKe53SY43hKW/+dyB1pKcg77sHcidFTOMvXCygQ46pBYQTeRQP9gDuXZ9tTNZBcJo4ZCTn
J6nB9UeZncEwQNuAKeYswJJ19JkiEAsBaI+wGalCJ1TtN+gX1M55lQIu45kdfdHY0iFZ2eBnzCAA
yOoszV4osY0Aj4t/sF+53f9t2ptMm3agqZ7j00BF2PkLwS8RPIoGRkbaVQpX+IegCEJ1TrpNFeUc
6OZTVdnTrRZP/09mezLH2mJXDfCZ1al2mk+hh1MuXkS+Rzp76cDe6fKlOgh5oZnZVwZW+uu60K9A
RYUghKR7lqDccjILWksi0pW2/aHHr3SAR9nJvKkxzbPJ78MSIip4Zm4l7bU8yDOi2VWs1f5QLOBn
xvg4UROPImfcYZTLfsYFmA/P+34Hmklos1ohgKHg5GCuEOWhYefHkP/VISu6aRb3NgkA5L1fN0Yr
tFahfFc98y6KOebSyLJbtD6zV0aXyH78xmfeVUk5fjktezSob5uHFTxVyt1N+cHlzL52Isg9U+TM
oNXvJuKXmOm6Sned7zR1oq2ntgX/zG9wAVjhJOSzQenoIBhq4x8MLRzxnCXXQ4Fn3sdm0B2+9PIJ
4OQH8xixUohjRJx8XrTlRgIf2XJ7bJx2U+mVAhrV2mfuJ70pUtuELP1/P++jhYZiUgNgs0bDwBui
6G/eGcXg7bOBZWBS6h7CJEIJnzMVoK4fzPfU/dFhGV1fNn7r5lZqsTcPwFLSfVaUOUFzjN76h1CN
B/u6vIs2B0OeeqZrf2xoTrisdUsOMci+GasoqU3PcO8lzPf1h4tkTZCX8IUIet0+R/vWpnmJnVJX
d9HtAB9Lb+s1h2us80LzGAELKTfAdHpfs9x5E2ZRJSpLBlDCfa1Jbz4Lt4CVxv8Xl0rCczCxWEcp
RpOwVWlznggTF6mZESZbFhRGysOJgXN9O6jJn36kHW2+5604UXWTmBKdzwiChgup4O3RY3XlNicC
KIxOihanGc5UjDvNAj484MiHDaAo0WoDS+QI3Jlzm6OB3FrNPqnBMKyZyxXv4K2a/o4rw1vVXU4n
M6cT8j4UobLN101YtIyf7zSyHhMJBizFG72L8wzD6WYJ5GXuq8PssV5S4UJWFpV8IruUnOLRxMQl
4G26LeVhFItajnk/1uwYu+utlr+Qh9Mz/n09iPYen9I8WC9Lx3SGX53SXQzyEsHf7drkBVFoLA88
in8ec69I+tGZRnmW5OxxbCNIiSRkKTmZUtMTxyFQ2WJ6T+DC5umL6QnPrpLniVcQ6qo3MMw+1Qzl
lwe3zzCRoSxzPDH+CHYsR3r7mWcIs+UpA4tzEeHgWiKJL0Xb6SOCQDvIRKIGBBCAkkA1JJJoWVwA
/qVv73c7on2UHkV1HpU70XSXJrRHIbzgWmPOmh0dgZoV/ulMTmsCQgiER8Miq0DCO8gY+BHs/Uvi
j5+XaPIpLvNxR2xLms8RDUYqVMfU4OWcydQ9Kcx3rSucsT07Kp+mv/OLT9YzgSP8sMAgZgcnQA2p
iYDx9Ti4jJPMfWBDEC3aNFF/9sihTp1YYgyEg8DIR6PAhwA1SOX+tpgLjCQ2juHECKwYgrecuYfT
us8R8iuIPeQS8fjdqMvuovhFHQhUh+tsFWbqcQrwXIPemF8LX5cpxCxB/orSJFdkyReTNlfnzm3L
P6CEvT4kGpIIkHOa8VQ2NKvYg+gq1j9f2LnTEAGWZkQbcK0Q8bNVzVAMhALe6jAp59xf8Z/PnRNA
q+8MPqmYH0Xtat53wKuBwkvkv3/EHpWOC9BRInmTF+fRLpOAxU6rLcs5AFSy+y3Zf+xW4ydrIzlD
1imEHlTy1bK09XSb0D1ipl6ww9Iv9tEUpx+BsHLjeDRL2SNVPngJ07PaiO4og1x981oB/SCklb1K
4CQSOQPPInyyvu1v4/TtcXlUieryyG2TH3jrYBMBh6L5YxEGqLB9Dxs7SSSac0XI/xWOYeas/780
nt6dJDRs1aBrgcqpC/tWfKnRkeUx0G/bB46BnG9bvDzFz1sQ/UVNGRQt57XDdxatwPhZ82LHyMFE
qMqYJJyIxhwXsk+6dZLIdBdCAnD/mD7x/uF/OIVzwDvO3SwnElbX93EoiRQT9N6IFJQ/UdPY25qg
ahqYrYqfA+fvxtpiVLM0+IdPOskIcUyd2snXvsfBpMLPUQTIAaR22y6hWp2+Ve75SMTFHJdC5+7v
fOCWPLayhdEKuJC4Kp6q2V/hRVhRcwQpqZ/7qAaDjU8c+ajSJ2FibpxoQalqRn6Az//3Z4DB0VX2
3eHup8GuoGywu8gwZEdqYndYeiJbZXJgRe1Suk7bfhRwPeHiC6sQlUqordQeHeTvSp9awaCQxYbM
UA+m7otprMuJHvOMj+KwEda01Tr/yWT4qX8ogUWH1q3RFSnHEUvdttQdp+70kiKCLcusa9PXKn5u
3SyOMdV/T184eLoyXarbiwXUBCIWWCyThergjQbwFog8ODIDl420VC2VPUlv3mfFU2nAMdmNzVLc
oW06CL60N9kYXbsHz+bbtmWwlbKu6W5VMVnlP3SxwLzMaZtTo9IreHwxU3BZSmptEnYX/xVQ0sUn
FuzO3Vj3y9SCclkIsi/Dmhc2XB6dndz081mqueebVQmbtrGYH/xNgd3hTZF/D9qHxjD4J1wEtb5U
Hta6runiCSqWSj/OwjWSi2OQXyxI/lD93d1/QGxRCYkZQAATieEO/2Z/6qC0eY0/RmgG76YJUygj
eg5lwrktKctn4OBTuAzlgw1agO54CqrCcP9sFvWhsga9nayv8D8omDcVILvcwW3G1fXoYU6/1xxv
zNB78r3uMkGEp0xtoMsuilqLcLced6lK9CTecvrJ0j06n1FzVKzpkXl+kuG0MPqpNaDatmbL1dYm
UDHjtdfKQnFUoGRuaiBq6ERWOvLEB2LX4SEnCgRksa0xv4arYcnM3bfo0XpQNv3rh2DhqMih9Um/
NspclzMIMuEBhs8XWusJ+capHZnqs1Daj/KnoHkTQ/DzgjFsodOL4UhNUP/RXYpqNQXPmD5iJkU5
/WTotghG38MZmjz7qcfZGvTR/T621WZE3i3/IEtlhZwfduGOsEYUgO0G4Ru3FpM8dAcqFtidP8BB
Ht16O80dY0MjTn8eRaBWW6XUGd0ST4cBpE20BjCSfDEDDnf/afv71rgSTncIkYULMX2BRR1O4TMR
JRRQunpv1grI3a8QZglEBCR1MOrWBkeX71P80cDFwagvYQbMqNa+DAhNqjI3lF1aYJP6Rt66WObj
lwAFkpwBBTmltJ8IxXdZBCoTsEvSnrAfSn8iSnnaWI0rNn4wt+1T9TSkqALnhGx9eW1+YEDP0oF4
6aFAlw2PtaJzpYifNtWlweuq2ImRo+XydxY4G44PEtmo5r8kkCwfeyNYLI0O2bkJY5wvjOHMUf4j
7i5DIt63TxbSVqZ/6daQtVucKpwRv5vsmQbYjIV6p/qqXiwWIRN+NhMEj9vYuzFgDZSEl1QoI9Q+
PkD0cOcK6AUh7D+ZjkDhGLUhpYVBCLM5bRdsP5irSU3mjlaVlZenZ1odjwwVRPxwqjNJwOf4CrGz
AArTitkY4ZC4/EEU+9Lm6WGIyacbhICvvROI5SPhqNacuC2c3HgBMKCAT1A4m5/xgrOsMrOzNlkG
8MI+3XUPuleCIzUWVSbLWbuRKqgTbDPV703Eq4/5NH7XrMm2Ooy9Uf+AcASPg/KqIaO8sEQGKY2J
d+KNg1Uow70Co6Yy6YmlhEtc5cOLvhY1RvUH5Sat1q78xDemjhvdVVsqA+IiiUgHE3gKPKLtVM/B
3JgNfHMpanEMgLMRkZuHz2MGSfIsErYsV3qZimwFtTMAJ7gsqV72Ur6BxVGqVgWiW7RUp0F2U/fP
dRRI2a53eDVwjT3UPAitmc6LJAT9XE5iPOjq7noySXaBVbxZtp+4y2N5jN0olTGc5Onohm/bYMxc
Z2GXDrdExOTFFJXwOC/71ih6VuoQwhUgFM0a+YuRxQcaJE0d3zP6qEzRDAaxNMeBMqJu2d8i7DWD
ELueSUfSMvrrgmNxhLhUzD0fzauYNVmrAlVTOqGGjnisBW44OTEZRDwlceAAiDYe7vt5fKZer2vE
rQKxRS4WRhdGG/Pvei3Ns3/teTIMYq1LIakdZukB92o/B6/sYQix//nC8d22zzV6uKVk235b5fvd
qNbHZjdbN3AOdBc3cv0/2wDAS6qUtoLqChkm3bi8obpqhpe1jRhGeHvZCpS9QlAeDxZ5E/jl9ylW
JYQxEQlctiYTI1Y6s/HUEaqDTrUYqB5bSb8q9qwLLjVrQKdAC2/3Kgslb+IGebYG5azpxk/9ex3N
LR3uEbTBR2c2f5rAgAZse4gV1q/1Ofa5f0Qks2e4vtcTdf0n0GHbrO9DutsAzo5r3TT9zuWP5eLN
P1Ri66sHu/l1Ge7cHaSH/fxP+I1DmkrPSFefGvFgRBBgQuIcEyh7U0TjJEzChcI1/rqlQBrZc7Wd
qbeV5CRVaek9PamwkmOkQpwbE+fGnlEwiIZKXqGoqsUBLc46UUfq1d/IneiBLtV3SmnLUPAqDEcE
Wb6+tgN8zBYhtKFZC7ednPN7N52j2SesHqpBC2sP6DY1AezyHExSct4X0XAomoTQz93+Zywffo1l
cRyGjgCDMnZvxZoHlg1dZyq/6YilY7T6Yn7o+tEuWhCdH+she99sbxWA83uc31aw8R7FnOuaqnvs
TBfSoAPudmA570N+xnfLHIy9V5br1kPPM0ZIUAfQWpdx1wTX7XdFWGVIpwhXuJEIqQZzZtWUYIkt
6KmCqXtCyEaoKvEC+iXUUWRMuC+NYCdQCfxm8B0KvAxPaaBSCRkRWu3AOqfKziyGpXTniN3FpeUL
dCmMlBLXvOhGu/7kh5Ug9jD+YzBf8nW4PWwIQrLZFCS01A1TyeIxLFR4oZ10PC43SiS9A0ntxs91
zuRW+h+b4IQO73EogegT3gWjxFb6RBTlcStig+bYvQYDCkQyzmOcS+ujFNCODQ+tudnyOgU69b9b
NwPT+gjjg52zvtmbFK/0t9CXI1FPVjbb7EqfJoaovGpFgQ1BMo8+eKX5B6QRlvre3xCKILs5Aa37
+hNBNkiUrQj7RNBIKLJcdXQAA44M1i6vSi09jD5mMerGuBet121/Xf6F1PQJzNo3XhHClr3O1P4Z
EHbDIyhzuJp0arWtjfqMuST9zun0isud625aM/UUE96G4WSM6CNNcFG06TgdXQplSiJPYI5rWsUH
cx0AEiDL/cxc9w1rsqui59h+vbDg4Ra7xVbNpOlYszPSGt5Jf9DabrHpVwn+p9HxZ5kFxMgPBJBA
aTQWH/pA24pAQOZaJgpg2E1hPzZd1ygB5JTeuFE+V625r6LM3MZTS2VTcIMEDyKWTxr7Hpy218yY
dahBAI4jakYKl4kcT7bnMX2DFAU0LuXG5AcCOX3/oH/awT8Rb6if9gKJDuxwg3K7e7PtKE6j+Png
6OAKvuOKjHWOc4qojFnf9AgMPmMYYl2thJtXrxqcG6vphmX0+4LEwmucfdpzEwUY2irKiPM756a7
ZAs1SB1JqiCx+Q+ZGfLy7Gu9/wun0uiwy6kC8ZyWCY1/XUoGBQ+eQ8T6S8FEJlF7Lk8yM/OOLibl
Ikgi18Nx6TSKkqqSDdw70Pv3BP3fN+RCh1o1zkPfrivYzKC+osHedh+dHgTU1RAhxaQMrhSXT+zi
c+GJfC2kV8lDZ2enw1sf6qybGfd6LXsrHbrAwbjh9cEh/E2cNaMJ7+uylhatu5n7S8hXclrwup6v
LjkM2FF+bJR60yC6slskVejeGdpLfEQtWPZFVWYpIihWrlfWmVgIBXjbMUCGcLWScDq2GmgmicI4
N3feg7uQBA00kDdbIbA76NzOIeuJ2i3Dd0YzATs282P/DaIOO0tRfKzo90YaN4nmmn+Emj+kfg7x
zyV4vmxKbcV31YJ4WKlHYnu123NNypRwj1Ea9autqBL2JYFqEYV+B26+bepKAYhwo5XD0txAy0oV
RsY3owavO8m5EJiQX3L8SuF0/NG7RfwllNjWzUdAzWUgNgGK9JfzMz4l6eZdA0lQBh4ljxhA9/7S
syArKqK3YQm8aZEpqriNZ0smCPChSRFpqDFdvNcO5kyFhjtY/rCtvjlhuBZ/WT5H4EEPxmCxZfex
KkVS0CmjWHKM6VkvmKdXqHqKesVWVuT1EjGNGKqRoXPKGHl1DYesVMhga/mUsloA1f93L0MGthnJ
mPlS9x1VuW+urbvsE6vK/ioTegPSewMx+PhYfvSdJ0ez7UdQcqSGv0Nvl2r1m1iitpcaNfHqGVhP
KwGt5vy+kh/yZ2vp8XPSQwVWCNNyofjnw30QIrwoQ52OF4JThr9snR5RfPiHEjA5lm17FQy6ts+X
//cmwVvXHAZ9HWf6G2Lvmyw5idvKMAGrSKPwio4pWoQ+rfc8L90Nl84fCi2UplfjT2oT4F6rHHVh
NhV/aB0d306XmZC3l6A3KTgVrRR/CxicioJRDNodsNUPYAdQ/rdZ3SHYLgVhKvlT9cdBQjUpzQhQ
9t9PLNlO1tVpB5r1G+BldkkO9eg/h2VPlP7KPM7irKpm12NTebVAZ5jbcANXN9wbxxnVz2Xmemmy
NOTkSseJ9uawgPKCYwaBrTCDwFiAjyOuGulUVplc+rt0keuy3QY7GQbLfOkgxcbqyA3DgeYwtbi5
W7LOAVqsScT/T6ZDPNx+ZdFqdGgC4jP6uiZS4wRef/C0xJKFzM5FtRrWnWWXWTetiAo+YyS4RaV8
87h7MeD14vC/LbW6tMFC7FV+mcNDtYnO1egTyQ0YJyE8Qlk8mKMJyg6tTHpajljDuc9tq0v/NFhZ
PTUkbIiwv33r36DZbS4sFxb5Sl/btcAPGbuzW+DhplgqyXb8UU5JFZBikjypJsHehFQzzreqbiP4
DAzcZEMwbH5OH0SONq7Y9DmmRHefmWuEOagyJQqDpszFykMn0TycshMg8/8VtFoStawR3OMda1uf
0LP08ty3GxEkfIcXy1HLrzPLkDQ24nFTNA2sWTGurHNsI+yVlvD6AQMhWYDy9KLSk7hP4DRsuYh0
BK8GzhB70iugpCGxqngywmnSjgHVDvhE/WshRRs4rbFm2HJUoW6jTj2IfKqSk6ai8tjxwwIz5Zjo
H4C/vUjvojSTB05w65KIYOwubebqKCg8h+u6kDFs/WlI3YB9FKzQefOwjN1DMnChEQDP2FLoQ02x
X8pOQpT2YdC18uhhEPYMlexmk2yt9pOkiXTc0Z+XAmW6ufccP3sxuzGuCkDusGU8hC/adPulYxpl
V0gr1LEKFhgUniEZ1EtKxh0T8rKetZbW/cnbczEMGklesCzxmEMgihN8t3jGNMbLfWqszEegrzkp
esxfx2nnhJDpRakkQnbcoz5Dof7PR9bl5NjJL/MyjEnnum1VunK2UpJLRO03PqqxBDh5OYtSLCfn
aOr7dQxz6qSpPzyPL7DeHT4gLwCqazxVh0uIRUWzp46ezvQHrA76hJTK48D6JQxTGMpyDRBF+dJ4
5AyblD+WR6PBNaXi6U3g+DgSvi7pbfdcSil7MwXneK2/PbYHksWDZhYeKR2QR1j6bb3ITE4zQvUA
yWjTl38iB9oVZ4Qtx/ZxuSx39FhOCpGHOHCHuIZVHHN4hKVTQIyfvb7JCD4er4HfbJgUAR1rjMkh
Oofc3L6xF0oOe3Z7yayGHZ6OTMlCROroRB76mcUj4JpmSPTUD5KkifYmyPH4uTCiWyXH+nwuMXSx
vp4TbqC5etNSt2SHaMWiy3cT7a/j8dB9pPvGJp+0j6CRhnxub733NW7rn2w3EeyRgjE4Bxz6cc+2
+vNjkJbIA7V/doTjgpXsO7eJRtjzLnKAbdgHHSWgJSugdAucTAs+UeVbGBU3QXuebE9FEdDFOlZb
hKlDNONbHT1GQdvOtVAvQdtvc5Z/joyJkNacztP87gpMwaEXWEOZLf0Sczk5pX0dWL9Ok5Ys3WyW
o7DC8KLfr8TsjSaGsDjQQQNlcFpP9uZxTmAj7AyVwAgiSTlmQyhDfyKp/4zQmSnTUfnmFwqD6UDD
+jlSL8/VPrhSF3JA9clhPNzL0nGrVGppRoK8wncEoyFfoSLowFj9scVEnB+lR9rMV8hw4UFe/WGU
l0GIMeY3bSSHLy1h1vqgeGxNRjbQKmArYXGh5ZbYVjv4I9r+rYohvPPLFrDrr6EvjkbMjaGTpwaB
Qo+SxxRs+6EXjuangUlQFzVOg58vzUwJhEFXQ4QBKdUyTHYp4lMxvK2ESkICcs1ylsRtPbB+g+kf
t4EPxGBL2RPBcFjXDhWNh3fXEyfstLH86zwi0YuMVhuZrVCK3HNd46rR+5ce1BVXL0WHz5Zd9OUH
8GMtwO3G7ZIl6n4sUFE3QQMCuMGPEcSBDqgjpVQDi7uncObKw12KgZA+U0Y1TIclyOxP29JJr0Tz
ku7+2/hbfoSYLuhl8QoAsQ+0C+D90MwLkRdNeZD8kIKADA7j6QWfMAgQpxr+aRpH5SOXKMOLcpXd
VWhxEURaLBRjlAUQm5vY/c004M2iqKzUhw9TBPQfgnLUfgZGMSSzTsR0GYsVekBd4Xa34IpZG+ve
rz7rdDlIxCDKfidFnNHjSw6CjvCdUvAvU6Mxh9MDR5yuDyI/B6oTAmLAwvSfmjCUso2CboeTfoqY
vzXm6kqIl+p4xjL6yWRmYBy51jNZPKjWNutonwGhj7+prZs2XgnTZ8GCcruPfZeHhqTNvwQ96FHA
zDPDnyod9k77lUiadbzXCXMihHNQpE2zeEMGabDbLKgqaBUcV1tKxEsgkXt6aaTI8mTSfUEVsrOu
0bAWAun+kE+HzAtKkf66IDyPGd/yJ07gcecCLKdKNVKUrBWK7huApL+ALdkVG+srvlFHXLH2xonB
pJLdKz/LlSYqLA+QsRCf/kWbyOUlvYsT7RHZsNf2eqdPhPpDFdf5tHL5WhfQmBO4GcIBtmYjCvYW
6uvSXaH7n9vjxlDUdOmrQZEO6JOCGvEIwttdBw6XNKjrU78kTrmX3aE1gAztkGEeZL6DY9P23aKQ
MnMcbR8dlxi0yKb5pOUuo8U/OTCXOag+vkIp/J8J9F0G4eAXdTmu2sVu8r5gA23bdd96/z42TJN2
e21iVKhoM44KsJEsuD8bqX8yeQzwTUPsBBnzX63NVUl9wTBXsVEfA7xTTM0586ejj6DnbWzjKCj3
xkJqs0xBXsjlG1mS061so0CGZNi+U1lWCOrGnGBaAUquHQexr0EUSh4KmdUQ8NmJbSPAq/ECQCGV
j4Ut2Ourjy71kPdkaEmhPTQ/iy/1srWmtF3e40XpJRt1x/rfd3giVpNdXPI59soY62t2Y4iL0KMS
pkxedyH6hhMSTpGCEAF8BNfICDenO3CWyVJVIw3hxOHJlCO4KveZzJpWHmADvOPgIjr+HlKdGnpn
WfyFdz4rNLabwaYwSQd7zVMX/KwJY4RSF0L+ROB2xU++Ash8s6FZAtyATe2GscSQIzxDht5ltkYm
0YEw1+bYEI6aR26Yl3d5XG2pW3ay1dGqctiGl4EKLZTe88gixUjmj9UUtw2rvcxwsqWUJxMGxxL9
p6WdHQJbFWjkVXm70uHppcrn4AgQBcpEGhQPJO4YRLooQoeKHWQ4Lmb0RIwCFcscNPl1ShJY4Dju
4VdXiky6+St3fhl50FPvWNluXn6v5ozFnpd3y4AG1qrKHkLvxG4xOmKM8QKXbYveladri8HA6UDI
V0lqI1SBG8fZmss34UsTw0Ui487I/A4lPkvHbsiaT/wtd83bGpnW10YuQ4WMAB3pLPp7MlpgPOqU
drJKLWz2BNRmbI5TOUQwhUDU+NpIgsw4/tsGZAXPNJGaeijoDs6PwXl/b5kHUSgDUAjfXSR3IWqd
LL8JIdtHuxEUS30smNsb+73GnAkGUBWRefShbFbJ14tcerbLlTYxfU/4a5Wda6jOXDXbZ7wJ3j6g
jJlNW9PPEtTkzqPrXhtspzq6WkaZMX+Z1igBqZpXabwnGVYCjTVyeDedySlKguLVCU8YHn7v0ZEc
FxrwAZFFHD2Xzlvm0nvodT6pwBPjH954A+k0+5c85GLXJlAAKc1bJo+GB9z3KFrQTu3Q3v8pGbrV
BERLdOIho9cTqxhpU1bGA2NJli35gR/HCiBtMJ7PtlOAHrQYdRD+qrJaMDcAHD9dlZIBSh5THgrC
mQJp2kz04VNWBQJGNepdb1cv20uAwMw29rTSBwVGyJjaKV4BzW32Kt/uOLRCbuo6dPUH6Voe3+n9
gFqv//sx0kghfXRYkmWwNLrKqRCP6786KYaRtI9J8nEuU00Ej6OLuPxaxFy8B0XyOeVQimZWLJwF
QYR9MS5hBSbjq6s5zWJWQqW9TPTQn1Rfl/UhONltLNoZZSOG8iVTw9gVXrRrqfd2/xG316WckoCz
5rjgMSx8Wqe8iiqgIEQCgazzf8l16VUbsDnWkfeJr2UvG7mN3OIS/tgUGjNKJHZHUQ5KDlvVcMFA
pWVxbh/vRPHEqHfEP4X9HwgI8MXkC/xoHP7cqtFooIdpGT/24kMTjvT7Ks2EPB0OJLdCWVRdyKz/
oVS9A/ND8v7z5fXzfgGf+lAtylqpA8+o41yV8ztq71ecXFQdnZv2ZTxscKIbM2w0CQQLOCpknnxG
cQS+vNddeGk2ZdzO7Jfo3bbygmPc9d/ABx9ZjVCfiFHSot326ZkSwDQE329mWBnjFsacw09vNsfy
REYCFYWS0ZvByIAqtRGIZzS23n1APmSnXduKrVg9sehMI/QCgp4GjRJPuOfWcY1zqgnUOkN4+EBx
OPTXBfsa/iee3fEHH+gF+HPS1yVqCX9YP/qlfbtrelRE+ZD3kdVq+KGFlHj51z3JGwR8rd1bfujO
nBZd7Gd6/6YfnzcJn8/6M7skEVEAxwKZWD08rowSxeyn8fhF7mTI4TLmdnNfnOIQ+/6c9MWmTiQG
giYyNNcooWi9g6v/lemIXuTeAgrDKK4QVSEuL4dKqsopkuOY1T92JlCNmHJXysUSYtd8DsJ+V1Yq
+TsO4bzvIgAs2Rvbgyv3NTEbG75d2sm+A/uHqb8yuN1i+Ocru6wAmKcST95vHzYvG/PJNFwesqSs
HR11gfsnbUoYBdoxjFnTRhij7csrm0jLCmQeI6qlo5qUNollWJlQ7Qs50z91GzfRGfnw+u7x7zQs
zr8mNVsiyLWr6jBSTzI0OKqyuoevHjbPqPMDwH7FkGpZEXdeu8h9+EqlzlMh7frR6et51Z9vvfaM
a54iJAid57XzDk4wn1CKkbu5O/Wl3KsAdmFqmWAY0yQV2FyR/z8CsCb8ufnocW6Rm1SdpVd+BuUN
AikG50spVSWXKfAbZeRrPrMiOQAZp72fanSk+Q3FvZT1w7DI5aS70Qj/rq2pLIfDBMysPOB6wcKw
hta6UAYsvwLcQ+yKsRAY6naS84V8KB5dgnXudUcfC62Gi54VhW6MDa7HS3GUg6+CSqTKLqhM81a7
15NQKWfycUYMgjpUaG31WJGXth6kzOBypAQ4XfT8BMLrmHj2kxij9R2koXvPwKp3ZbJ2SsPwboWG
N9Nv46GopkvPA0wYQlkuAH6Xy0H+sKCVJy8SkLDStDxZdSKCrCskJdv7OpLMrIJNyDBcbLJE67mi
MyZzgAoiMPF/KJUkDEB6tZi+tv3Ma7Q1hAobrvqEJj755/a1ifmwDiJhUITKFnZ7v1BjitfiHVqq
7fDIBVZFYhCuIaScK8W6eN9CnnHGFW4KtVIrx/8ghoiIxVV5N/V+iQ+AzHrlhLLeMJ89HVq+lTwG
HGsIAu/uURgPEiJ67TDNwK0wsvt6iE2uSaKEzey4OL3sGNb2FtmsPX8RjsXhD60tXztDAV+5jovV
WRLLX9n2u02WR/ODZQsJ10U9n26T/aTkJbfdIXSVs4o3aUnUJlKYZpbMSL6T1Enjj1HNZhUDWGAg
jfYgR53GPLj3vFLmCBngldq6bIE5L68yTWlEXQwN3ArY58HS6/ZuXturzm5uT8eMwAF7UJjBqgMB
WcRyWobhTtuEbLqIfBHsYZo3k4Q4HNlneFXe1xsdBzmPChsgW40A7XjgFPsukYp+uM18umLuJmIA
7EysJ0JltcdoeJs8lFzu1Y6iwIHPLmJ4GdlrnE/wfb2yjZXc+UibsAenN5aPSgekh5EYiFEfBnTM
8ZOpEx1GVLtObADkrmiQGGsm0HxlWH53Yp4KqJFZUeZgy7vY3RuVcRr7vLAviVu1KZuPE9RLjLcQ
fIhEnXzGIDsxJ/1QsSc4+MxVym0EhHKGHl0XyrsuJKpgCXAWi1Llu3ctWNzNMhLvoklA/aQ3742N
CTa0jgxpgHQz7C1cJUaOK9AsUVDp46f9CDOQC4hiUeV26m28v9bAkGvwnPU8CTQ2CZ4Yfeg/vVFO
xIR1JbkFSEmpk5htm2YLc6nn9eBiB/v2jJbu+OD12IbC9elW5Zhyzecvt4MB/jmBqT/zPUW02H1T
1kyNA+H/ihE1tq1iks8qzDNZr6cxh5n/hDrzp73R0zecyLkRFRvd37HvXgahqQasZ0h7l6t4S3mx
Qkc/RnvTw+ldH2FcPKi8WENhxoMhLxgHXkkARfXXZTG62K1Dr/PcztJTwzYdK1ZgCQfc6qVeOVjt
yeXZ83s18j0h+TzOBY5rjQFQ2ANsf1dilTqDwtcn/JP6iW51iOXkmfuFNdk6s01pPY0k3iDYrvp8
53ZtFSsoNNc1koF28e1IG7eP81JK8tJvY+Ruv5mcBHbLhAY0ssxw1A8fQ58cEE9bHvFt2pGiHBND
w/JqSp5k3SWLezDYNVIiTiVvivJAxbJdrPafZjEmTT+E568CZInHLRy7Nwc/dQDyXjUYA5bBAeli
h01VGSaAajEgW4W2DIDiQU4jJxLUkU0UnaYerAd2wylcJFj4yWDort4OQc/whagAVScsilsaePZv
IpEVu4EaoaYUDdzoB44ZvpBK+74iPSzx7BWuK6T5DVm6+UwiP54R+9avb8CgmPGACGKZDpwO5zrB
h3h+31YZ4NMTQqFUpqiqHcQtr+Wu0bgfdkteeZQMViRq5POuYQ0zfeE0vS0JfBZ46l1zRRmEwmgo
3Y16vxV4pkW5MJaGnFdtTgQ9Zgdb6X3DRQdWAsirqUyRMTVC/Tf+JsN007Do0K+v/A+LVeiwdI3W
keXG+zodxO7dNNm60EK2v5fIK/XqH45tuzt5Bka5AnDuq8oqnfLv6/P/wcp+aZJLbS93Db5MuqdK
dlTMe8iVJtdgOOcaXLkO9/s4/yd+0VsbIrIRIqjm1UNupqe1gHbCxWXyy19syyeSyGTQSXwIpOkW
MEhfZkJItMsdG7o9XBREYgBclKL3/lpUIUPgpkCKQ+hTxihX7oX05yD9RZ5E3opaOrTFGr2mwSQc
fqRA58UichfSLqLW1IEnWf8lrPBbc8gMNERZy7z0JQltETxp0pwqr3k8UscnIG6YVkGzRa6GfkJO
muRy+bfuQ85SaFbzHjkfBpidl2tg3hRf9EYuzmAp/NCFLXKurD11m7lO3EiC8vmhA+Q+a9k3hc08
fd4+1cscXGX18bjyVF28yCW26BsvV5d8HLKtQDO3m7h35zaniH1nZo4FfYpiSbzjkxfazDFDTw2c
d7s5RNZWLCTobS5bVxnY8tefh3Y8j8bxfPLwkmGEMfxYYHv0CWHtV4Tr83RKb1Pj/UBf10VXkJg2
0b/NXgqgupWiQQyvMxq1CWchR3NLYeD4rN6LGNluZgehE6g5TiBy2RGiN9glZnYEHI/oE2E4b4qJ
o0Lh33mLZ7Dnuz8u4fHrkQ+JYZxN40AswVzMu1UyaUTHGjp55cHYhb1KRteVLZfwAzkEjukgR4wb
prR+FG+qShr5nE7hxbzclcUWkujftXxwv7cfzwWc261dyczvbrZbL221LwXmEGRokEorLjnWxL2f
69KfFdZnXG6uEdCIN52AGC6lIDGZAcE3vrZy39bknzPI5l5ZKCTWac+Kd4G3kGndAhyR16xOvFL6
ihzJtjcMSLg7YyCumWEKuNFQpl3UGGH/I57tBabgHPNpmm0RywH72igJkhr9Jh7EPRqxgBdmx1L+
pcq8CJbXiaxjtyQX6cajWxX4UoooPz/VZuNsHyKmzlyxxSmWr8DhQhpFtTFj+27Cduu8qwWjj97D
IKqH6mUaYckymZ977px1CL6J/OQpX8AaDkonATa8yc/x1WmMni0n2DPK3UWnm3laM4o2qbmEq36Q
KCYDzaqp45QhEeG1s8mxkisrHnnaF3oQCuCf7a5J3ynxYzR2yuG6BDRTr+iACWaRZYSxqzkHF5LV
NteqY/LN6XlWQrZ8FhV0bkSNLnoU/PyAH0Dlg2xDHcTIMdp+wGQ7SIXUj1HCecpVkB7vqgx/2ntZ
8kpxGlRPRQJtHIyrzsjP8TEIsA1ENyrYjreJ4NRF5gKhpEQ8EANNOxgVWQH1mVkZced3kxxK9fnI
D2pWXPa9zlLatdcxBcHjHeJ6eWjB6TuvOyQj6eLXxylzXe1Ej8kDsdAxqZCPoG82CSXYMImfGLju
qPHH5rD7ykg56czYPFPWAiaM71tG/35HVplpGahpmiwc7SwmtEVg/VcC+HXYVclq9Ld2oI5B33d6
tQEG7BgFUo4q3fkMAHKUC9chROXbLKqij/Fy86QyTpi/qJdsi8v3RIRtcgF6X9V2NpFX4CwjiKpr
fdZPI99lBeuy9TTgFu9nGhW7EBrd/4Pqq1NmuHYmQqGbZ7Ib+WXE95hN7ALUTsA15x0hGft76z+6
odD6aOa0mHxuO3SJUkSmzBkHXzmGF4tnK/xMKgyJUedI6I0vdC+y5eVj434r+Cetr/sDG+Xm5MMi
gWrf/NHdFF7eWJ5MWbwFBlbovnpfuBjktsz5XOxiMmuIF/5VAZ5Rdhxhq5wqQ2hvnfnV2Z+uWhS7
okWAUyRUIS3FnEV3bf4L2EjBOie5u8jawUwpzAVM3fGeTRMx+AvaEQV8T4FUjf9z0s5faQ1COyyn
cQYcX8SoTqUGJCop/bpDGzdRv5CJP5ozM/B0sUpGMJBdBmRXio2K/78dU1VAH5RyladlhFJMIClq
W6J/FgT4qSYwD+duTPYTXrrVhOigoMRMtOgpyF9qQgYmpTob7ygi8shvYhj+S2OP70Z56WxChyBJ
gVPmBrW2GFqJH8hzPJc4AnX3S8nvoYycxE4dKSWOuU0bnX29eyNMyW8sGNoBx5dx1iAME2IZnrJj
3A8nNVSd0NjOztqgkppAekmXHv9lvH3bH2pePXIGXEFf58sDXcR9dvU0/r8Ue/+Zs3m2Jwqvlpc1
qBzamGO8jA3YxN5QqEfkmNLLy0S4wnuXHFMb0PM9//RMBffhEesk6FnZbb9P5qPsFBCZU9dd7cRh
ZoF6dn7MnZ6Jv1xEBKk2CPE18OcvnyI5x4QrZFe6fB9W7lJ1AfqQz7zCO50=
`pragma protect end_protected

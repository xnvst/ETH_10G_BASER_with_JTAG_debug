// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
TIPtY9Ockg1ApXarkixPR3wOeLarYdzGxTro8nYPNyE1GdSjhOGjwALCAaWus38WIw6RDAikH/Rj
hI7nzc9gSZnXQiilAtRT7sQRCNxjGjta/3jxAXAsIRdMfeCg9kuWKrQsijWHc045OIlNbl8AoNlQ
G2sQmaB+tdecACjwi3qa4U41HZZ4mfItJJCxSaOEY2ci0pFw4lfNZMRTsP9HZQ/dNFv0ptQea2iF
WSaZtFAJ4NnkIP/SPXi/yp2+Td5MjEM0yJFaXyJrJ1q2QvVtiIUR+cCBUfK/1q8mSd3uwRNRS0dU
LSaWrWwLzu1ppxPu2Jn2LPH6MWSwnpl5o93ywQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
nIpK0vT+cjl5ttzOj/bFU8X/2oKbVO8PlD02n0DFrT2rrYJ7eXaTldO6a2J51DrHRksFiRxiVHi1
hOLuuTBUmcT2V/JeRgfLPDgfAC3niZRfYi+8+3v1agEPsPyk3ZV0YlgqYPIDurmBJ1lrU9BrhWJK
RlIvsSPrZQs+CKf1weU3peOsy0S8YCBt82XxAM63mau7xUhBqdNr/jr+q/4QAj0iE+JjQeCoaDGW
pZGQ2PgeYpKrxd7dDUHyXECZd0SjCff+CK3hFfP/GIRx+D7Gage0M33Dr4xnTUfx5App/SwiJ6oP
PCcPWtFRRiudUsoU0XlrtTMVv35mfe8Fm43AF76Jeal21QvBvYIqaEatY8MBxWHV1TMZ4D3cJ/BQ
94iXj5+hZnAaGIiZjyhPdxYybaaBkPuxIFs4+5gO8+atSaD0aorPd7CY3SRDHJBfpWE6VUsnrllE
Hx99KNcGRcHu4/iHrbMnv8a8rJ7VFCYeO5N10AYu3NgH1bRL4/2tWhAef9iXW9fFaVtHzsTIb60B
1MaiKG56oeRkELC6h8/JmtVwYnKqKQ6oTt0BFs3KWov4XJspt6YsKDuXdaVyaF5zquTdLljksTxT
3lbg7SU02MNlQZqqkjDF8j7eBjsIBTs/BvF4H2UKhEZYX8TWRzLE2u0XoF4TeUpLCu8Tt5R6zhgp
u+tyPne5q707nGXYfABcPk8Kkkk1COO3hA15ZVjzR2pE3ZOT67tz4rc/ro6Ysao63Drvd7oEAD/4
lfGimI7Uz4ZoHQoMyGhfzOBkhXq6/e6YgqpDUt7xv7dFgBGI8fCH6Opgiy2v1Og80c8Fe0SN35um
aomAP5NRsFRjfWCdjhauqcmLF2Dl0C8f353KDRWBp/hOQaz9cyh+LIEBkMyOk+ek48WD1/TfZlcM
pWi+EC9X4wixi6ffveGiuQDdoAuK9qQhQd97zhhgBV5KUV0CvpU9lLd0E4D1lq7VG8mzZ+vTkoUJ
wfm3qKte53rjvtx/3rSuYfoU53ZreXPimCeFOWKyJM2XKk7UyRjNwdlJzD4APNLyTQ1Nf/ZjKSHI
3R38qf8T9pDhQSl3m7xNJJpoa5avVRA9aA9vCKHODI/bmogBHFSa1AJhHCMj6Nsq10VF6sGjDlcJ
wczfPU+c42sUN5fXivO6j+/5KRDwgXePyVzht6rx5BrQvIQqXVJCjtVvC3fIJNWpQI+VyKfBvRJf
2GqXlnry12MrW1n9Pb2Mb/yQja1+8DW6z1TsPjd0ZyzM7xmz/5ttR6CruWYx75QgOPCgAbXyFpgg
3KJHCks4AIV+4E3+gL+PJNqmpNOifAht6jF/ZF8cTf+hH9NJd9qa/vBCuXaQO6C4+yi3l+ZdBTMN
6Cb65bvHf7Xe8a9gqrnDb3oMIAsXh6Of6B70BsNIHatH9FBKI5WWGSD+jobELeWihvjMPKQvJ49B
OWTX9w5jWf8wp93hRVx396QSVdV1nHgOnerIME08LOu2xw06dtty6yKyL2K2m9piPg2gPB6d3fq4
j//d7Z0I/qA/HpSL7XF7dO7Q3jsEAS/QZ/F9XtKwWuU8PIo+XfN53HfZuGU/0F9Hn1c15x7+z3n5
qP7jWbadGDD7yEwt7mslm2wwKZETojs3rqiL1Y/TD93EPBEXhw2FoqjKQjx2mfZCdvtIQDtxcCWm
vHyTMtPhBO6noNYlyHyLRA5sCt5aq+bkpIlD65JODG08xbR77fkFH3SiAnNVRDH4SxzTqxftYiyt
sED1YfRYg4g3YQGXQrP+feDJofrB3vkVddaSlDa3eV8vkPTiHe7ihKFvqnIqoHefyYtXmKQlfIZK
eOWM4uzvxr5mM/PL7IGYIFP2ITRkdPemYH0vPgEaLkGHX10NTT3depAhubDjTeJ6v8S+5uPzzJwv
OlHTR4+f+SMSkkII7onC21gDZh6QDtp21ycu81tuXeckzNHVggMxdBBpFjZq0UtPtndPUjKZfWao
DXw5PtzE58LyUmDBV94UyrbR2TIkz2gtKgszB6V6dqSEaZqW5RMiYFGe6QBGPyxk5PVdxy6txwlI
TVlcHRFAo7CXaWwLi36SL7DVRgaZAaxkCk7etrGqNTRgelAfz0xZLnpG10sfDZHPMwVp7y3FNj9x
AwYuNPNx2H0cA6C1PLa2Kt5HQGbPRVXOIjzLqvF3j8Z3lhmKCjAwg8L0wlQUuX/itD7AvEvGHXxi
7xearX56oPwEuBIJHhvVTqm5G1G6VGWyVShJqlf9HYUNNxRmAuRhRUDWarXmBdYhDMJiCB92icc3
flTy/ymyX0RqVV8Wbau1D79QM3ha1p4RvgFP2UVNg8j/c6tmpL8iIA8Gy3HVN4LHYeXaTmPoeNZ9
K7nFL9MO74Pw6Ynm4Ni903vD/XdsTkr8hcMo7vzAEkEJfEJB4UAEW8aT2W872PmzxmAa5/8abZ4F
G2LMsCVQIRIrmqsdQijdvi/9fBazDbW69IEsDY6JhvZsHgzMGRXhmpdmXApQF+nT7XD5k6z9a31V
zMQ4wtos4RO2HW/LLahQUcRCBEeGxxHsK/GaXD5d5UG+iY72ZfMP3Gvf+7pddulI7H7/wIqVD6h6
udSjsFcfhU9XmahvpDskBotJEBvgMPyakr5Nod4WhOITBjDiuRu4Ww2LAAjKtRExPPCD9lJ0wpp1
66aTIm9zP5sZnruEYxgHKruvX9pqTAR+uaAfoajGZcV2hQorhKdgTQRdJfZPF5RDKyhjMZj3AM9I
TqNy6ZNDyEy/OBTvPWh5dnePUSxHNdei66Ux8Zw6T6yOaT4hfwziC0g9lsJqxxg1uMs6BdWZBoD3
7pRJWhTGwx8pHNhC+1RAMER51YOtYMoCNKI0W3lP/XAQ7mtqP+BCqUAn3rRU4ocwuhqvSLaX9N2A
zVlb7vvVhJrwF83bTw+S58Nn978SihbUabOtYeHSgPp+fXQalil3uuA5HWad+h5QrdNQVWyeYqWO
x7F6A6MVTlffa0FTqnHliVaJeBfOhTvNTxHjz92vTs4npPpd50KQ8uZ7/PPOZhgs4IwOH1MCp9sL
DtQyETMvcB8+oiXVlnuIl3xOWTpigTppNLdl5923ULYb6BA/+mPfjtU7dwReRQ17GSmqJtJdmDpq
Oz64a14Nv0gfaHbt+JRBoXU7N5qs1kj1dT476I607B6zuLqGk0lPEv/Sfnn/wFEcTjihk4DMSwFG
pgYmesoj6hLTVOqzFLDBaPgftG6poaQkGtj4mjkvoprmVZf3VgyJCvvAstNZDIV00vVUg9kPYGVG
1VChxHwEaXuORub51DXoNx1pQDDQsANcud2w/weeeaouzcoLB9gb9heFkzpk7M+tjbwYxcq++r/q
dj1+M5YGL9hoV8xZR5TwX/EFryV7Q+YNy4VtpWgWxhbOSHfZbzVmpn3wT4IeewEnkkZtPlp6Nwbq
lPjIldhXuVqez85bLoLWk6RzdLMOdv7LmB08eogQVJvEdOCINlQ+OygzN6ZIeBiv3m1VIHHbsf8J
TLf1UerGeMkp4tcSckc8SmA6Fm5lK4ymJp/guR6WROl7djHTFQPB59sEAzAxSEncgEPg5PWQ7+bx
xMdRbBwNLQraJhjK857N3caHkj/OlKdWwY3D9XpmoJgTS4Tpi0naHqDO4SwrKhqnWQI1IAoOdLAS
FHjLxoHEGPBwgddPNWXs+aaqv3ech7iwbn1peQsL57lUp0hb1q9ghVeYRqRr9+bJ1azX075Jnx4c
eytgn+gmgY8uthm4UD4hujbe+c1s2QBusOUFBDo4uuGlh1jayb25i4siYdJVpEhO3vjBM21fCpMf
N79rX9xJZPLMhaBgFazA6Axcj0SD3izNtduHzETK//VbUpyBCS1KD7MYWWXhcUSRrpygtjvxX1J4
rGcr66BiMNVgQlsUJwjFWCXlc4AwwvYLvZ5T764hrhsYb5kOh9NHcJouoSq0KnTCcuQTvhgsu8nk
QX3Nb8lpCaTupBbzzGN08iIfrCsPsH4W2h6kihMtboQOlCabTawmxMY7CmrMp0ncCdDLnLv5SFTy
P/NKztJVFwovXPYKbkjeBt0pAlX/iPbwtazGLXsqhPDVVHXVkcfZGRyYcJ/hRgteo1dbZWAQcycM
1jwCuLcnRUoLLJf6u8UEayc/p3cawtGGmMth03poIdVuP2qGUqIssSX6MGjEDvpbWcA0Xwr3SC+E
X07HWwwx5TqxQqZsVeyTZ9kHHBlAvst1hE9SnsdYrFLGNhKkQjpPqQ9BLE95wDgY/Kkwy3O41kLO
F1T3/DuZiIr4xUEzzAv29Pb55wijuhl/KA9xfuK3PslExwtMKSmIF+wHQ33rZNkHoNxX6YAPSV+t
29XMjePCIy4EayqH0yO7QbQTCgGIAaQ33iM6NWwn6vItzJyhPvw7GjYUK35rurKgqbd7QnXo2piO
cOEjBebZgVI7FpY4CfagP80a+MkN5UrRJ49gM9eOxD4pEWSaTROAlGUJm978J8MNT+7riqSCdG0u
e6dJUSSYda5VX+OrwUGlnxfdA7rd/WZOUnDdXKHukJphCORNOczSSwvdC/An4omuNs3Dx8Y0DTPc
sqwddTrpydz/CJghwzmwW6DEElbWEyeeum2GQihJCy7q5ruZIBL+3PJNf0nlt0IMINXAHrb3GOnB
xhguKu2zi2Wleo8rDE7xylUC/vCxJ5EnsQa0h+2c4RnyLgcIBZUbHKyI/lmm40Yo/WlHO6iL/t0I
abYPArFdtfoOJkH75nnkwxYFebU905YF4RO/91BPnqLW6EzqdvND2crJqh7iPuvHqhAA4uaLPWLz
YiyQrwy8Q+txu/NqN66Zu+nRyt2merG1UU/1JL+zcbfgTS2Z7oGF3Y4ETFKA/onu9LB2ajWJ1Nte
2lglBkO+jozAQgC3JLmRpvmh6qiz9/8MUuvp+3NK+ueHmaO/rmLYGaigNRDISVF59L8keV7TRnNX
HEAZR5T44CeOHok6qjjHcb98y45apzogm2G4ObHdJ+IVh1UZkiDcVVcR7dw4zXtMvQnT/uPkNv/G
ZKO8xMTgyB3+g8Kbq6AGxq9R3Izn3y0DVrYDCDkxipORtXLBs7RWskVz+jWKQcVDww/RbZyv1qma
1X8jKzpkH1LAkWhyj++MK8DrekbOZxVbT4MBJq0DnAp/dXapoD0P9WWybV2zPjAV8srl8tEhVL0t
EtTzrNTf4gS4qTEsLdGZ767k6gqHYg3+J3oDV3Vb5gUMhgzqC+H90ZYHwwcnrYBX11ClBpJ2krHu
bDzvvHZRnCFF90KLMOYm9wuUvfC1XgKANhuxcZdQJ3FgH/DdbiTkKMTNDjl1Q3yXnE95zMUNgvn+
p0LiI7YFaU7ofM43HZatLDDPioHMXefbMXiwGsLtYFDwFBegiIQpQJJKaoQevmQaMisxaIJdF+/q
J3ZF0AHrkiu5C10jTtcxQESKc6Ik2PCG+uxM190HVc+6X2ier/5WL1BqqHoqtAewYWPsRFS+eHrB
vR/h0owWmWxFUEBRl2MLDXgezSoNWz0BSDjptlQsjKkzI/2K/kzmoKY0FJ01en/tZ5xowh5oSunR
496nDPMTPYFXEBLC/ZJUgkdTFORHR2KFP4Nj0nZReEKSOkInBS1pzF39tA/47wKyXXus9cE9Nwaz
9JVFfysn4blow8ZvLtjka0FY6FX3noeI43c6FHOhZa/zq1p4Om2ByT5C8kG1GLQKBV0xzvM3YZe0
1E0WKI7fyv/Usg04RPTaQjGJFNF33Kb+sOhFOMv+MTjnbCMspM4MgWVhCHutEPMaW3ngv5dbfDpT
hZOxvO/DC9lIOVInoEPPe6/7CqXXKpd9MuE9gS8zIgn2tdVjDysNsQVYGkTPpZ1ATht8G4Tct+Fj
qD6O3EAXUmfSWNWIVspjzvdyyX4IIPJmjeX/ojA9clwLDWX5JUuIcSiaFg8h6OR7UnVqXDqkJELj
7h+oTSH3vks2t/2FHzJK+4l0wtSMesQCw3DUgjxCvNp42i+hybf+oLCclpeET1ymnRezNdXThF7W
k7ykzQq8Voj50udITK7vpRgB8lzD3EkQE1xsInJ3YT1XPZcoBkaTjUoYt2xPqZwIFGLoLrHDFqz5
qzKpHkIqNsbifOBD0AkcSZ2IDjurd2CV/Wh18UXzi6oVAixfaH61/+/X//FJdnfsixznl5mpGMEL
ydnJnQqTvPckAjAjahFkR/0ST2FfIg58OENbDc9wvgqF34PH95UWuTsMH2TeQ8UEaEgV8KrPmxrR
zxDSmOxdXpjLbTCtKTJfpuw0Pg/5R4L7EJBMHDzn31M4cmkJBQKgxKN0xs4uKW8JiYojf+3XGngD
3SDfoz2sX//Ww72lRonoCD1ofnwf3UyxtYA7ouYIk2YHmVfR5v1eRiGjLVNI7Vay/0xssOpLrOJG
M+I32rBYoYRS9skLKMN6VvniJ3zhI3F4WLuJbEw2TOJ6TexNutc/OwZcb4kiv/4i6CyjLrITTW2A
he+HB7ND7hrUG/zRqzCMzexUQePG0ZMoewoVuuiFnYTE/EsPgQMwmPntCY5sDFRvxfS7AXUJB3vM
ON/ykLilA1Mvc7bxa+6zT7vz0F/jnrQJZgkkY+3JXQhdnNvjWjaquAa5jemrmVtSZOFEZm8Wfd5x
dhSjmffJ6paUjvEF76/AK7uALyrctCZv5yepFKUKw+/mg7up1AqdjYl1SLYEAEDcaFyu1eUl4bgn
UBvRwFq8b6gs2K5LMBt632GywFmeIqqNVtvfWvGjEzyibnioWxhStoNlAOODUR6b5G69wZcMs/Vb
wB8lcUUZDDHcdgA6u67SaD5gXWMSKBLvUItuaphtc3Z29j3mLncaUzN7p5To/rR3keZkfPOff3JD
dn83eEgOHc9JAZzovT9+yPPn+l6CqNCg5Nin56ZGBBMNBnuoSpbjk+dFfpmkLNR9z/HbtG5uUF0Q
vHUdAqrzNNsedJiT/4/GsERkHEzubg1PlLNLRyzDoryDbCYRCdnccXs7/aS8z6mnBnJ//OACyCL3
JVMFomn1srHMgGDztR5V5LA1GSq2NEbZfdDxv6muNdqeVyVAbyedwBNyTfqV0zC2xCnjNtrum07M
88hm0yD3r0cfuMOouWRE/TUzZFGwtTUkGfcYnvSVZFr0RI1gCZP05REqNKLDWR4uvQNLiLgGKviz
/subAW2aW5kDGTYnttReLRJfa7mLW9hw5/ts3dpBbRobxqIAYjGpf1cwSKmRwfC6UFgUAAZsjaWQ
d7472uaAYcj5i6oT5yzpIKhl7cQhH/vszNVNC2UEvSSdiQ2j0j9s7QBcJW5ddcRW+nsQGAxUbUc/
tvtwJip+d+9t4o1EybIal+sxk5lekfpJFA0y9ua7O+NuQoybJwVHTodlzb5zcsZea3E515TdwMZ0
Lpp0svH9Gc1Et14Vo/9UTyQ5ayWqPvUWcJP2O7RDmr9lvzw9Q+uEhRKttpx7/NGiHVreCQruCDEe
8r08Dgi5GdnZUNFRMeOrKdXT9N019irSq+sWSV3xP3OMyB5Jx4WcnUq9rY/84lyN7JeDEFhctNaf
pnV4h7+zftdGuD33rrsGw5PCpd2frgR2Sy+0TsnPqn5MHvvYxSsz5AAhfL6hNuZyIQjMSG0/gQDq
22cv9s1u016IxW33t9AIFXhwWs4UVxM4cLQrYoCiS78bMFwTNOVIx0wMD3EabiMsp9Qr0RYEiZsU
KJRxNhUlf5rknU1SZuEpGNarEHxMuj4C0xk8K6FXkZduN3e0ytNfJowApRgMArF4tq3kkX7KNrsR
HwLHBHIn+WLU87+KDFUSNrh22dvIHyA5wzgK04PtbZe22lHIbBU2DA5gJz8meO3Kw6bLYaX+QtYX
3we2OVmQtbMRbk1sdSLu+Au1BfaVlaMjFK/27o7Eq+FZcJbGMbA8lUciEzLLOm6y2QOulKW5FJLV
4r4YSDrUUOD6PgZgexxsTA1FqIoLo3P3YhEaHcB7Lfcb9ymen9FQcpJJv4d1/QNPzT3llFg8RoVQ
gOq0B2kwe3ERhTgMO/kUXeolR9+Dueq7fHDHrZKJ07QGMDhvESZVs7mtgYXVuoNpNk3lWGJ1OBZ4
SGxDjg3uW9ma7yJKh8A5cj1mOjzWorjNReT1f8tcFQEr76axQfxHPoXYJsaa1OJyS1xMeRnb9Rfp
0KsSPdpc74w5az9RA5UjHNuAklIH0AukywXA/o/WySVEuCcWsAn1seJ92NR7RDnenpfKK2F8JM2c
zkKfssZ/6hYk43xZ/gNPkyuhIgedoRyhoOQN8PFEYR68y6TqMTeK1XMYGt06R64wcQU//T0jIw5R
kQ2Wnrhp8yqDtkb1pPQiPab2V38rxrow/5Q5VfP3G8xXZUFJxg+dOmEY08hvALcdSyRdGd+/UYUa
hLUM5FXdDF/OHauvUuyxkQvHv8def95F+cST6pND8FQ35swTdRvwh6wAX9F1nBwZSUv69z7IlHNT
y+2Ey2q90yiqDZuDsKV47Hw7WDDJjjzqfvmPKl8EVQ2pjfWtGB9pYlkzwczidgt/4T82S0KrKeA9
miAn7Amcrbgui/T2x3KsDV3zmHk1TO4xBgFKi/aWMpAxbFOB3tSoqjIW8bi9CLEsbdpQbwCf/MyO
bdMfnHFC2Arzzq9YkPlkuQctqHbgA9W2IQUIADHfFiUcJfpD2leD2/wDLFlC7kVmRRGBTSbvASf2
vncYAnPVpIh92vHPEL9NhODhIcAa+n5ZbWZ6e61DCLmsC7F60hvcPL8VHvzxWD4QxMo/+YIRXkQq
A0BSh4mgfcqKz/i50MutJNHAN2qnjXPZenk22i8dVmgscX09jKj5OI013JWTPnnEEw1sA7H4HJrZ
LcDvXHPdt2+5+DWS2vUzOop+LtFDf8F5DZ9q9e1LVOxVU2GL+RpsRfJx/nEyi5Rt4ws9baABV11n
nubPoxXhjS9DfS5kZQXCD5ui9XvzQa9CLmTNnRjItzPZLh/J38K8Wp055vQpSRqRMsNsFlyN9nUB
1JoX4n0CUf4xiZemzNmwz0qr3gikwFxdY8W+nq2r3Q9tjYZ6p0DdukSM/Qbz9eJ9JSipkzLjmT4x
G1g9xsJ7iKbp7o10E5wr/Wm2U72za/o0q1hrWK/Hc0twSSnAWm/20r8tZl1cx4tqeYAMo6TuRAeD
8QkAbDbNRULGfbZPKQ7rFFnd/QTwjRksPol2OAbdSrguSoDy8rJ2nhyEfK7NTbN8aN+uufKNvm9o
QEJCwgDsDrjyt1nUpa9NVLgLKyBKzFeN9qJe0gRqsMeI7Iuuw3HkMrF1B6iEwrvGL/aFIPQ4my3A
wmjezPysAjmbOZLqxIM7V+DHeF0FXc4v22pbtvZ7t0WgrPAUxb2kjuSOz5s1RtLOGlHml41AiPPW
yQJLR+sfFXa8iXnUPJD5iwgHNmoVf4qpY+SSH/p6qjUnN5d8IEKN4qHzdRRWqxfdEw6FwqVUWjT0
yzixjjYh9Y2vkPibzgkJFukhcLvDoR1u4AGTifCNTU+4RoTBxB041OmtDSsI7/XJSnOhGxj8zJjn
QjY1eggB6dgFxPyUK5/O73C08BIEZfbS2KA96+3HbzAbVjM6V9eliNTLl2Qq9Af4E70OL6ISRY3R
MZT6LQF+jbnSe+PvSBhyFojzIC1inwLxb2Dd+gw3ZmddIRmRuR89CbBbl9axOmDa6MGdu0m+NZgS
7fWjMxQ205cAlyYYnSNwfmRo/Tkcz36iWh/H0gN39ZLuATezoEmg88YTXYpLhpqvnN94OwZAj6V7
c4Kk9hZpw3ayZW1QiIUKE2LNF04e7HSAqxWbn38pY5tY7kQTUqDnrFMLnxaTZNH/+VqhRdXUhJx4
CxZg2r8Ue0Zwnn48npXq8cbhFBIJ/eW6ZqyGWzYGlN1UR3gKOXwdmwF7WHM/kDre5ZUDQn6k9QJk
rS0AIlRoja9GF1FEGveKAU6LxC7AOlO6IW/L35uKiKI4VBHV62JLvttWflrSrlBWaTietgebxqdy
Yqvl1xZkeEpWhkDqImNquQvwtqqfh4QEPHWil2WUEOBAdq6Mlfd9wLVQw6wVIJcdEWDRywAf/DV4
q6qFL+bgPxJP2+GXznVIkIZuc4rPXa1K9FllfmOUh/XNS6OzprzUP+8b1jlBPJ34Ak9KilvNfjIe
iDN5mjKDN/zJl2DQ3kxMJ4XMCa2BDcNPoVrwR6S0ucIdiKYAqLFeFcGI/OiCjDJPQKEwY91vBibO
BHmlPplAtwWAWvzNtPE1ajIwz14KiC34YG0weLhPg0bo4r4Gi07usv/qCerruJtNjzOP1/RbxKSN
dXAN2TxSnzyDw2EEK94jlXtTQ0FOMdUVvxr6C396jixmkLZrfI8RTz1huhPcBVWwWp9nFGY/2fVJ
R/sSSyj9GfgeYmVU+fBTcE7N0DRRyxiDkGh2IsZvNmpV1xJtvnDa0SVrWDxuS4oH/cMpAAWtHOfF
ii8u24CIs9w6QHw3kE6LkLn/ID/mk4omBVWmOq4imiX0AZuvyqJcseUD0nRtwIZL+EkzTqqnkCAg
QHNI6uzLNLJG4hc1UsxI1a/st7opQEFreHPZ1iba+mWIPGTjfiQ6ego8HBMkmimjDIlD9Pw9qYnZ
X6Wg6Ywv83V/QTPMzuwhiSvaTvzPmTS1LWztrQsxP4kfQzSbssdCJU2nGkyq2H0sexkHlejdcZG7
3ookrmVUdH4TqQVpnrDCFHJ/ce06LV9XP29sS+JtWfCfmm801p1Eer7a/xUtrYdcWlIyVGOjz6lq
awfO62UMn7f+fk8B1iBPyRQoT2cHSIEdGflQp9yIOtOMRBZh+j3FCNfAwdD7BavaiTb8HtOUUXe5
IrA3I6H17cT6d8BqFTpWlvMrsWLJbcklzbfjdOatWIJsTrqsof2AvMfTrnvr8i6sEW04gBsg1hrI
XbaHOEfI2hy+YWljNxgFxj2jnSx2VShsSQpaCfOH3lXtGLGCbcoqw6hDsq0q6cS1ZeENgFdGmMtH
NqLftEXpcxvLwdLbg8IqH4WeWp7wp47xAwVPOb7hI0RTYPfia3Rx7PoBPm1+kYXV10yoTvu4xICE
dCncADSdiW/hbKqgxqK7VlC0INeLQkM3eaRbEzqtZwjUbsCjymhKblQf0UsLP/D0LFIGxbQeCIxF
z4FKenUIhdxgB97qAN1FQro8yLUmd8/jZD7D0BIVdfGpjE9aX3rOqqovNjC2KF4miyNqc5TdIHB3
YswQeaaagiw6SLEikfsPqxszdXw3mhyG61e8jSCU7K0mqg+NGWaE6lfCIRm8R1O7XyJqwzuV2LDG
cgLe8sv5EfqBoJha/d4GbaLLTWgdjk7+N+fyWpvkDUJwlzV29IP9vK2MjDAQ0M42Ga13sETmVdjh
2/4YFuS+mRekM5HhE+I3iFaFwOrK5mCQpOyX2STzOyHKbW39LwuuHC878gDnr5YUnfHBb0djdYSv
5n0z508xD9zuylE7nrooBC0tkTWjnZKCsfqovJ1S8+wIIudNgFxA2daKohR+WCkJLSKLvYw8AHtO
cAaygHiUELlpMRwhbF90CIY0cC+s1Knbwnqbd0vAP+k4rM/aAtppnUUtpFYJkOAeUTy/rG+g2ivA
Za0aMWvxzkuciaK6YwwWn11pG++AQAp4L1tmnMay77SWE2Ug1BKHiXradsmLYMBhCmf/+DPz23Vg
d+tKavNZcYaF5Y8Ie5ViOnhRdx/y7lUAz6XUMrE5njEu3hMQlUBjS0kmoCYmXUYfl2ccK/0VA+Nh
hYDIfOYdytNINM4QjtB0An2GnpqBOq0vomUOTmTzjKaABeNX+V+hNOkbG9P3PyQPS5QXiIEMxGQi
qYpHaMZbpqzLw6+EAYlko0ZAVDZ4Q2Y7b/WiY31yjumIRl0YElSsUz6tBQpUt5ocvDi0WD4aE2H0
wgisMlC2B5OKbc9HetEhRCtwSB7rLJg7/LwZI7M4/bW6VDjrCrG74vR2V36JpuN9sa93XQGtNQYh
Rw0bXU+j+rr2KKhmJGbTUkvvbz2nworRmDHO7kEeBJJG7gyfl9SEMo4ybmpEzrX4UFvbJxAUlfjn
EBuCVtjUsLwqOvc8ZRiw1sE0jnSuDrdA2L9qJfGwFCyBHjmHLBPIPUP/hb4/ISDR30EdyKmWejJY
YTz0fyaKQHjSsSDWoDMuKKHf4nZVIyYNz+0S0cdU9+FUw2fYHgA0BkmGcjE/eeGq06r7y2i9XHX6
Ia7O6aDyBwzP91wiDY91GtT7I/NiyfNRnTWSHNvQspqWiKDg6bqDmFSRlWFBl6U+CpOSybfhUF6o
F7h55phjljo/W8qqXI3v/INI7fKuLhdj1NwRmhmogwTQ3NNGqzOlm76MHKJHpqEDVqutc60a86gC
/EzX39CVeQMEQsZSNDbrCXiDQMjFB8DnLff+Q8arakO9Jyc8xBrujFi3azNaCB4H50q5vXrrCU1n
EhzVWJe0STQCxMqTk/Ha/mOjDuwddAkBjc6oC2n8m4TCxkkPV12v1qRv84VjKM2GpIlqQ2M1qXKj
C2p+RHiS8l1zBa6eRU95kX7YuhCy0geGzNizd7MpegoARI+d3L1PABgcfDN2zKiRUfekgUK+oITh
obttUbWgDuVvRrrV9xfHGMWNn8bgh8+fGIWqCcthtS4myH4Zh9syEXuZ3EdnTVx/ViQ9d2NDvhzd
fwr/TX5LGuAeKF0VmvQLApceJ0dH5s1lrzwsDTQbRCKS1Y7eV0goHSCocELguTPZresDnDOMR4y1
7AnppJEkwSIt9ef++lYQE3aAWFnJHYR/liCyDkLC+uUsE9RyZiVNCSd3wA8jEdgany57bXHVojr1
sZis7EPhlqXLki+9d3iNDbZNTVKe2E/IMr1iVP0P76eWBsWuOmL/uyE+cRQ/FElbfwna3pA2t5Hi
y66Bsg8YFkW3ldJla56jcKRkuLQmdFCk/RsT5IDgU7Z1zOYR+IxktAfmBmNXOlIPmrSwTpfKe/6w
NIjjBfjQCj+0ouDGIkpUVN/z53NjY2ay4ung5SOhcclvdcfDkvCgg9xhBeVJwwETDU4XdoU2vb+S
2tYJq/JCwagY5t+/u5oY6Unt0pv342dgieiRTsTmWQnkMgN1Z6h3f1vduPLZxnbgPCCz0Rqq1F5L
kFZciSWqIsaaqtEapGRwdwV4+w1Zah//KRQSVlUeHQZsVWNwBg70QQNvpwvpHl9cUmZgLh89DTCg
biYI47DrK5NeqY+nVtatCBeO1K3wyST7GuvRelrJ3B1LASOqTHIXTQCsuFRxYS0oX85oq4vK2hhM
ZvdKopTCbb2OQhm1vHknyg0E5bVkikW8aG2obzaEjAeg9dhP42HkissFn+gnn40mogcxR45XB4+4
bdTJdTeWf/eZAhlZltF2Baq7QglHGGlcUBmUR+xdSOfRWeNpRXlm/CwBK/kkcD8acJ1fAUQFAW5x
Gc9a2kKL18ynvw7/IXD1o5a7Nf/2TVcCthvF1ah6fqOfSKdh81U9Ubi7+uNib5TdfU/UQE8EyyVW
/Qhuoem5Vzp7tu4xnSjwoNIqZ1kQFiya13sL0xJxPXewfw5J3RFfJNv0zUCtNMFwPGKOQDf6i4TO
jcjXX0RKPDKRcS51SWf7Qsx8iNlTmbXLrudpmk6hbk89Ly3Awm3X5gqHZXzYUIsp+XGRXxYBADgs
mNEbu96uEkWQ9mInPLnKBs+AmABfYyFKnL6sSw/ov6ZZ4ErjqwWftFfYlt1r7d2ogfrU5vyjRtF8
WNq4Ze/XoiE8PMxtOdEUhFBR9CjyAwm6vEnQCvkwvEbucovX2jlWdYDihmZhbXnJGRITHhTUrR+A
ux1G4WJU+dRZy1Rqfo/Abl9tRj6kXu76EJMUncw0HMi2gm9zqdROwsy39FgIAG4eXItRlKkaTkVQ
E3+S4JGLJfqMSKlVM5AKuSVN93eft0UfBZCChCzg1DDX6MfD2CWClVMvN09x6xA4lAS5DQtPRH8v
F2cgehEmQW9Fso+INjp7FiMde3kryX1v3t3A41OyBPeKotKtQOX5vNsaO1RPZEmg8LcgE//mof0y
Yhl5c/LRFmAte7PYxGATEoEs0VLwQWtIQKXmVZB9y5+ZHxF3T5IzWbfb0vJcCLpzaq5knwyLEapC
DmgKVgoVaj27vU4Bd5dFWLvtUzUdHRzKJWrWFBFFcTYhUVp+tF4qt6vCY3X8d7dENC5VSk9Oe7Ye
Ce+35u1UfuDKCj1V1gKuJu89uYmWSdzaVO28wNs8bjksCQtFxyWonwrFC/npbVpYkAemmd3Cufpu
4H/R0RuStQRsP5kvyRZ8lVv1XlAoDZvBK1+h4D9/0Jfz7eQLoC01PphmcAOm4L2fhPkQsKd9J09Q
s0IY/hY9uWE9eLEyaMW5gnEebAUMNPTH5btqjI2TXO00KxEPjP5+BNzaoCvKqqoaLKVNzakKnXjg
uAJbBQRKZarE3gEXqMeJVoURqSMCGAvXBb6WU5qfwhIykDBcKy3CNule9nv336IixyMFUu853hqU
nUMr4qY5DHw3pd91XTRBhGMcAbTZDQ4N6TRTrnWIJmqcIaGXOqmWKusk8tr4HaC/PPfcnpthKmrt
DQrnt/uENDXizHrY4E79EM80pQfWXCfT9GBoBiELWb5xnmpFB7pfbXv/AE+IWkxHkiabFU28CNHb
d7CmkrmtRbVrXMc4o1kKBzjBN2BAQ0+BsqSejL/FlvTVeH32tqfdwjuSokXAopFX3TkCQ0xVF33z
oVkk1tvEzqsFTTHoFfhgJSfz/GrjP5HZ9Pi0kdKkB+AfBg8JC0dEi6VgQ1sXl3QxNQvkEnZtl2y0
/AWWjZWs+HuZ8MaGgcIyo+ibcZK52ozbyjb8pi1TOJs7hLNrF4wpoguGqVfOOn1SliVmYcyziV6z
0UnDHFa0LRL91wHwhemwuAKrzv/pth7ZVn5X2Umv4bF3hfr+vAim4MTfX6HHRV9xNYMjHO7k4N9u
tRPZhz50V2MUQb48zjhbNRD7S+5L9ckcDnQy/pmvMs0rZcv/qip3MZJZ93IyYz0j7zrPP90mZF/O
hshn2lf29seEx/5aTd+erPJNc7MKXAsTTcEiHbwslbCzoJD7T/I10XMa2izw9WAdNnplZfsrJua+
dm2cIbgNekL0GSuaISG+DuBWSpihfld4Sp96+Z3c6EiYJToAEHO5Ppv0v47W/ZNBq0dtPjq+huM1
v7Wp8Qrr9ZGAGbVx+AFC7yXHnyBfJIUSIP7oZdDg3dXCR4PNXkPj2sg6m/BBhu/9gUxcD7XVSMNJ
liXXsG0pFHT4PbKbPAW77nT3XdHdzNmwj3QWklkFHGIx1w9kiq+ajXbFT00eW9QhAOFVyptHiuE3
XPwyQhbTE7in9vPlbzGadzoTtfPdKuU5sm79t4NM/pGPOz6AfzUIZvesND+lnsn1AqQ0Sy/uELlz
i5mNP090U/YLRb9+xyU3HF+r+DGvbjOho4NNPAOn8D3qZHqzyNdeSrfr1+qecyRuEiYdNzM1/AIL
HUtm5TdyMwBlS8LHeDJJXflifNZmn9eHeolLswOqklx9YQpETdTTAUCQsxIucTrDYaq16fFE8wFG
cfaQ9C+42Ete6fqPCByoKzn7Jr4N4rEw9zi6P68NQcnAs4ElxiKXFnhx2ep/ZwfMOv2h/cEYT3rB
1X1Lt9XyP/T2koxeUOWlZ8eaUKO6Jm/bcZx67SZAw9vYUGBIoTa2X943mkV/qeuzbzj9VorDHXyu
TxJ8SljO6KP+0JyeMxVayWtbYO5VLHeRCHqtgIwRcZtWnCeiXYpGOr6p+AoG3QRZflHU0xPQJrrF
mmcWgRUehTvGdvaewt0X+b3dNbf0K4LU7YhmSUwrnbVVO+/nPQmbDz/YwzFoZmgk0FYGmzSIpFBi
tsYCYQBl8LsYR2zITtRtQZH0xaeqMSpY7pNkcCDdl/TghhOH/hJnRvHk9p8N66P1Xx9sHm9Rjanb
eHCGkpzuDPKvjA9h+yEvy03eSYlKCJN67CWKClzSYNZXhKNPAK0yk0SGhC5osU+D1H7xBY0XHXpB
D5DaPbgpVPde1iaowiHblGbJjv5fwlJIV3RoIkfx8A8D2Y0Al+Pfx7bzTgv2O2CV4TKqHHxJik4s
wLxoRbhOX0FJIBuIAnsBGaGfZCU27fUpnPmct9T9WxGAxIm2AcRuHVXvNgfObMuDMHBFq4DzCzw3
oFQd2z8seYgjBe4xsTuN3shn7G0WSAD6QwS4skzWNeE/Xc+Sr8MjqlCO6ryOMZOgeuO7N5/9weDY
ERZwvHwiwVZK4bSdtuNybTyUewJ37tq4G9ya1roHj+cmjuxKNClwwfxoLj/dnHho6NfMYxpB+D2F
nQxIOmc6NivKq57xo6WrgHsOsuSI7YJm/bQUPA7F2mtS1qB2KTuqmh9X0/RsbZA0JQDPSyg4D0MB
53nZcqI82vLEx8YJAh6QONamxQt4dodjQBJBlo7eds4vMMb1zKFZ3zd6cl1NVlbne2oyufIA9PPj
vi6pq03NYxZuabYQyT6MkvDlor7JgqfPYVXs0EJ4srixFQxH1nl/ln8MQpIj/vgp9/vxcp2n71Xi
oCFf1hCNurZ/ris2O2MPHss8tuhOP+y9Tx20Iy0y/FqcEP9/5jO7VhYSTaumMt76SuWYv+QbrXUz
kMSaJ57qyQVCuWXpzuh9unTeekw2oog/bjO9Zdvy3ldCiz05J/dxWr6jgw9jceaS3Z8+nt8D4B9E
/h95QSWr/snL3TiRLsE0ixqtGlYfKzQS55QZ+rcOWH0DxQOEZtp2KMCSVVJ4I0xAEyFpKm5RXrkU
KyhUoPnQQUW4+xRyWO57yL0ImiHjKy/olvA6eXftEPRjrAe0vYQ9JdHean0GlbBTYEkz7P1Hyeja
wFoqqLK36YKfoF11IQ5hk5CTJ6OItK24Me0kTObGwXwl3SWxQ4LDMwAqWc3SCJRv6MftDAAGh0Zy
xCV+Eedy2w1hW+41VweCDqAGhlRO/5DsaClwN70U27zbUbH07OtA1lCPRneD+4XJQBBDqh7fpQ7b
LKxgszUxYH894SmMw8tJQCY1ojaIwR4T77Y4FMOg9BGjCQDqTjASMEegDjARP04yFj9s0Zi6roUo
qZGmtB5bNAueXOBL6txYVRaHunoo+LqsxCMWU5wBR/kL/ex+D+Qe56MMn6pk24jAwoxl9PPnmX/o
KeuICL55okn90/dyV76Uv/g2bodwWm2V+zR6HJ8pDFpE0xBpOsViZFq/LooCVw7Nvob5AdLhIbD0
mVVnmSwWJWLe4numH3bEhk+cYYAiFoMjbxKuJ8NhNR9m/2b4KkJi0lwheikH6EXJz3HjNMOg8szE
TjLjagT/nGWZQhhQg7K30aGo+ecyRZ+9uW//GPd3FSKw0/iadhVj8iTpNIEfeNX7seg7gHoGT2bI
Tc3YcxNsRR3dlGi5MIlZgTsD5bvsqi7LKo0GXBYW75V1hcuCsiIFO2bzd1wpdMdyf+ajPx5xDit2
qLarIyRHJWVO1A5HLWlBDd0//AaPS9VPS1SBHrBBoqAdmR67uMiLZOJOUd3Mrx2wdnYKBYPVW6r2
4EcsA9Yf3bM27JesPcvhSaUJIwK7+MyUBaSU5E9a36uNj6odY/LoNYSJDOMcJykOrm8jcdfeyoWY
mYeKXA9uEY/eAcVyJSFvWKwMhrvftOJiDKmIbht5FQGPNVdjdx03vC/Kz+qry6mSUFlzK/km3vxD
SJHH1l4Vr0aw7GWoNtJc/jmhFRx9GEdSb8Y2KpT/oWo78+E9XA54Asq0WXFx+fidjJaa0t2imDWJ
AmZlDJlTOf+kRlYY4A0esJAkmJ9RbIDM0txpPw2KuIaER0HRx5aRLgRQzGuLXIW8YJrq8uiZQeX9
0PM7lS6aub/hYzjuavP5rOT0P9455glQHKoiMKHUnMhFah7jB1Ql3xH8FrOZyj2mDAztyBh6Iome
+VeAyq6+/3sSlyc9VCndu8Vs973EmlbKqMl041ejBifRKyBiwrm83wqVEuNkAoAxJlu1qKerqrjz
uU243R7UsyNrzNQ8PKt00UbW0wc0LEUkxO5NE5zg16ASzUORwgzV92nzphZ2JpvmF/axBtskQWOE
Z03sgurtaChMylpYVjkRnyCQONAMb3mmed8FGU0U221GH4jJQmRs8Rgg1DNdbKOXa0JkioBgpIbL
tp0gvb5fI5z3CjOzykg/OAsUrQWsXiPzZKQ0RENIq+e8sJFrQGEYwHHyslG+vSmgFoXQy/pwqQgq
+6pawdJTD8MEbtpYBoTR+THqzU+ftc6FtPq2nr6G4uQlfKdUXjZWSH9omgj2En34z5jCwrB76emZ
p8ITTkjT/AQW7BMUW71fxrMNsmX31QacNpTeGDQSk6KsQRbiM7mrIt3yv0PxbWxZP6a4De2gZEIy
nb6PzHl+OeXXWR8o7vm5dQPSXLd4ySk0sJlCsmdIrCY14LaJgFDZalqyB0a6iufC3b7faWu49Epo
Y0etOxMEotdxuHempjIr4R1GT//rfSK/FDoWbgrnfCKNbuGFxa/FGl/7FwhNunEW27E1c4JbFn0Z
SbeD9gUG6AV06PeyvkycB0JuMUrw0HJHzoDFZYM4LZDJn7FxwbbS1j6vY+8ssZqJ7YnPcNcfG77P
QCMX3aRWjlEjtzj/uZjI8H/zvnLQpVvzmUibiPFJrpwZQiJgupFRoP6et/4kVBC3qSO/Q2kTHHS6
kTiAXg89Ly3BA9U59iozBmmYWzh78JVFINlkhRaXgWR95hzoPSzOCJpWwlB3zLuySh/nkkbGNU6X
fp3YDbz4dTChTD70evpzHUIedx9fkG0gUyEX+pb+OhT41OhPK8fxh3SmQwfK3U99KwECwEp6haRN
kgumEG7sTb0uuS8iO286Z9JJJLl6tR3nFX4g+tcnvmaGDr8kKeXOLrUgfARGoSfwfPxkYxzsY4Zj
YkhCMkEOlZc9wQDFyUX7uoEzxdmPU9iOvq7yiDnz0NzJIJYGbVoOJ8vvc/lA5KNxWMMujfONVseT
lz8aA8g+OTRdKb32MIPOYws2GtiRCbVo//09FqVVDyHTV+A8zlGjvZDG0wZKPGnnX1+7aH1Gp9m3
FK9qtkgvG7A5HamugtzbA3nL69IAmonWDkuS2XUSvY3GJt6qy8iorSt7g0CZJar+82gO3AYczbqE
qND+jK39UVJRyzjTzCz/wa750/MQIOx8pfCAmjhc/97z1MeUR//olTppb9U4h+N+3GIjEpIVR+/q
WVt3usK73M1BEjJEnPOZ5v5Nb7dPsKi1ap87YMDTMlywVt1YOZsbm010V74v/Y1O86g0PdX6eVl6
bwkqNv3Z9L1pQdUNJ0iuxmpdcFvmUeyCVtemqwDez2QpznxN9rzrRPeA7RkJLsJCpK7/dWvCyJJ5
TGMZlj8EJLTa/qdi6jxhEsJuAvmyYm/Heh68x8tkdb6G1LDNsUCKpLLMHClR+0ZUbAooKJAoWxuZ
fJFmuLkBrkdmauDzkbbg0BB9FC/tFxvAgT5pmBG9VBCjFYwr2c/tqho/LXFzLFoMUYZLPnhoAYOD
KVgYPyI/FfdMnIn31+Yj1Vw7b40maOMSSv2Lkr/Wpog0SH4CJ1ivyeEsh6XgQFKObsmxwfyeWvZJ
jjwd01/LoTuufxxrDrjAl2N1khmb/5OVu+5gsj5FGzKEaEKf6w7ZXD2JQcMg+sM3zfAYNC9mfCy/
I9S6BSkKDU937ElRUUdKCgSb5J4wpQJUbk6QeWARwvttDim+BwPh9j8TTTvutnoBznAAQEnv9P2z
pdxZkTsotY8t2YBcgHwPPgDRRKBOCqacgNjM0Twfr0ybmKeUz7Uagi9mfOsL0oJVDZGUDg92R/ql
CDbhy9G2M73ZWGzUYYJSPFkEo+GqhyXojgZwKKntonU/Gehlx5QcOsJR4d9Fe36F4gPsBV1noU24
lF1W2/fVG4UHX9lKUsW8XAkazooQRTNFX3FbmKTT/zHgEdXaTLpnSSWpMilyeLoOw9Fo30wdd9eP
l/9Qg0Y0SkSvNXAlm960ZXTeXHRM5Pcx8HfrxLnfXAqhPH4r9gPsHvcElDg3zqbh2FaFT6sT83xc
go4a10BWIaNBmuHN/GVvQOlKObQM7xBufmWihjmF/v/FotxsuraIc3TomYLmQxxXw1xh5J1msgpu
RbxEfTkvt+T6sizH6Gdb0bSj1+VW4Ht2NF+6zmyI0XK6Z0aHp+lRQnRJ4pLA6W/XZHgRCD5cjfGB
huLZ3TFRkNHVp6yCbOW3BFKnnztika4h/kBEjLlbqSpIlvCbUB1Xek8PPgbPQYV2aFZwIBlJqTuU
d2eQx3tbp3IU5N/OZREG3Z3N7QyokPDjjRmAh5ioaTQvesOJRcl3KUEnG9Vr1G44TbSPMzfPq7Ek
V8D6FMsIQPKRd5n+yIVx+mYvMJn5ArxpbvF+yF4xKqjnYwkaTq2oGPVs6BGQzbHspZSBtyYSA9Pb
v5JVAtmGXVu4KFkU4nXutqthBhD6dV7kwM5reCMXokhtXJ7zJo/klZZf62iE+M5LRjpEnKSOCcN6
6gC6MDQ/H5RH/YVwstSaIyS8Iu6Oqkfw11FKrKFJHc2k0kuyN/ufWkUjkl/bwMZbM/zRz65/wN7u
ZHq/Wvo49bflRrXSJ8v7SwpnmdXYqNSdAHk7fxx2gAZTChHYojrbvuqZOBUWTVt470mlvA2OPQy9
hWhTTFWSsKbHeVWfY3ApdA9un+1sND0GAcfG/tj85yVA9PnRnRDnJ0dGhde6TdfhXCK7mSj9IxDb
RsTOz6nt1hjmtneuPzZzaugORyDIATm8u5qCc1du7MXMPXEFcTefCoLbFxt97j/2taJ8w4HuFLY1
ezvOIx59au9ehXEoOD9ruRyDXPDcuXDPZW66J3+vawLoTiLNlykrE5b0zMwh45dye8IKHfhaw4ng
8R3ETI0owfW1CMr7f8IBAxJJ4NcTjQXsh+sIEPS5putf36gwYqu635s6J42rHIuhddCgSxkN6j+Q
ZQRJBbSbnEewTjMtY/h07hf/zD9yIMU2/MuD0W8ZlRtKEp2S92WPLXDBYwwK54zYtO6lBR2NH6Cl
lmnT1zIEBWZk+3BEruyr2pOG9eaW8MPN5ICaZaDW1hwj+/xFAT4jxdHQMSUcvO1BdBwx8rP+JiF+
bcPwMzqtILdN45CobdIhJ3WuhmW2awV+nQrHiaqGNYmAmgkLintHsylsjaI7/EqrE0PO054lmm5r
XPQqr//pd1ljVoV8OMgYzUH4FsxFVC0vZoSkCECDbQtQeNHjSbS2qVuYMR2zODGLS14IzgNih4cT
cbxuqX/Zvh8e5+RnZdAVJOdTOneMlBfNxn74o3TJti48WSjhq6hPM7iMIOU0vhGrDEkPW6Ess8aC
9iSCbc3GczDjaqqk4BwnXSHlZh39xjG/MK4gJYfSiz95HBid/t4PxF/fjedS79QzUgUyU1Uuy8Il
IvzNz7wDkGleKwJb+687g6u+DayVRpG0rZmtvrBdylLrblbKt0F6hy4ekkWCXwBQh27O1GfdR479
b7/D/mTQGy85VsWSqxOvfaD3HLUbTI+Tv1yCkilAxFXCytdv7LWLN1so3bgScD6fMLmCW0nFJOKz
C9bI32iUjLSZ8yTA7JbIXzL5B1pJZwBPu0CNHwxTqn6BJDYPpiK3RB5TlaYOP+PLyTLAzMLXfghZ
U0A3oXhsTd/KJJxZhP3ne5qk/UgmUnhG/RWrX1yyYqYsF3PLJzTOojg2E1nkr0leGRK9RbQwMROJ
BfRHh7tSIIJP1fgMQgMIZT4TUDT0xbHzHoLKJ0k1hqsyiDoS/Xel0ZTBpNHnWh4nnxYpo1EcXvd0
xumRng5MRFiXE/G15tUWma2ORozlkwHxzZO40nD3CDFoiAUplCm9qSxGe0/+AViOElx6Xz6dIPmW
VHGxOZc7BbYnRvlkPgO9PlfCXmWv8l7CHnVheZHTI1oW66S/NaRHdEY8yoj1Qbn1RwwqlxPFB9xV
WyUYVWniY/dTKt+1l9wkAvcvuinE8r5Jl2rfy1hMFZ1Hvbb+E74oHEux2a2CYJLrUSXTxiK6rJyU
OuejlEAUTQkBF4gavhfiCiwHqhVR3N8ZS6Lmz2+40aDoRl+srD4y17VugI1KsScFvnpTs+7KHOh+
glx12XwXq7EVyNj5bhbbrfNYn9NBwyvBW/rkLSBCB2j2kHoo+6v7nW3TNviB6QhyPUIjpC5et6MQ
kmw5pptgVRQ0kZLJYghAO3mhkpGoy0jq3TzE5w15NAJDUJKGLN/Qisp/rgs8XnaatmFkq2/SPdl8
jkIGzk5X5/o8Eo8b2eCiAQD9nvXO3wps93cge3h18O3DuoMkL6hEi2i0OVItS2xzxydNRek9EZwV
rVqHYIP6voJc8F2VkaMSuxpw+N/brN5lwbke8FPFMwLMScksYHY6u+XhjkZHJ0dhEC4cfoSiiCxw
C38tr2KIEqx5vsuPFGmn3FmTawB3sDUsd9htKRJLLOx6REYegZCkvuy9M9tzfvVhbZn3iKJ3s/PR
t7D4A2XUpBB37YVRZe1qpWxeBqLTT+kfoVM7SBuCprlMDFG8CMdDTVJe38vSct/lzJDQIXVb5Kbw
Q9gM24yBhvhb2R2aKvKdnhqLdq7etiFUmACLa5ISWIxYU0OBzZO//mRNBUCLUs0xAmni/D9xGZli
C/OZzytz6kYkmdgx4W59PvDu7ScQFRH8F9Nk8s1T+Tkhdqkisu9b0w0aoZSgA0C6TubtM6mM0VJz
lBn5ZpRQXbfbXoo4dN6IKGJgzb0B8B9b9zJDuziP9PKQh48qEqDFeAODAXhX2SwLxXYVsiNVd7u9
SZd1THqyvDQbSXN+usJQkxQ057hiZ/POF5cOrp6ZMu4YxZwPVMy/PSGo0GHZXKnVCUnNzMPa1qZP
hu+JxhuSrNdupdr9BNIWA1XVhnRdUW505hifawFl9IXebpTS/wq7XUGANpSd0IZdFObbo4bX5hDW
57YiTKvksV0nll34Ko7pvkK6JWHdspInq/h8bFVavIcRwEXiPzmtIwVfQWW+X9eN3HAPNWYk7ctY
VmQeGZQpQtUwFh+3c8w2DgguzrgyuFKoyf8NoK2ggWkdYA6W7QgPVXi9XmpqVadKjhDKY8WdFpIK
RuE3SBDMnCJ6suG+fqfVoNdhYiMBtHFyi1xo9B2cFfmYNg01WLKztVCMGbd/Im5Jg+d7qrbx9cYO
ZNuAfMdizabEvbJ1jfS9V8dsy5VtCUzMK1x31Zmf7xlb9wutgWKcR9j9Qj1Cj9w8HV62sMCoRLuy
HKf9EHLUuY/ZHrqoo6x6N4ePiQSVrBurPpslnXiaMQiYx2aNT25mUmYV6iRIN1kXJ/hGM2nir4f8
7yUFYPHjmmRUjUtXedOgo/Qi7HLCH0rILrouG82kZhHE9AFzeWIOFtsDMmSyQ6M8Z9mE7ZPikbu8
3UJIa966x5FpXmU1tgsuN4Vd50in9eHbRoCoZARkDrrNag5wiblQSk9QuFhLXxXR0XMNUnTfbtrl
uZoiHwCFXXrDRWjk6/NO2TTICSIToApr3nkXEcIF0I3CE88e1KJ9m4r8/NWgEIXt4sLFNFDkAtTP
e129spLIuBdUUjKcQB87eym2bexTw3jpkgiO7+7vt69mCo2AOGXpEBxuiC4jkheWTmtNT1ZvVSHa
6ugBk68YIQ+b4mW4QrHNTr8W4pu8Qz8GtqOAk4YedIIMjewjGSKNDKWELp8dLBPUglQxcummFe2j
9Kt1dJYBYb9KfAYtPoztkib9We+pytQ5+9bIj8CjUdR6UudLxjZTq3ZGRi4F6aYjm5uogoMGzK+m
CLEsen+5WgoOdHL1r0j6vbiYarKpRFQM3aJ0AbMm5KFmKbAxrHQLs8OJbIrcIadHlNqzAviMxrNA
fpW86GpA8MFKkrkBuO3bRoBI0J5OIuhBN7hEQuHr0vYOCvHDjxiK7cpLQPMLoxHoyHRBnhUqC2PC
TrgzK7+UdjrirgTU24q6gHSjUcxcmsWMR6IcvSHSBgCESvFEqbm17y0rHy0O7PaFHPp8PRtP3sRE
K3t8S85FxCOOV8N7OMwTVmfZSH9fsP0YuufOsmAeHhEzEJ6b9oSyhXIxu5ywafrZgqEbjoa0/MFf
SIj09WIv5TAbyy+WbH4Lhop+XjwjOkETU9SRW0FowJvFbTQiIIiLIbPWZzed6TkYwejXgAxG88bq
YAtSReyGhDtFjb8ukFXajqX/0v/yNpA8x3jIplCzr4VeCVKqZ4iQKMVQjfFhHcZz/w6YhKVPBoS3
UuqeEyuaKp6YBeZ16yShJMWO3sRxxNTs0TYXNRUeqt+sq+FUk7fAgDn307Kg+kHOGuYYhxGewy0B
t79FanSxsJyjHz8YF6JzigNeaZqAZSG+pkOLE8hHxHNgEp01LiBt0NG6mvbI2QqpIhQyVuCby55N
m4E+0xgD1uFR6oeSrSLPMenKFW/SDhJfKY5EBukB/qAbIX78vkSEMg/KHDTnNnYnMfdyDeY7stbf
3D2wX75mvGWNs5IddpuuG/Wbx0cumcVkfXY5Vy6uS5TFEsUAI9xMonTpxO8+pijjlH9CwZu/nLtD
DDliGC5wp6IZ2YeZrfxY/VCT0FgzSGSuMCiT5QmWVPe/chMvNWTgKN7zwhBUFeiqQRz+wDMG24jw
o+q4QO1zqa5aRiu+4Bd5LbxUWROMxOs5Ixz5CUCEa82ipegCKhBKbFijOUXpc4KEXUIhj20vVyC2
1zwQe+RJdaEQgB+YwX84EUsBgK+CpW5SCVsFAI1tvYrb6HfpSnRGqcYR5fs0LFXrUKTqyotBZ9C8
kipRIPeSPpu7xYtW/20iLUUpbyTfEDflJJLwM5AN6gR5Ny9cTwKPOXGkfUXvADYEbypvCZHRVQaQ
JHI3UaokAf/6yKouFsQVAJcr56nzphyD6FQW8tpJYmUDsz4WNrFPLF4g9s+bD/nM/yRHFJTptdMu
essGz+sC5D+yhJBRtD1fA1jz7IkC5wsc/fIUv69C5B2CZy2JZaKG4Tcmj6EWvPA+iWjyT3oFiFCL
8xressv21EnhAM2noAskUA2livJDTqo8hBkp/RKeITnPQRB5aT/hjeGbixjYX6oqIFdH+NyaARzh
URcr0CO+5DNgGHjnoTcOzMEQoCkalRZmyIkeArIlZtUrL4OOBD3ZZyx431BYf4q7Wo7W88rAMWjg
n11j3ZmOUtqK3wODk2yfhLgZi7NPsW4R1wXKy/6T1l+TxDyPv1Y6ZZxsvCz8D9OPG2niSi0OvLdf
0EaBFNYOx1V7G0KF31NLlBZsAmqwFoopYGhTJoznBZwIEGN3pAwtfIHqzoRx1M9i7dOa2A8y9YmD
qM751t5xSV2lIbvM7ZglgC5UkVc0mYo+Zvug/ueaQ03Owip08sGAe4xoItbRoVLh0W+9aCbQk6ed
hVJgxLfPiD3ICBRfc3FbICs2nl3OB9Yt9aLkTenqplprxJcIb5gyv7cVvYz0KVIQjMou0vvVaSb3
i7Ol53iX4z97BPquYQSYaxPK5D/wWeBfhJoXQcXoxiCaSvt+bj7Gmoufi31wDK2St8NWPmqF+mE8
2DH0Gqj19d3XQbmVlARrN4GYXJOtsSx+0I1WYZ0bSXy2lch1NLnePo4dMfL1upQnT0d2oCBSRECR
3FaIqHMmvdYbocgjEhGlrLvx3rTo3gr8d5fscTiTGOvA6Ibwswsed6dkhbpzXRPFvbTjKpw1sE5y
K1kpp3jUJxF1fQanFknRA7DY65dcKuTDmECjtiXb8Blks6Cqah6PZbuRX79pON+/JdcnQVkDLhJq
x2Z+T2L9HU8sGgkSHG6uo1Pv1Q0doPOhA67nCIX+ufpdppqb7oiIEjrcVx8y8IyoCYuIlgsz9+1D
V3dKWO3ihfSMOk5e4dwPqkywl9UzvGN3w1nilMhfA2HOdBsrGt4Pm64jNx1aqBK99tVNd9l6U6wX
uROY+qhqF8saKHmRJht5gdZWbw7jlIzuB2MsqQq2PdO6eSK0z9S2IuOkHSsFBYMsFNVMSQU6LFFv
v5EYEUhG/W6+j1Y/q7e7nQ/Tz5fKZM269AywPoEid64ihyATOu5b40uycQQ+9mvsVsDnW62J2wq4
VXG79msRksVPaCI5r1VMoI2C70xrgqtSOW1blYcO7CrswbyKr7fE94XdiXRq57waZCkMW0eA39dq
L8CEezPemDoq324xL8nEBfo1yXU40ye6h9tT+//MdiI2c8KUvgwkZjyxtDVEpDMyRQo9EGpSjdKK
6v5XOSsYaTxt9AscNPDumPfSUrstVFfWWg2TrDVjpbD/KdTQMBgi8PG98ueptlHGBOOvu8VDxKjf
L7A2oLxZtCGXqzCCkNbwja5n+SK2mFHmDod1wHLXKsnkRaFc7U42PKzRh9urb9ws9XzOU6A/8DBm
t6hPqzPAY9R7wbCqM0U2UC+2BOseUxB2MZHH1Rvsx1AIsB3Ly2YUzl+uGOlbdftKalqZ2jcryTce
mYh7UoaoGgK/c88xdPUMDnmhNaL7++93YST45OshC3unSKIVHFT9bOcXr98W1laazTXfQ2JJmf8L
qm3h9Wh7DasOiyborqDasMw9b/x0mFOyPoy+XU5QHeDg11QwVjr2RDD17uW3v0OzBbknyAdpRUlP
hGgBOvZ/eIusAJnL3UPOMVDPlb7XImvm8cCCtHgWzirVva8oyjS0jmtCFnd4DlwiDYuUcrgAysMP
6A03f5luhChbdyRT60FDKB5xDMZcKHxY1lBP8/+tpTUIFSfQRc/bbXkqF/MXcMNxWFrdPkuERRka
A6JvJq2DT4qBkGw7V5zk835ulBF0qixU3wKQ4tpED5EpsLuK8z17Dpc2DjTFhfvS3zIJDTtANy7N
snrt16lcXmF3ZMJ/a2Q4rZDCXzFmfRL3R2yyTU9dglSgogVrq7+JFzBWjVzO4Ro4AK9lpb9Dczgv
mRqIg6+mVPKRVST9sB3zG05wT79XzHVCrEUU6QhA2zmR2/Oh5gyHfN8asNQaOm9pt7NnB80l/Elb
W7rkjmbgQNhKeSNlHDU+gIIFBoe0Bfla3Rygh9H29QQ5+oWc9I2PX9IWY0mMI9oeNRxe6aIVo5o1
TCvtsdk1wARoRew430OskucmIcY38QHqjs3YWFRYlUfLWmZuCtRZ0/AJeQxQuWz8D95jgzxBC0Nd
hmgEZHtKIPplumOp/ZqfI2PU3kdTr7deGDXbOf6b23JxTtbpIwZ7BTT6LXibKKigKluo1/tdf1bn
r0NyMkkS2k7TlZxidx5sev50pbiu7GUpRYJbW0NamIL6/P/yonK7ufrCwDgb8HLUGQqLoLgpK3EV
/x0GfC2UNsVg+FxpRHdwdCMcXBeAkA61cK7lSeo02+O3eqSxtswNYUh9+pgCftuvTJxPsCIFVyhw
zFEAocSQzQfNojIV0iPoLLtqpNkvxfE3RzHAoR0IyXjJkdahGK37VH3Jl2/9BnAU+0u0c0JLY6Si
UoriUs2JtyIuv35/cZU4WjrWmUUfyJOP3FXwDILaYbyD/DmPEt8AIMaJsTEvNZdmyWIWW5R9k5YU
8apdFUfH2pSPOTiul2cT/XYHicc1IL8+sw32JFFy+5PnGiMDwaHzUQnw1nO88BjFHximuKl0E3O2
e+AZj1SD6En92qeAZ4eQZJI6LG43JxISG3+77+9+MDbr7JGNOWQRmnSvxPbM/7hfBpMv+wqM3SE4
ir7UrlaxdWpTEq32V8By2GnsarrXlMrgP6jg4M+yt5+luUdqH9A0NPLBq5PVY4h/74odLaxHBVUb
Gi8mOc3ZTLBPPbM+CTZaSXiucjuH0MYuC1ldVhG3USqKvt58GCRDVWYHcLV3iOmK8o1WvjPzgguS
WA3yvP26goEzBepFRHadQTGM5yxPPauSDLE1F3N4uPh6Aykns8CJUw2IzSyYw0sOgJ2DS/pl6vt4
Hy+wkwKvPmTvqOGpYR0IYgQVj7IhPnJIbzXk0nUel0lJY2PltlPXWbkFbqlI+YNKxneGd3MGGyeK
DQr3AUQACrxjb32px5vX0TqoxCNKs6iMpoK2vch1p28Yd1vgAxQFq0D7kXRgPUR6joXNo2uW3jET
vpEbjOy3YSDmYGPhabcHTypni94u6K/95eEhRwYxSenS7nncLnbU25QTmznI7g3AyYnLvbeeXPeP
uhYcbVxt8q/Fu9PUMMjQ4JMl02A/EUkgpqERikBuldAtG1iVBHLMMYSlDaFSmDTD7pC9/FgXEjfl
jW4K8JIGTJgnBKKYz2ppTzmxbt1+HY+cxalnStbYBemefTICnbCCM7bIA36CH7mWVDVlrwqXEpM3
uUGqnD93/bsif/sXkndMzrZagLPDGLKjsPUBHZPJx+HrAL2xdfzodO83JOpCvigAp9Zc464vNMJ3
osLew8tWm9MvdSHci8Auf0c9Xgv7rpcPErPKE2QJuaRzU5UqHy2FHvz9EqXHkAiEuJGw5VKfCest
e46xxzvZMCF+lSryckAJvrF+QJ58ECkB/IDB3t5cumsoBdGFe7zcUzFYgwCemLD1CyFzhYPZWm79
Akp2EvKZMM0Hx5StuuhIPnOgpQLnW7QGbJ5hVp6rcBVasZOTBux4fxzIrcWDq7F6DZAgngSIrL8m
omzUBC0Zm8sWdqjUaM/wA2Wwz8J0g4vzjUxce7ZEa8jMtdfRUneF5o71VulTnHUR2eR4OLwgV+lO
tcLRoWSbA9kfG6ukQAnNkqeUhqPyL5MiqSA7FlCqDxUYwbSeq4NO8rVw8YUf6DiWuyB7xBw5ji0h
nc3q8OhFhZaX+9Gyoz9U4qd4+snUwOk24xb9BfqdYjXy+y5N7YY1iFse/pIQi2NH8MiqyT17C1lw
0bWXsbliasl8BBYTUKWZ0ai53Qzoi2nl5W+nOc4GRFqUVUn/fgDgzzoHmpJjBq2h6LhWnImtvCUl
foUa1JkaAkfbO03B1XMJV4U8NLS7fI2U9/ywCmwyNY2r8uZkPr3Aamyi3Jk+3RmK/7yBy3RotdI3
ewTdxbGkd84p8CGqRwrD92ujUK7XDJ24pDSceJkl8GbR3A1xc1p6joDOc5lyDNCy3U0gxHEzlFcE
OBNXBVckI1YfkmkknJJ05E5+CG4ZIeGyNIamKIAjAzHrBHFzRbBkEqlDNMAfjVIhE4GLEpZm9dhr
cvrWOldilXv9bE7Ji5lLplb+Se4V3nSwsXASUmFy/JrPu+vaYCGl2IJZau0B4qbrDsECrAySxTH8
ZLFga/uixSg5BfgEwBmFiQXxrumL8LSuCBTCamjCIR+gif/+OB5SMAxJ+7YzXzOiu4aGFS0PeURN
eC9lFXAt6WQMQ6an1M94RziY/MhVqzu+qmWh0vilJjBohCcsFxDRs9esnx5YqRhvu+lMG8VQTKtd
5SJSRd/8EBPrhEV+3VwjQ1NPsq4kyyxCtYQ6hEGX/SsHn611ODLAnonwyS6xLxQtCGmWYF5wETMt
jqmc8ABa8fem4TlI3ksmiEJ1cG2BURFemGNgHg5cQhbX7P2MT7tFyEHtQxszZK/W/45oAaaPleKy
NCwDEIgdacd0loQcJXg/3ob9TPz87kJfWDXJpWf5Uw/OQNpq8r+QiC0B+B6ZJcWiuep3F8cG2RQm
uUSIdxYGUcj7vuDMJfu1d0Tnu/UT7SrL2j1AXoFeR/LK6P8R7H9B8F2TjqxW4tLcsTckLErkzL+I
Ez5bpc6fRS5j7xAqMJ40CvzQPOlLYryauZADqBs21/XxUTrzAtMINRII4rnRMGqXd+DHES4y2MtU
GTi2/BzSBdAFZnF+q7RVv+y0blGvazbfB44eIkKEtnaUGnataCacdnLspp1JnYge8paBlHOMuNCT
I1lZP9NjQyDw+z+/mrkwBcdns7zLjy3juTW9C3V1OYbcjVVJpnjR2k69Jcdei/lj4K01ohkaJbJJ
TdiVgV4AGbWEMSXbSVNPlVDiyjepj4OXMAFbNGdv3zI8DwHGeeCIJarI3LjQ3/PY83bzkp19nLdE
7Cl2J+33NpF05n/vHzAMjj+igW9hzzTE2DknkDOP0+hAjfq2ZonUlbEr68jrYEg1v/Rk7j1oWKbY
PCMZPVdOg57gBATqsrVnQAHj6sDpElEDIXdrR1rceOacuL9yrslDCtzSIAvm0vl7IYP+mywt2itH
Rg6wSfNbiB5c7PVlZD33V1l9uNk35kkEplzAYwcqnVhMSvDNiAcE8TqZAw1+bc78Q0bYT6xBpr7r
nKwUXsjGIgJpbWEv8jjM1dL34OzsfBKXw9Z1iqG0yzVVNi76zQas+VzvVn0meIuYSTRdydxM1Wez
0ypMyQB2pgSE8eGgR1KRMvFJGE/yv9KaA5p98v2X0HQ26WvWcgb5srLXyc2jxoCl76DlIQxCy9tT
nwtqUCH17n9PSXMtQ3WPwXMxRcCGZsxsCARCwovI64ypvcmEKT+yjX7FVfw7yoesQE++D1cBHJYI
418QPHM2vtzNIJ8XUZELGhwdTRniLyl3CmcoTLpWg7qikQQv/MzTx0cFvbMJBXjXLzI2VXDFR462
6Ezx6I45DTT6Ejd3yh0FQRFiR8Xb5Hoiqcwo5Wiqaylr9X5UR4uOsTIRjJyS2EY6LZWOW5qTlN+1
+MKCjx1TX3f0asApYtzf6q/6SYi6HuPfyUThtXysNbHcuyNkAnYx0wKJ6VHHh+1fkIteG1AXokGC
MFWJkKsRq8GEqEuIDe1Ct3V7mHGlc8VdydHrYSxMTs/thivPrvg+ER66Q3rmyaw8uxWF52aMqZ0n
o3tEjQq3hyYvWnfNZ5X2I8oArBESFimUiJB6gBRbFpBlPBn97sYS2Dn+POfb0papI/GFEuq7EVup
nJ90bvHmIjJMPvxptcF5hLDrqtsfdAmV7Kya6oE3WL0Bj6L01pSJ1E395/5NHdseIz5mBRjMgYvF
yf0wjA5LHKEWS8KbbKzn6odaX8tHGOMJ/mAuzAlJTja5v81gaej5IgMbrHtqE+4i/Gd1hJxCldLu
Ltyw+1mlNnfExg3q7Tjgs3Llp6TWd1wJNA/kMLFXotq3As339iBZfSwyy7TUETmGWrG5jf7ZiReu
V134PVSpjdk47EY8eXZmWRN9lVnvHuEzEjflUBY8TqT5lKR+1LEim4kwE0tpIFcsbIQ28wpb6tGa
bw8x0gaH9nfvuFztKb8CvIeuW0+2eR5pdMKhUxnsT39nXl/uII4agvQizdyHD+pJbaHOm5x+pIJ0
bTYXWn15jMsUFZjv2yBPZaPXYY55LEOyjyj31LK6R0MIgVjea2Dv3YkcLlzquGbudjbW/2ZCs8qh
ChcxwYt4oCATrAZFiT0vxutA6Gs+P1icpn0wTAcbBlThI3ygy4ALKzpTpu4YEpics6isv6LGRjVD
gxZa/icw/M2nqGe+Ro9/lzrKObeDdpfB9xZapMZJwIUrAoDuN5zWENRMsHE0jYmmXL70v3IQVLWP
KEL+WiBiMd+ronQ4iWoQEzZ54f1C73UGgPPQtD5JQ1nJ8rrcXRg8uv+e3zHWxEc5kIg5vPG0ORwQ
AZhgFRMYnQtS4LwrZbDGmUV4+LN+CM9zyDZcbjjFig1Cj+Q5kksG5Ci6D7FPbybRwZIs/+1HG8bS
wppR7hAIPPCaOv0zu+DN1Jm73/H6iIQKACO6IJjaHIBAFnzphoaYsFE80gV1XJFdxF+o5ZkvQXgf
pcYxfqs1Hq7h6TFzDtICJgV4XtFBPkZPBZUreUMYp4y5/5Eqg5h9hGiRJqkd7cAevf0hnmpgySIE
QiNLoYqyeaUjoMvXD+3rUALQc13aNh4cuaSIrXx2z+fqwHb9Jt0zTWbyWHYIJ+LB5af4s7u8x+vr
Wb0VHT44GSI3xXVfL3g7KzgmThM6t2GWqhmsQgBntcEx9huyRnCIeWRB3N9InuKZE+4nR63JbImL
5KmyucW8Zw3wQeWkNqV1S8+AQmlSDHWdipO9BzuC0g17bu4P7gCWnnAFJMUYmp+DzN1yvPjj7iUd
Syk0uuSTQpqHG8SWJbgygGnXAVS8S8DjFNJeeVOBA73UA0Lij28nqnAFGG3TJNJEr2YJ2tMqQyDC
zjGvbEcTwtsfdMiFSIM62fGTNTrLq00NwLZ6SbKXPp0tKWG7MFkt5ntifxlrKlswnkO1cnn+hCun
8mlYIF4dKxp6IjlKzstrEFtYcjMB17Zs9kAsTwSDXkvO1MfxNPRIR3Ac5ZHzCPgkqcs7YP0+9Trs
GdLakm76vL1mvGmzd++5hQnM4f/hTVo/iB7ht7XPfaDYqOc2Ye9d9TfSw19txXiy76o8wCbam1jH
7dQjhT0axJWIqYwR3n0toJnHUGIZKd/c4XHQpLCG+HLaMy2SehaxPyASHKk+NIQoWgOfY1ZY0aYZ
3q0PyM3aXjtSShqMUNcPHJw2mX5U+k9+AhRaGuQwuij4N1Uf1MsdnNmlR99bwfmzdzgC8LJBHqIy
zlvptmfW3KsUTx0/mUaNcta0/j7aDNEEfgmXGPiWYkst9cf0CFIhb0Jucj1l84qSQfEfXm2zyqiZ
7T5S+qewFlIdK1LwrmRQQzSrigMeiggg+CuR74IFsN49y1WT7fZDUPP9lLOA8qZrQf91X8HQ2VLY
YAS9B+YmWOFgvQ3Y1FcgZOiMUaQgL8wc/a19+9xKT5b95BWuDfEBwrcNMafinCheHnLZCLkAZqdy
Wr8wVbRyqs7P12wSUe7jvv696XS+FsOoGyS0RqL4Rb0qWfZfdl0uIYcBXMAOWqsAtEqhEdrg/z2c
OYpeVT8257uq/DSrKF/h7grRsktkQBgixwUVjqigBrsd8IbU13FLEWwZ/FVJLZzvdywt9B56Ylv9
r3gw7PWFiovIR2mQ5FmLMe7AJtKU344I4YPSFpDg+wAit9E8xjpFBKc5I8uHVJnteH1sSusKGpIL
1ofWPBDSvde5hS44TfHpSeV0Ne5T4YIKYRqKWbgJ6QGj+rz1ClEkh8OPq0djTsgLq9MYQ58lx9AH
Npo9S9X1RTQvblpGjFKOroXYVRM68crNybEWlXkgPumsEtkxDH/dfWkTZDVzUSjU+4T+U/y/ddzC
bT+A7H5Sy58VQueCO8uy+h1pggH64zG0nClLoGqKNVzOJRAW2J7XguaXQXtmmH6e9UmTWV3q+n3V
15NyMshGy3xE1wW5a6a0J8F1OAakVA3bi/tpgX9YeJGUEg8VC2apmRxAyEgdiFdFWEbI4k3K1KOJ
vuo7krYfT9pfWNDXeM1FC1V7Z7HDRy9dTaVI+TOBH8ufwA+hqqKhKItcTQkI/6g9G2DU3L8nUX6i
qQXaCMQuqbuj0nB54Lyg4WaDQ+Ghv9nQqrgwKKtKOBp5eMLElOzHckbnt5FS34IKSI9b8yWerSgC
2u7aGn8e6G/u981KHJCHnVkUw9RF2SZcHrRQ4XaJt7xnt3fkwsXAsUE7IMFZVZVL/pLijmxiAAYW
jY/9MzKTWTNklQIq1EXtPKXrAXIVsG0ZG98anX3Av4X1QP49N/xSk+NZkyUlqlNUQnykx/uRcaw8
kdVZsEZJ47hOqACp4tIXdEWRCzQrGzhwOEHTXyREnoOislA+HCqya2NeLZZN52ss0qGPSA+55WwD
wxmlSLv54kBRF6tbBQaYgYvq6xwdzy0CbkIGUJNm0aEMdF0u4e0PxfazoqXy82LQMtfYOiCdkzhk
Rc0L1jX7GnsMQT41/kbNeqC2PzNFK4J6ahhO0OgyBAvWn4Q0lpPuFs9Ut+G7t7wkXKxZAHOob9KG
9bXYm+LioLP5u6IG9fAKGnTZpKs3XSWgSHFbmxXwv4FlQbQ5utugDqrkyOEvIHUSEdvcrDNSzL5t
a2stST5fiEn5MYvEXW4NisCiZvLWwPgPAa+4qHixmrengkGpkKlazBj352j9YiWQgvb98kyoY0IA
G1G6MHCNs5MkUwIvRaF4KIoOl7xhSBehT+VVRSWuCY5sILcxCE1NdH15Qik/wCRjrii6+Ljx5auW
HPOvwqz+Yx4CKEFgsJ6njJo8/1YsYLbJEsXClgISQBIhbcchwZCY/Y1VIZ9j2u2taB+8iyVgEQta
gd3CYmmjXUx2hdAREFRmFk5hOJbebLIDl7jSKM16SLA0wyVskN9rewOLWoIBiu4JvZfOMjRNAFhR
qoNtLgsx7LA+0/GvKrHU3Syi1PFmGjM86nbyQ1UO749MxHt97qDmmsv1RwyaYlnvhmSkrgytNH6C
X34TlNKsIRjZCL+DyNy7d54kxuWdqVjqYHTiPRyWyGbe+syzlGzp9CgIRbeAtCyfJeoHCQ6E3U7V
vYMxaP7DfIjuh5adpD05suNcda+rBeEPvnfMP4O67om11NzdjbOwO9hv671fOl6qktCzpTQ27kwk
thx+xs249L36Y47JkGapmO5UqS8JF2i4geE409vOcUuNiC4xROwU3Kudd5K59M3zQJFsuYJqxN4F
3kSGeprlmC5y5JB+y70DpAIlLJ+ynP8fDo6qFle1Vl9CmWTLpOpc2wNi3PPkKksJ9udd/vW2CnRt
X+NJBmdBFknumhcLuFfv1HrgoZP02O2kbin//6jOYzMgTi2ouWZ5v4zUnSxIpQ+4ou30P5GkJPG8
2SD5Hwa8VuzjAQmaRRRPYYxdSPkSmY2pjvtDS+PSGn9uXUUvAUF+TLNupliYkPWFujO9UNsGPvLg
2dK7axWWkF9NBCbzhIH6tqvwP9JLVXClBbBYWeVZm/ZpcFyGJauNYyZ6rkqDSjPT6M15BT+x76FY
E0wuihmHFObRBexzahYY3D3tCqkUJkraTFR5eDVstr5mrlSJtUNbxSC2tboUWIEd+1xpc6UNVr5E
17mdVHmTGgpZFG5PWw8anpMEYO5ixyVpCJHC3e3RJ2kYI/wtr4hy4NAGMAnUlaPJj9R9j35gEY0+
Y5nN6BEJfRSHmzu7pDgcCLwcfjatUAbGG5YKTrTb8ClsX78dW69vPFDg7xkoI+PX1VyUmq/J16DD
wHcipsyOYVYGep02oHpZ4y+8/Nr3FLaTWik08Viy+h4oTZurXawAJVtKkzUvd6FTnq6NOsOBQaiO
Ha6OKJb+SNVFOzNstoTfD8+guTb4TQvIPmZN2YO/oPQiptvqXoTPYxiSftAqKQJ0WahEgKM6yJlh
Tn5pc3epZi2z9FDRN+vWEQB5PMOmVryZrUJL5d3tmP88XhLofwU6II7SnF12UJtRwmuVYA/+fxik
thCp9l2D0AuBiFyL5yeRooCdEoLxG14ecpAAQlniERvpMuO4ilPWAM6J30n+B87HXkHKokhGc/Ri
GNM=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K2T8h3dyt9TOZCdO/ps18I4KDBjgOxXK0GTrjjbYwZTLQ9icYs5/hFoWbXODNJdy
Cpgjip0hMWmTDYIpIDuSnh6D1bABHYwcE0atdxhSx4B1Uh7wE3Dn5IwT1nLvd+y5
+2xsk+wiPK9vcBzXO3r3bY1bXXMVQvW2zMGcC0NYLjY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30976)
chkapKJ6ddNQ2Qdh/wqnHFFw6SCgMpdvjPWR0uo3QXY75Wo465OX5K8MGx17qP4N
DbptQCf86T6hIaiMvggc1dAcjNPjJpZVQZGLbklNFCQqN/z0xmm5Sorw5e+MJW5h
vFOIkrOPwKCaJgrmWJhz8vkwtN0ZyB+0aJDQhUlTB+n7ZoLmpJb61C6n8i7Ck7Yo
Ye51Hs74z3lRZm7ZJDvuWTt+zJGz3+sL1LkzATcFHqNPi07tr7Qq14K6TJnteEeE
MtVNtA43PJlWkNmO9kYk28XhsqNnfxfMpinOqDOIZE9zrkP/CS+FxS42IqLlsSDW
aezW3LBoyLx7sdWEvRMlHmI4kaZ3f31CIrf60qffDLrZhenbr0WQnun3QhcTuONh
f6Q7vYOEaCAcLx9WOoBLPzFgfYDMkn4GxSQVrfvjOxjTzdTR3+lO/QlUYDQIEIH7
quEp+lUN1OLLiikw7twuEMYcOyzi7Wb5OcOyQ4nrJi9FjFmQyQKjQWWmj7HNtZrE
KIsJ6ual3SOUWq8qIzXyhj8nz2PMq/K8HwTYxqtak9w9me9e74TZ2PztiS4Qkir4
Bk59Oobtxh5VLu8egPt7peFYYjl4u/5Pp+MhzgULeg5ebreOOfpauX/OIOOuR0yJ
5fmrkxmMOv1KdE2niUQQtYw3vd+wbGXQJbY/EdD4yVPRCq2wh9dR/aMPvqUtC35Z
Lu/TDkMJZ5tfuNZZEWeOUAYv1TEoNdb4Rl62xJoMuGQiWNwmnmYT+7Tc9Gk0o+h+
V5PEPKaB+DqkZ0+mLhqeofJkgru4lWx1xIHSc5QGidNmEgGvB3nxCtgfhy3TnWsJ
BUmMj3wI22eiJE227upSvF9TLy8zwba8ok1INeW3DMgtSX0pvdv+X0RMqHk7sV8v
a554oLFqt92+ssVOt9FmvutPqrRXBSrnb7HkC+IAZWZkwLLu+aZGNZAa5PJWpLAf
xgZv+qOiUebvB293aCaoeTCzjDpBfWaJE4Tw6d4KqSTGv2D+xIXdxj9rJdfKthOB
m9iJhQHWRxLVp44n603RlLZu+xtnwpAT+eJp9+pFgC3u00bKToOgoltOIr064kOd
MjZu1wXqTpFJBD0eGccbTyP2qxAvjolNPeshF+mvrMSNdx5eGpoZNSVrA+tUug/L
4Qe0Z8D3EXCDwiV5p4NzToAqE/IEEXW5xT63zXL99UHg9bUl2b+QoDamW1/FvxAq
rjF8K4Qqs0vNwVwp9bgXxlWu4KVq41L7CdRr92hqaiEAwWCQWmiz/WcLRq9L+Mj1
DTKchHDXwSqa06KaeGAvKirAr84emUNDmBl4U4hBPxYDDhjZxn5IAkX0iEdg8RHD
pksBJ9/s7A0b7pwIoaN/6vw/yhmWRs7m2q/T1+w8cV8OrGSxMWiLsxUflJ4KvqdE
gb/Odb8R9jjrKILW90Ix1rXvGUnjNEO+wwBklHW4yUgmHV0yirJoZVW1MNslkFK1
+YiYjMImRRPlSxOcCbPQFXCcZFTJ4QpWwb9OwODqvQQvALd8hYts3s2xovLH9yt2
vPz6haH10jdd71fnXdCsNhY/43ENrfBPQ8lXRc8+Mfa0lPWn3prtp1VSOXfm3YKj
kOIeaY4a2pUg0hfRh+fF/GkNMYzIMQxNhVdD1IzLDBmhCXXdunmY9T215cFVtGM5
vNeQkCodg+eoaDoG6Wif3bBTcWRl/BytFEdCxpII9RBxq8FABHtMbj/1S0F1Cw5f
c/IQ1TNPbA7C4tPsBuEf/+vETezHJ7Kw8p9ft4pUy8udNUlFh/GdSRdeobWjciBN
z03JgR6lOw2ULqoCthh+cojlU6bM0ENF8yy63MnDATuD00/GAaEmP2A7IoD8XVDs
7ysvrNf6Qzbozo9lViXECyPibsECluRicUQJmLLL4b9hUUKP0OsYYNsxlTP4A3/f
dqRMyrdMVYi3gLgDrMSZy+6SDthpmofGNJK3NqppV/ZbwClHVgMjMtIED8aMURJ+
pKjI3QfTKIsK3S0rtOkGC1kxfvNqJBq3qoaF32yXKwVUwWbLTRbt96n8bJcb5ukV
X8N2Ziw/F275CYaPWmWwzOwJ5TOanm2EIdInjnA5e8bYrCM32pCRV87bz36PCfk6
2dCtRZqop/440cb66Zikm2MD2YiYS2iWua4n6nDTCmhlZc+XTAMote167MtpH1Am
Lz+b3SkA310U467L4os5b01sdkBLrVskMKGvEwHT4LbddJYrzlVyYAGc0YDy0GMp
G4y2qmQbm75DZ+cGnLPvmXu0gAyilPPjluoCz+pt+SvRO2VJOpssSNo9rvgJficw
qmXNDqtuz2yG91mAniCQoQDC5DvBqub4M46z5C0gZSHUPuuiJnrGwZJ/ERofhZZt
JYw6xuJCLD+uGp30ljitNxf/UvVDymFfTSOIqyjwYN62za17Hw2cJjMTA4zHCgAE
TM5M5svB1XJYcOhqhgZPmywaOASGw4rTbhmrZs/qkBx+nAordwxroIT5AIHC5Pnb
IBtJ1bpSR13QkBfccCgsdTixS8Vp/3eIK4xkwzddpiQSdEGLas6y4Mq8mK98RUFa
RnG7Nj+StHtnCf7OTZvBsbgyHLBzZbv5amsgaZMHfLx8hMRZEbC+2XLhkB6Jsv/k
dsgdSWAm7MKXkW/aWGKOt9bm11g/9pg1nzulgH7i76wyu6Jiybh3T6i2InvxIrWM
eV7NLGN5Yi+vI/SSRaxcksn6x45HtLGKKNhcmBl58XAtPJC3jm87wYjL+UFvbgxd
Qcbtf0OX29Tpc5hvZnawKswhx+bu1o3J+rBmb704HyZdrNjiU/wGuSfbvFpaJ9bg
F9ogNA8bPP1nI3fd3buySmRsADhQ19pLD43UxYxx5puOz+RfxZF8nddlw/59V+ok
eLGhDAxzr0bNcFR5b6NPHelbbr8oD7jfpk5Rn+r7ZZ+BCgvoc5B0TDK73tF2JnVA
pjzePnE1Ld3uhZzC0ULdB1zjF5+f0FgK/oW8NJm7tiQgisVvlu7VnUxftdu0Wxbx
Wyw51Twsev4E86uEh9aoHTGXvhSE7n3+25CW/sL9rZWH43Jpk6E+qz2KCfXyNrPE
pyG4EwoovloLwCOwZjzGP47OuHW7HO8dM8au0ieHLqR3dRLujMkejYl2KlVEWbNi
lPUrH3p03IkTpnJOlr4JegIy4G5J7/OfbRR+w68//rimACbbDqj543eRYgiHmcnd
5LZb+wZyF5uESVbJKOBGctezFRfTnqv4uGhb4d2qmDlZZqB+qIsG1OUgwYBgKwAU
hqJhEXDNm39QfitTtx1rKVrSOVnNnxmWPSgPuLs7IQNGKXnDBpA/mgQhHmrUJMT5
c4adPrDj6/3VK1XEb+ZbDb7y0zxnsX/e1lNUVgVjMpC4dscoFfP54Si3um1sZ7Nt
pw7POCSRXILsCfnW1VhsW01ZPdeqrzKuACdYxTox3pldrR5b2QzTSxBRoc6Rnipi
G/m3zbSdWvNr5XU89C4D6SG+Pvk5IWws7/kRb17ZUi3O4/MbDZ3e/61sfeB7bKMN
aNFCF47jHC7Erv1EkaQNsb+Jd9iy0/sCC/Ifk60zaoVSGAjqslovwbSlHWbTTQRX
keiiH6xbe+l9f6UTmvbGa3dH0dRwDtGdrVUY/ZcGazrSKyrTzts0f949d8MXzAGv
7advPGzdk86YrYuY2K0tUFudJ/2F97IFXgYfotGQ2fa7m8CBs4w4eWcPssrvYm3h
8rNASmf9rPcOnnFHz1Cj34W5CrWB1lIlMX7kT+kQcqLaEe0qRErqv9Uav+qbhZD/
rBStBogXxkI+wfZyaKf0XsWldaJjF7PTnjcwewAvs01wjQYe2z5z2jJQTqRQxZ4L
dbNcckT/aDvQqBmEsNJNbpKJyGRI56RDaVHNxfe65m9oTAf0qAQOvltIx37JNSsI
lJpYSS52huwEop++oqV24k+UH3nRbVdbu02gp27ZhYBTUSM3IpEUBzmWxBmR7A+A
hQZWH9yUntCaZyP2zA9qWfu2D2k9PktD9gqPLItrX73i8Yfe+wv49r4lQEhWe/KV
2MPW5OkKnbaTS/8Pc4pgXd5DQHLtgSZbf9bC6ktuO8nrtVh4V9CrTUGHgy06V2xU
j5R/syB7Zu7cHYG4WvetOoazL0JdezIPdxXr3oQcuce8K9WQ6Eu+Jv4f4cGMH4ab
H7HRVhJwC5M37D/8YFCjOw0ltfDEjqfi9EJJhibXTPw80ur3i7r8XEJoTbV4PbNo
ashNJkBPP0hQlQA/tPS1TJifB9f72ceEaBj+NlXyEOP20pgcAxKx/xi9+MxrFK6+
P8dyEUJctxPEG5COmSly+o1edi6IKkzAmKD/OwLC1NYxzhlDi9+CCo/kExtl7yHA
YDdjJ1fAR5FwOmBpwO1nLpM1J3sxouoSIB3lxwNedCRoAD+arrF+cglfJb/L97Hs
B5NYrzEClnnEEfCEKqD1/ySR/dXEBkax+an4i4IB9K8G6PwcQaqY83GlCDLCizQu
jmvUliK4ifKes/rMCk8VpC3ZN5x8AKi6mOt43dPZZ0H54DRAYej5UNexdyIVrpPm
rcgWXCLCLw+9nrnPOUWhdtGsDd1XNlC/RR5nEPhPQB8bzZ9CDfDQQOpqq/dL1wyu
BT7ii6lmGjXbdMU6+U0bhrUMTGI2QROJKacfGPhymc/PZH9HbOmI7wer/OhmIQaz
RWxjyesE00cuDHypKRsPddDySpQQ90sIKfsTwtsDw60nKaIQ+7EuJTgyaj0RIgLF
TQ5Ufg0p+XxDiPPz28aWZmo+JWuSCzdnS1crTt9QCona2O2uNgp5q5wrfdfwzEXp
ZpGvNDLfurETCTHbk+Nwx3G8KQLDPY3xuI/b/csFCwRKW6SgxvqO6ouQx4dzeenK
H7ujQq4U1okZS64wSbj73QfoAujMt3vMGWTRL+VVf5lLxU8TPgrNeqoUsdqP32mf
98rKpTkgjNArwSrxWjyjQSFghaxVrBqNVcG3puAZ/pRBCp/0HJ91znM7HG6sz6SR
E7ZI7cirUNG5r/5Ss1xaT47SBELNWLfH+6SRVC2oqtoyci3Cz29MejCf55n+va4h
yvAi0Cw78muxQsr06HdO0/EaEwD2U1RZhFAt3/C/N6B98tfZuKe+KGqLWolc+x+1
gWZ/w1xRrFcKH5zJfO3zwicUhvhYnZc1l3qdorJy6nH3qXwqdyxEm/RCCOV7PQBq
gv1t3B4o8Mvh36YVJOOgLpImWEn/F846cAWz6yNuE6BUHJFJ7iSNfUKErK43P+G0
9dxaDUZlRrrcgEh1HroutUod+3BJcoglZCfZSHkjx1k+Zl/WSkw82CqpfGK9jnbe
/NfYdXd8ET36eyBzFMHoOj7z1JiYrW9ZNrdF6IHFey1Ygy93rfJUWUsoBJWz8ZnX
YOtz7pFlwNwk9NVFd7O8cnXuQWxIzr8JFQ55YiyZiVduXbvWyHCo5tRT5vt8S283
jude882UfjTi0mW6QbARRZmYXApAAdSkHN+LoXafwo6la0JSxYNaMsNnJ9UAWy83
Dxc3x+xrZaUKfgi847vtdvwFD1sZ8hVABHr9rlP5fmg4SSQUU4pmjh/BC+jYOsm2
6wtJcyT9wPDLszFlmt8VFmGjJqQf5FossLz6k77KjEBZOFt5NxfNQK7PYtwwzp69
DzBp+vCeBk0q5kFgDU9OWGjG1Hd5j8aFUT5WKbrXCsk2Lq1Ju0RDzr4Svi8oCofW
jqcpDgfSGxFXr1YjjB6gbzaKu7ABiblqG+LYyeLKIse9T2f6S2zYZIU3sGfURhYj
yqftVpzJBtEeQzQmrZWxM6ulHK6kIbFY0A60crsp5SdYoGc+uNBfovfKdvmhT4qK
VAjMgnps/CWNmO298VFdq9kaE+SaEh5tMiy0BO3mlmmL9+L2XHnsLTbxtrXfdbTI
gzC/zwffTjFx5921C3f/i6E5pbixVfzAHBM2dc8P4Hth1pZJlOC6Rw9JGkPHXbYy
NmNViMsfmrGBhMrqSIaMzSItNaJMzjUYkE9qLFX0oaZ+s9qQ10G23iTs7rTNou5n
pPRz8mPtPTvd8y7r1Vkdl75l/eS9Y1QGoEJQMl3lTeg7Pvz53ygVCqliEnmkKCqK
4ZFNzDrJQ7zJAJ+TDud5ywZDfquQU4OETgzI68d5dYdLj/lySiSoW3O4sUuSIYVc
KVb3TgyD4q7KhoC4wp+Wbdc5zivlYEVGbH0y9NHU1KeGT+bG3oZzgcoSqhgM6xU2
dlk72v0gGny90+oT37JTA17vh6Lj1JdkBrSAivISuCFlwofkvgmbmftgL/6wrFKx
6wLgxen66PyMt54H1PK03cTaksxO2hngFWJRajqDMq9ccUbYmdetNpmR9RFOqUl2
xcoAto4wSxsmAiZRe8IqJyIA0ERTaBTVuRKKfgSw/BCVdOAl+xfyEuEQCcJ/iz72
tQqfiYxCdHQhutyaouV/G/BSx28mbiwByZKoWD53JZqy9E31ezpAewwqW3L+PIUE
21PfH8HKQViL4LhuMDUe4VGdVnxgsZu37ZH/XJK88e6jAVe+XBjdpY/atisKO1hP
+wooiwz2JXZc+dUBQ7e9wSx97c1Gm98xj7rU6VtAZw3GgbwQIphi0o/lU4CWkbR1
JkKpx8aHrGNdGZIoh00UPDWyYQcx26pX2tAvS113kMfS95RsiodJm08sTEAZALqu
nFpaiUqw7hz3lzvbVByx9828lVteW+GNAtJcUopdMGKFxMg5SA9GHSjvPsdl+Ada
aXOPHHL3OG8XI/PQjGY1OJqF2sZBToXtliXJTfOA5Ej32QhRcm+eWzewrwY+Dh6V
EUTxImFPsJHMOPdDw9WBbbQ75T+MN6aJinmCH7xUpFroIAl6VjEArzc1gQG8Tjji
+MgvK6EbFGgWa180Way76gpTWlva44mmvVV6hFOqXLP0Qp9C1h58PiD9Udb8kLio
RWER+qfQvrVb0Jx8JD+6g4GcKLPck+QKRh8retOfBRFh8ZG/LXi1eiOv5DZLRxyu
DXB/0cBuwjQMlbu4fpsl/aazu25V4Cpb2aAWM3g7liC8JE9weTy7VcayRQEoUI/b
H4jbjSifzPPSKJDJ8TMwsGxTuIwQXUfyUttCp/cAHMOqeb4r9T2RbhSh9AoSNyJJ
kN6GF8Q2Y7n+Oegd5bE/5+XnjVzkoQS3wPJjMyO8IxuT/35y/cuyWAjQQvhZWnbk
pGuayfGHLoCOBA3zn6gvgt8VsPsEnczcAvwhMAZz1WS53voMC2cqtjketnQZEXUv
P+nCFMs9sRKbWi8t+nFkWAvM3CDwUE8d2XhhBiWs03PJhs4qFN07Bbmx75UXGo62
oPfO923ap8AMfwOY211hREeCVA/nvUmif3QUN+pwgBz8F1isf0lau/4LmusP3ULk
GKbqjSpWR0J3xeuJ5PpAv702PKfJdxluuk2odERIR+OzUoyYglYQy45P1AAxOA1c
rLRmAHEVJAxyNYiAP2ZTLVbKOyqbuZZexWR+DHpsTMI+cymT3cT0KAI3WK6q0z92
EFQU2dcnn0A6Vo8Ea/2DP0JHtuQbqHq05kUCQW1mpapKeSzT1HLqyZ0JzeLG/xVy
HBAI7MK2iMboeXunGMgonj3nbYYuTkLZib2W2Pnu121WAYhCdIBcEsGWZ+7Vsk+z
XQzzPbtjUwSdnDKEy/18cOuduxLb+5Uth5kRafRo6Qy4g1N5CxD0ruDECkkqOEgp
hEsxPN/cwkZOe0snsCQzqbpY+EaOjGyzK77FpZ2Y5fqACBLsxTHImP3KjdgppzSl
hQxsdZJlBcjMHqXUPiKNut5bdMu7Wx+a1fCSApoIry/yRE4CksJVhci3674EjfKK
418LHhrpnFcbLz4Vu+1YCIEbteIPzTC60btdI274na5HQA281Y/tXS+tcKbMo1DZ
N04Yfl1lJR9MZfiOggY2AVXBKZi7JfNzid+3SJ/nT5mVvJVpdmwvApC6S06E1UpH
XU0wgi4IriL+ip3t6vKt8akRIaOCts6pfHf7CxtAuGM091Wri5cRIXkEcU8Wb7pH
/z1z8O58/XuHRONyhU1XNrALc76jhnsCcvVEmNFVxR9LV2D4pC/bHpIKMt4d8zQV
4TGJnHk3hjKi6/gFdanA+sW0qp44BD4XAZcEqhk3EteYRnrQ2/AGBUk4GawCI6LJ
uiRT7DW6zZhWw7fKA7nmg4RIx2+CCh/uHxQOKQygqXWKhi6cR6nyh3fydCC51lTO
xei4XTNFeuAbO+wx5NL9oZbuH1nfWGSOEy5hOqAZbXAlO4dVm/0DkqrrjwFwGT+I
S2G/OGwwsCpa71k+yTY5i+RvPxo5n5xT/MD/JPgHF48bb7gSM6dJ4n7wah9W7DWc
s47fj0wkVCRbuI3lbTH+zLh/+rwku+79X2t2HmduO9sp12iUSdFe16iP4aN9mXo2
Cuz8rMpO36/YZzKPPzaIpABSccyQK3IG7HYQE+F0fsqdZWwio+OsrDDUZ5lI/VVL
KiIE+15LZGBFxMxneM4Wk/Edaea5BlWAcKzLGHfm2RVatptREwR6r5YLF05ljy9a
rubRqV5nxPTd3bZbyZyynnUAEhio6EpqWc0p/uuP6FuP9kQywpwKFmfgwLr7Xqvl
meF29oej0Oj+xo7sel209+5nU8b7dpP4W7c6a73VIRU3Qc5IiY5+TB1uKa4k2tHd
Ybyp9m8PFZ+xP21NFexLCg4mJG5mO++L2cZ+VoYngVZ6iUfgoy54xv0nKjnOdeOc
R+NyBtyLJYD/7ucDt62mIxx0wzxDtwGyPhWONwIPi9LprpdEYg5CD7PxfJ56pgQ3
pOVoTg+vmEoAS57mUEd1V2JK7gvF/At1sN6d2Ka3NMFSX6X1WwA2We3gHBEXk794
VhnlIrhNRqSIAmly1XEo05pSM2ziQpwUYD9N/vLSnK/0TyJrMcHSQgtGfHPCP7xm
BYvwo2eOp+rgUYMzMyZqBlIEzykdtt1GQT1iebcPewdw9xD0hbZsulSWcIFkKo6d
bS2AscBgv9LMGOrNX8daWk2t4rNYnKW+JJ4RqZDftfrG5sFJn0CUw6iTAMXJaFwW
8L0bZc7jd5wTCVKLTvIWuIxL69rBEyvAa+GfTZJciqHI5j99uFjPJx557uoSg2JW
NVv1AJb1a9RGiotArmWi748omf4p1hn2vOR7HCj6bWQW7dAqowA4n1TBq9iitUcf
0X1ogCxb/IIqgxc+wr4cah7JrZVK4/6F4PxABRcbS2isa/nE8xk9f23jQ3QUoElq
h6YoqaHYml6aDHJcDTyPPzSVgc9O+KG4bcOLzNH4Fv3DRtpBD6C6o591Bdz64L7d
omN66OLiuD/6cJRJdx0L7NJba4iE7yvs9POHAITGxmKYv6BoggMfh6S82u6bXwWC
S+f+xunpVctTgfN/nPv6kzmc7JivIwpwUJEQUsRslB9TvNr61+DkGFV0IlHru9ig
3C+k1AHtPWqgdyVvyOGvXeH3lujX+SMRtyyB4umO49mGBYIgShla2cqId3q5ZrgM
NA5N3ZHwK/agef+wTx+7IvFI83QaLO1+si5+dqHnYIXnevX/fkkqZTDTRRiPhZ/g
NHMYGZfm+W2NgVO+I21ZBkxW52Wqjaw3jlNJhGtDW/LPeA/O0h1TNoTFtbICTdb/
TSbIjQDZokgdTtYwIJkjKk/yVETG+Q48CmwJM2ZHRDr3AtxAdwJdKU18jkRDNChJ
U/bvJAFyNK7iS/gpZJRxYL5TzVQ7zWXh9PVNlqqYi8eLwT3z8FoLIc/F1u3AiDWl
5JPKi/aOATz9gQK857ED7NGh8YKr8N3sfEpBHj1RGBu3sj6fxmS4ex4N2mLQgIlN
BlMb6o24fTeoE/kUNnXZ/cCDHDjpUunKqrE0GxgeunZe7P0qrFstI5px8KMh0LP2
EnMqjo66B68z1FkzuxDaT1L12RT3fcG+7CtYRbrLJsgwaAuNXQUFkamt2wxZ0DwA
5sBhFO1f4ApLV9i+Aeci/JSx5Uw31LZ5Ett6wBqylPkd3BxdxlyI1RF0oq80otlL
ikyXCP2VaovlrNL3s0bS/dL616PccVXzLp//j4BY22iXnPtX2k1UVVxPcLhUB5Wj
viA4viWnNUJVFHTJ4jaJ6eNk/h02vel9zjy3q9skOzC8qxQTvAaS7FJoru7d3v2d
hFpDdSjofDEbzgUHv6g0LTQFFFMKfGO7lmL52M9AzDJBcAEKVZklyFbb8TXQDTvD
Hp7NTaKp9AOU819e04SjPy3XdtGXZ4YDZKmgC5LNE5Anfz3uHxmaQRj2l4OanPsw
kCtfLeYfeAI81/d1rtz8NILnUO21MqFmOeSl5AHC7bLXrp1MnYFB/w4etfWREsnH
PSEyPWrHM1wXu2geDZp7j4jV19RptRJaKVb8tHq1NK8RBYOuyimv0SnbclBJfewd
DljYBPz+yl5GMgB5JCcToY8le3YVj8X+QoO6m/lnwueJhR0gJBTIdcWFZWKFnuzD
MkUztp2f8A0nmTlu/VtY3gWTY+IMu/cJ9V5f0TBm8N+chEuM217qJY8Sjj8EysaD
e+aUWD3pn/nq8AuVDbG/nRG0mENg3tibfqR4ybmaw3FAsXsG0vTF1ShbAJOEF3H+
AGJXOiVHW7HPpFDM6C6iBH3zfWX/XkHiKYm8dhM5UePx2NzaKJDWqZ5+SVjgA3u5
PSLZiAOR3ax28ELVs0hrC0Mbe0Sh/AsMvhJuWFSI4b4Q1Nm/WZDcYSdBbvu3+SOt
w3I8Yg8UrgbP6V93HxErtGFyVzMNhN1aBsgCTl0Ai7kZfBJKvMRAPh50Zre8jpFi
0bGbkSMIdF9YYYhU6d6Ujw9bqj+JIg9DaE/P3N6Bl1aaUdGsIxgCtqk4L88kuqdn
3yIpTD1kzrGppmWqHCwC92teuLLTwEK7uqHEl5ZMrf/HVXsjhPf5RaKaDDojbGHT
NrkgZ6130hsnHOihdyjT9oabi44+Xj99kercIB3iLhSB1fu+cjplwyh3suqKUa+m
Ase208HQ5aZO53dmMvg1mdnFsSynCgGpnc03AJqfCkv5Xp9pYBhAUOCp9cenxqgd
RvkXun55JKIL8OL4zIqaw+4CiEjxua0mRHuVSEWv63QsbqqIWOH8/JC7b8eF5xF5
8x3z7MBf2URxUZnKnq7fIj5tZ9mMK5g7wW4pgC18R+OwSQGbEWWuIlNGIRzEcx0y
eOzPJjojfQ9fVk2gu6zZvrqXi2mzIqeNsLQVHuEotcspct08w/ikG8ACo4rc3YGH
8NAktgJ+GkeuyRKJgKqGlyHLztuUNgUgPjZOCmHsVf7uIOgaZlP8ZbGPZs80t3uR
nMgFQHacMQP6FzfXIeUP3cqX9wYDdjdwfY6ioP6D+Vs32VAVrzqO8iTYkH5p5y+E
YHubfqWvhyPQjKz13+gdQszoEg4rj1byaJb5NnS08fNSCJMGvSyo8x37lLWViAbm
luhkIRB/JUe1xiAT0Z0NzInll7RT5i1qF0hCkKcQMwsjLuMNC03EM/PKMYSiUmAT
ah1eC1JOFoweiJfTIVE4QAgsGDtyuvIGppseTlAQhupCeVMWnqBeliHy7n9p1uDZ
bXQdNPpi3eWRaZ1/a6J0TZybwqA6U31IM3jStkctTx+5dntJpGdCUXIv832+Sutn
C2DQUCC+PKEYZM05Iia1urWFCCuyx3ngDiOsOeelrykJOv8c6Gf/Q60WbPpKWeFk
OlOBJZCJvqOp1wksZWIveCOt7TlDgv41lp6FPxUn+wDq5ZfrK2nMburceS28WGac
zkH1elg7Or/aqGrwP2HSq+QMUgXmXTvGVmV7Q1BezQUICjrFYN55m+TqnFwybD/5
1i/zHwYYqp/WFC997yG2Zpm3Q+BUMh6fBegQixQDonKBE4eFPQ5icCFSM9ZbK0tz
qCbZDJAXYsM1ZxFqVai236K3kUztvRHk69cEM2yMsyyMYgwEqJWGCnkc7RJoSnLa
9v6lnTmi37uE2BaKp3MuxaSTX3nBLlAKqXcLfL58lh4mrzmmQoEKwF0Y5j8jTy86
o6Adnlp0ygZz72awKPIHxz/VO4DEJiTD2aYhv4zwCXXaaNcRKSl9p5PQxfkGzfZT
Vt3Dy+2YOEoWzXZO1p8yM5UEnPbq9v3mIpop7t+j0GwtXHJ80TJlGQloHDH4Fd5m
AzcXJu27+hQQHc+EDtQ1wW3eofK1dMKXvxPYHB1PczfBalad5pMcP+YEol6usF2m
f5mZGdohFGuUY6X3iaW1azkhoR/MeEI/A/9cY/1z3ve54/D6cjxMOn8M+SudhdpY
NKygz0MC9ORQq+JGwnMOCuJvb2r74fYgCYlKh0hLEQgBFAt+brc4Pjg1Ss1ORysg
vG2t0c13dWk8dVwAJ8noOyP/ZFE602oUaukd5sKlGPes6Bx+Wl11IJc5r3Md5vH0
WdSlE1zpuJsEPlNpzQT1OpAbFUh+zmC1F7F3HTzxGSvvL5RIcmWlQnC5V6H8Qm5v
sKc2/q/7IPfTUCy78P2PRrmlSfQnhEMUnGstkXpTwQZAT82aDQYYkUF/RBZ2NiSC
vQI38aBSWGNzGpYI5uXJcMd4NbZk3ZXHgWyWWl8V0JikrRzhK/cG9aCGhgonNjYq
mKXLm6K/cD84UNB+w6oIVBJPN65Tf2xGC3mY9Ar5qoekSwS1VLIytG1+k3S2DTSC
AZEUazVKKueFXWDcUt7OFlyfdGa5V9vTyGVRjd5Q0WSXPUlJfnLHZBsATJNiUzVf
9yWcMr3GhWu+MCJ9LHjY3w1MA591TKQOorfho43esIrBwRqIq1L7sczY7HZIpvB2
m/pJSyfcBVVhFf/imZvPVm5RnXMVVIHAWpslnwL5aujdotbKP0scLjAHrqTP35EY
8AUZWdmlORqh/TNuP4BEWpDcPDQasXTD08DtQh92bwsZYTal4CflVRf/8eiZA6Wy
ssr9sGxtcheV2ibR+XRnfVavxEhrrKEUrBb9lnLVeOIgoSp+Pu0JDy0eZElpc2Ql
s7Gj5MgsqCFJ12ecFBi441H3hudV/AMOUlWWrkJk9w+lWQjUs16nXY8LDuX0CL6L
U6UXkV6RXizho49rhFpyuOoACuWUzvFlVmxueg+LCV/JIgBjX5i08kEnPMvruVRc
ZucYBw6qsQzFYfc2Pz4QshDz4FVSvzOOSseeq4Aopm0/yGxNAP976/4dSZhccXaC
19ysk7hlQTRLzZgjmVbA1rE2QQD8lbNZCFhorVDUgFn5ejIyEas6Lgc49BvfobZ8
pdL66QoQF4It6eTuoP03QBtW17xouylb3Gx16ED+KcLZTsoiRToYeHAgkDJs8nlK
lBWdABVojiga4V27OKfU+wTcDH/JeSwdsFwKzsgsz9Jy+rVbXNbJScqI62P8j/c5
pA5tBoj94iLbYDl5QcqKpbwFJ3UnmUz29QvsDtUmx3pdi1D3wbwfQoeWv0OsV5mm
tjOQ63WCFnQ42/WSB9QnH9VruokEVjYKMEgIYz1qT8jlfICfVrasfCCMsJGhzJfi
Y/R8ovMA7K2rO16+rQ49g5qs8+cTNgNPd7YLUdoZ1SK0tvgtfXLvfLozZtumjt+F
HQPTJHa92sfEGJdUmJ2VQmaeso1krwB23LiWSyZE4fKIz/eRCLXYEfdrN2zpsUZP
UX/c2zBcUu7kk1zkiY4svV7PCnWnwpdbfE2hhTjbGnxj0yFVgTaCz6n57EcYAYfx
9AcWayeZBctgQTygFyRkx4eoMoaZAClpZNyBOgYnI/tSDcE3MhhYHbCFHHSM2Lxa
0pk3LI0Vu5HRLsSzM6oz62Z+EMUBVnLQcFEPKvxchGyT+yp6+e6g6u3b7ze1wZg5
2q3S0lpSUdITExTnKGxy/cx3hJqjMctzzuEn8eMHd7o0Epel4f1zHGMOyuibNCpT
dTz+aeW3NGRi+TMV7cBXnIDuWoDyLFL66Gwg77m22+E1XV94H9DY36xJ96bcp0Ka
teIjWTCcuJeEzaA5oOXkf6BIWt8dHkIMgXjQze/5t+xFjResNEgGnjn4T7eh5DA/
BMtI1YA4YBDGW6sxB9fwqpo7AXxHM/2gwUt0+OVk2m49hsxQg69RWnP76nLHlEgu
KtebBxQ9+xW7jKz94NRYIIvftEA/eLZa0gTC6tkWyx3rit1YtkxD/BB+wfvkIQ1B
t05cwph5IUChc6P+3v4LqD0XajVj3FHh9s24LKAXOmYFnCbWOR6uuPI6MVQbZXs6
7e69E1vWA4YujpGqs0IH4p+mSOpwsXbH2B68x0cXVZPk9e4xohkgzA5dTudC9sZR
CRr8wWQs3BaDUcW9sMTY3tQxwP1WK4H2dzO0wuFfNfj0jK1DU0ET0iqnAE8xbDx3
5r4jq1bSnDCO77A/faonPO1DNprDmpr+pw8yOgy/C3mILjsVG0dD87r7WU2c6p5S
AiLDT+s0lJhnFu91U6IyvCy9Flss/6o8r+6NCp5YU8snjUNO92SzAXLLAb2WrYeI
Ffp8SIh4HfzrO2JJrLvZ+XGcLri4TGpn/XIMk/AgMTFhDj/hEZycF8uWKjh5tuYV
cVm7GWSpGS+SrQGTiAOwl/gJe8yJ57HNQ/5icc1tSPfQypLUA5S3rM8azyI+tp89
cTLxU12lkqVsDWe2ni141oAMKLIZo+rtOrSSlGi2bi1QC2gAbtRay679yENQCgDL
TVF2QUFc7Kx0FW+fHTLBQndinHuM7sO1r/AR755muuxyDO7n5D8/9eZspIFufUOX
yQkyyhcbkTGz8Znc9b4i1RpsO+aHsVqCkdUEQv+N33wl2PkEIx9a5DAkH6CrGaig
oyR16NeP7jep22By0kEcdocef9OWEAoT0HkCyq6MV9tQ4aVuAObgHG87bU8ntLnA
Stp5b9dwLFcl0GrbD7wPJcgd75zxqhCbiXYulteDPtaYsSGwBLWhUElebyQLXVrP
FZB/lljF2MOGNM/248Dln9JR4fmh0gsSscsc357fPNpSnX6kPG3T1Xjuw+X3sdlm
ErFCujkIVsWU/hiTIxUTjgx5cYmnpQz1wHF+S1cLocBi2K8McoOOw65Ct2MN3a+W
3O1jB4PJXQOMD5ExJDjSA+xhrXEth8GO/gzumpf6JSoxX+rTdp2I9Y/mU10552tw
AVz4oSpTAMYGOhddm2eU6VRFg6LNm77UnzBzihHZZMz2jPE+vWTxUONX+0+fu8XF
6tMoiqerWXYXZr3VNBU4So1fADIvs8YtDVg94cszbal2v1iGnkpzUF+DF8xd4PGZ
4U/IeiM1Va/eUFWKDxefhqj+q/KdPLx93H3Gu5HMbFMS/Uc0AXJ1KbpmzKFKATU7
3Ukb04l8teMTqQC0p3+q9mp/TSC7gooAzr4atcrLeOHwI9eCSSYm4Li2F/CUC8YQ
XFj/ft6K3Xife4ZjsvyFpRq8Ix0A7kS3HuzKelmuuXhIZu9TjXiMdaqBGkb3ftiH
ZNS4/7Fsmz/lj6RqjKazoVhNZ/H8fvJaUnIvIgsqxf0C+DNF4JbSrMtTyR1KNm9a
ekY/s5CH5+2kstGA7DwY8WgOPFqPtFKK/X/OCxEcPC33fpwSCNiVdWCaZYnrCkRi
PvvzxJElSpWlFridSpcipe7Mvboq94sczvTokkOO7v9F8ZqVsGyY+51GVz3CXHza
v2iUKtlpMBZXJtsYYjX5rAP08kieQvTK2dU10AN3a4P6Yd7Qnn+bxajff4X3PWcC
6teOEL7W3gUW3pk7s0m4unWMV2C2K4yz78bqn1hl0mZ8b1IKk2DO7TVWNrtrd2GU
BTLnKa5p3NzEyRqKkhN3hOhKnr2r912syGzHvfYsmGsFY8ol6S7RgvadbqU/94Dh
RPHnsmDI6cNYZHXHAN31RVS+e7uEmWmnpeoAE5I2qeH21hk3+VqoiYKFyZ/Rs6Ab
OoIBhKOeT4tgOryScLjRSbe2vJZ4Upbp30BNwW5iemKmnSo5u9AHPkq3ysIo2ESk
Qt6hcQvMFNoMTDnDIKV1Aqr+8fh/eS3SNV+ippbd9I2EENIRbuCCYGk1q+Al0wAo
tU7y8k99QNdROnLMRg+DheEv5BufteSOuuwXeFymgY8+Uw7U+3rXZQq1FqlBGiv0
y8tv8o41aiicv51CfxPTWMeBzmGFS5IKd9/WlQBBlv3d91RU6XlusqY6RQ/d9YeN
JQXprGyAaOCfYKCgrpFxtYMfBV3iHmMD8b+ECEtm0ucLDFRGvFBrv+MfE2aTtRsZ
Pb26Jh0W3YLq4ZUiBvWe4KUk5Uy2RyqCfa4m6tEjfMQyzLIYM9p8OtQfQXbrRilf
UzIsbuafmhPA7e5M5+jwTG3NM2UJyghDRVQ/U7T8+Fpar0vO44TSv42MjkToeNjY
DXFxwiApHO3BN0DyaIMLxCHkgsSu12HBtFdTrWO9H1u0BMfG4VSfsaxBo9YkHmCC
LUgVuz1NdbT/OjKtuXLLYMSzyAppyk3IV1XGZZeSOQ0QzwmmLYaz2BJUQKdtZSA/
2u4sYUiW3bkicQU4W+1hiN/kvrledG9nvyQSmOIxgYF1vkPfurVX0u/n3CrOZ+Mj
MZAQ8FbPmN3P15E+oOIETqbcpC5VfS5CTqypjAa8q1MDIAzhqve9IfNBmXvaOr8S
RNp80GvwJae3kc6ijdUFbyWN9zNnWtIzmigh4CYKwVNfKtuEXx20YsZ0wAeuEO+U
unnFiYTQbDbdwaN0+/SREnDzMh4S55FGcTNgQL7eWKx/t6UtjAz1l7rv4owMy4H7
I6kcrLV7E7peZMhWp1nqChgyOHAAdyVJreb3F77CQGp+9B6/d5zcGUUfJGlrMoWF
hyWBj+tt9IixWjbcMCyVIe4zQZEhjFuA7abAtZxFKkqWrJn+HDUiAWFgC2EYwulM
LIjPBSfIsUWaQHA7bFMCVSJuhQ632hGE1DLbjCN4vGihjmde7tHip9OJn0EqHi1a
nt4mrc/elJxiV9IlSWRNBGXaqvqCvcFnJWNocfqfnEFpxSxQAqD2B287HIF/Py59
vHdXtdD9MHVBYZr+IydlxJ4y7PIbngfI5pK3IrczMtbUiBPsfpFq2mcB8Yk0ZE7P
TBwKDgmq94Vg+QaMUQ0sBX3patyJu23/XILs/iJBbSzbbcWQNCCGOrgUpr6ow7Hb
j6fJGc/AplTY1YYap1Gjsq89el2np2+JdPn154m3yLB611p3eFTeIucSQ6StwpuC
tR7U8XD1GzipU4sXiuwszE54kxeOx9mYIe9jU1TVvbub8VmwXOHgkgIGwenk12/9
gQi6aY5AKdcm1BslJ/Bi9b7IcjavfW3eNPPBnA4Zbjse5958aalbGCArryABaQst
NbmFE8hIpacTNFvxvoLP2ye3011UhICliH728ov/oFQ/Kq1BoFuE8zXpGFQ9yDU6
5WrBkChONT14mAwhHn/AEqwI1MZR55JkuN+mpOUxyTNGeIsB3Tx8cUFwoyTRFw2Y
WQSAgeorS1GCkopdJPEDPGrXg5QwvPMhxX8p/QjHJX8gwZQ+KMAGCYQgzrWfJtWT
Y7Bx5mH1seKMOKWJNiuz5Ip7Psl9IFsxi4A5rohebgHLBg8lLF85XcBrqW640D2Z
pgTf/pcHB9OUdEO1+DvYLjKYpe7TkdbPmZdrXwpltozZ0CY8ZROjfEsqeqx1Vg/G
Xe9z1k2ONKlrK6FzyzoIRQsOq0dNRcbOoR8r/XYt+tjO+kqUbX5vyDtwsrl1ZdjK
UfoZKK+M6W+82tod4W6YJFIjFJzN878UjLJRkDzQ194cQ47gldVRUVnoTnHJsdC6
19K5x+u3DDtqOIfetmTuiq7VIFcoGYFxKh1E+2CgFSA2VsH6PgnxodnTmxa/ukwf
eoNyv2pybWmLB5CCWmYhsPWE+QwL16crKThwhLWObX0VMdvNdZoDT2Blh2XfPH1p
Qv2K+0Aep1GXu0BkzbhZ/nQwgp/iU7suwZGhExAKHUPa1+aTeyAO62JuFDYnFkl0
b7PHtGYkAIHnSwVuQtFCTDvsupFQItUi1DWCI8hK7VxQ+VW2I1Ot8gic4yHT2OOm
PyGbsnn3TF6gRp4v3UVzwZF1GrRgRh3bQEvAenYS1L9VoFoUTrnAa38eA6+jOGXt
E3gQjV9mKq/M39zbs4p2lG7GqV58J0f6WzzlNIQ6gGebUyPF2/2xDy6TQvgvoCyQ
tBsdZnTg9LiSdKGRxhiuMzjUURkgpJF3WzJQZ+XEtd0LVtCeeDnY5aZsmLxoaXGC
UB9qNZpC+0k8ISLRx7M7K5H3P0bGJD5JxWgQnsL8O6kU3tGr1C1BI+mlk07GGIPv
oyr9VkB+rnbA/aKhiWpQFafVkoIsxZMG0UmjWz06vtinzWk7ZRTyMFStneppX1LC
QpoJsMfPw9l+F34+1CJU72XMENqIXvOj9GZJG5YIRxULZAPTl50awrBG3RInyuRa
ReVcICBguXn4KoBn26lr1k4Tsw0Z5z0GDPVZt5qPOI9u6oC/jblzG8Q9XAKkeeE5
WSvRTeU5gCt/1TYloGV6fyYbzu3z8RpFwyewJevfAy3C60rwbmjy0wQCOxRh1bgP
P+sus/i/ynXqS3QV8155Mfx+nBN6XCSW1eouuvz/gY6ffX1TsqHIBx3WIr7KrEo6
bBdPW1HPhpCaZqhi/thqDz5QDeZ8OTWvidDgPbO8zYotxZl2wMR0K8lWO+E2KHqP
cdp3fNHjUInVX0N8u3kPyqFIzSyLLpcJTWwvvDgK1K2sEngt7514I2zTvqqnJPmZ
XzqUjzYt2Tyjh8cnmbUU0/Ol3bIWiYP1yP1cwPrdvt+Sug3k7s9wWsq0mq5MurYv
8MdJE6UT7A1ZNbIHA9CQnzEUQp9kmLntRTIA0LlrMmT6J6+68oRvLGM4we/A5don
VxiYm/vi4nAZMiq+SUJYEq5BmTH3axfYvEdrs4g/17xSkzK8w0KqgJo04h/UxUFw
Y+zZM3bCia7ednqItZ1kj4AwZ4nOyw4znfeIAI5xsjUq9CPfOaOMtYHcr8crBe0j
v8k3rg8sgXhbiFMRKRrQw5VY74g4DJoIFNoHXWy4IzGZHR5KNEkUBFRy63eV2VqY
a/S2sNkCkVKcPFQM0Otmc+eFjSH03YSOYPbP7xVBwVM+utJHMaugBZbegqyQSPvq
qej8S/+UvEXC1hpYL2kKmmk2uJHqYKcutGfmDBi1B/8kSp0YydW+kKBaJr/5M5qQ
X0qIpCM8u/3nL5KS50MJKeDckdRDXokY5CwC9ZBtdVTQluaG/Td76HwfpxqOGOS3
AL1W8pGP/r/ZkVCI2Cfsdhmt0AAaKBnTbF3vaRDIvf8bbadfJpRoKrh6dpc+HFVr
N4zdvh7PlvRS4qnhhTX0HMqyt95OuvWYCbBoDKg7LW3LSNB+IevTgqedtjnWLQ3Y
/ce5GDTE+n5XNrEEQsfsQW+PNzOOdR4qE9YdhIke/zzz4pYQ5/Ax9MVKNo2HXA+F
Gg0IDxOqtso+MTnJ+c/ZuID/jNPCRZU45m1WItpVwCIFLpd4Tavs3CzXOD2E65du
iV5Y/DWOum57J1PHHk87MJkGibFUhZNm97lLI+YldncQ9Lav+ioZM3jPJHNKfqBU
CC8hH/bTYahwnvWewR+nsgjrohhLfsFzoVP1OnKNdHo0KYwvRcT1iSab1RsPX6cn
Pvms0/7amztXnx5WGx3kz6j186Fl3vmmFDn6KXcnhfxzCTjM9ahFMV1YK4T+zBfR
J+pybqlZd5KxM3C3bntFmu4CzZIm/9uLSISAlIxVq8NQL7EOV7ZNyClaEoBpgUFl
G34NHHSW2vvlWumejinEfHRHVfDcYYQ3+mUtWBSSvgWp56oH4q/I2917znTtaG1X
VTYa3J5l2utx1djfyH4lhIIs9bjnkidFwEWIcR3LVdOyFcaa1qIwkFGSe4FwLZxQ
OJWI98mZxupOqEaQLkTZMZB89ARi/UWhnk8V/8zsMGO08UVz55mqz3/9OpJ3G4L8
DdWodbPXpEOuNysLxwclgoMcT9m9AVcVN0x+UzQncR70GXswco35EdXffqyyRB+C
1h2v34MRNhoJRPBXBR+/7HwanD3CiO6dXbuxeOvKoE0i77TW3nIe8p3FJodYVdYQ
YQOGvr09kR4lMIH70lS+a9Z/JopsPpOg6zwJX77WTpntIYM0ehr/rCM0k7cELBMc
k9vceXYal6XfNn78lZ93OdBoca2juM16yrvFx2ca9MRaHEdZwyKz05czfGhsV7/Y
N2PVv/dUBoc+Er05T1GFuqVrZV1CEP4BlkWvPg3R49yAIsla2CehC2d0ZMEpqYs3
zwf9ZHBj9zDgl6KUaphS2oL13JDpd6fRUxtC58FjO7olA90HW75wtXCw1LMskT8X
I9kG+L01jE9W4QbK5knb2ch88w7Z0nBSsN3G5RYREeRJ8GQMnzN7HEeV3rCFwGF3
S3feXTrcp/4j5slIXuYqv6rtYPYestgI8PQmmKDMh/eYbtVKGrOGy7uU9TpMQ5bs
FIGArKQ8dfMVfjQWgn+4fU92DioAaPizixUOHYrvqqmyyk+CH0VZqiCUcDJK6V1D
cM+9Dp9kV+Aaqp9ccSkIVCXlYULCJeyxPbrBnP2xNKbnUujMGvQnkIPbYELhPqEy
obiKXBRnrE/Zn4G1qmV9JT/uwQD8RfcWkiV6P7Ud79F+5X1sxi4y7g1gUiI8XDgO
3RT9KI3oqLtzhwX+xODWt/8K/fMyzd2lob3FwKhWKeL5qXpOdZVJ0I1NvfsZXgc1
pEqxMCYgr7EJqFnSkM5FILeuja8sIYiSST0yqj3ysDoyrya7zob2ehMrcQvww3GT
/clIgFCqe04cItXrl5nyQ6mjJECH5fpCh4szVeDh6Zy0k42vwgJpXm43VsaNxkjE
nPn8rep4+aJcI6lviCPRT0OByOgP1YDgjsIJlOnCMlZ4muLVrxkomHi5iTs0s7Fo
eRD4FsQ1OG93Y/Pe2OVnS6Uzb3ofZjR+11HcIPJ2z+C0zwhGWms51E82xIhzuTO0
x8OL4++HWiKPYG0Yft1nSiozoLvhsw6CRBlL5U6XjWEklVPfAKw21pxPc06jNX8x
jBYHabtFg+dxpeRIp6LxeLUhQNa5PdYGC6PYZDm+KP65EeRdGGFzSvayPcIb7Oq3
x/zemUbX8giSmFbX7ExIPOPiQaYgN7MTIPv0wEHZ9hqdgggnLE9qSItsnPBCOfqU
TrpR0AHVENQLNTmA7jcrYMtygwYTN0MJoMhqcBKoiBYE1lrs3doYMi7a1uUwn/bB
FRsen+Rl295wu8SNCYRnmkl7/VnLmKXy1FvHJ2yTrowR9hNEc8cFqwbsDvkuuUdj
PFb0r3tNIPs3wG9gsLrOQKUON4nsmTC3Cv4aikClKJVTtMHgxoHppRVJ4lhyBnKt
WCtMmzxbnF3y7VWxWKrwj0b9FgqcsIXrXPaIUaYoFuPweFD+dNM8Nz3l7uDpBcn+
M9aB6lPDpUslA618qVazOkMssO3q2PrC34aytgq8JvyogtejCLo+GCFndImK8kel
tYAXoqkXJg/Fh/a3Thu1843RpiQ5I244N7NcVkb/TS05H+s1YYkj7GkuZ0RRb3Fl
KvHYVU9hAfrgW9qB25GvAE09VeIQSrvtyw9uEF6GoIa/yzAa4hVPyty20MQHWVyn
VDockTjdaNkm9+GY3CQm5zv+nJU+wcR/ZLWEtVM6Gq10bcIQesBliiFBYomJujyS
6xzi+wqsLBVI68AxD5ZKXVhw8QoKAReqZQATEcxfn08RzxwCbAHG0ZhGhNAcvwzW
BTdGSNilMYbvfrvDJshV891kPsbY4Jf2Adsn4qO3YqNOQHWWPdoMXEyjf00xBkId
P3pC5IAuHtO22n16e6KPRy1KJnFZOy4AHjMuSgdlyeM+/sGSKM9l+28YFFtShbv+
CE5Xv5l77F+xbC+bEyA0tQj7x13Acmt7fKaqK2u334ofRbZnmQlLkiexW2wCCzvl
kUO5lbtzZiQUuGkht2eYY7JLMYdLkplmpRZ5CjfAbB6f5fmrPJv0AxkoTfzJ30tm
/hRm8z+6BV18+W/yN43qenCTJaArnGmoMh7nms5Eum5oCtNiaNx4iuX/IyFtLGYU
Wv0WO/FGHkBrhGekltfEHBgqLE+kVbzoDjHCLss4X1GjcA7y0dposkUQYhm0hTPe
4XA9GLPOHv2C4CYh5cc8eStg/M7D6dGioIS/usVnUY75LZ0Zu+CgCHs0rrTMnnqk
eTEXjCBaBmNlmNI9vz4i5fP4gR8F7804ex/o02ZwA1nrAjTK2ds8f8g3a0KMzPk2
JSak/h/QipxHsJs6g/R9WKgkdmuHDlc3zpqbZdJdMnlqstHJagGiTsebUKwiUCCd
RZiVVjPGqElXzadG+fMOKts4NWk19f1CyY/yWSqogE4KvT2Lie9npgMSTpuzqmQ3
FQtlQZf2e/hIlshmEOqaGKD5qMPmxLYz+ZEQw4FiRzBoidXYzSQBM7i1MrHnKq7K
NCjBBJ76YwaVp1yG2Kp5VkHtnhyxK/Mnedb2jAMHxpgtR+B61O1CpB87DVdw5TNF
TcPjqOrh3VG/LkZdDE9tWl4OB0b5Oo/Lp8aSOwcGYKunXTN/CJ8xUyfbp/foN1kx
c2XpiV1s8dsp3W1w3EDi2I4JOeNp8YMUjjSjo6r3P+n51Qx9mcb+jD3FnTDrkTim
hTwKBISEZhW0HwsiqMPDioBjyJcUm+TVW7+34ARwTeC3g4TO9/SL/Vp9mFYUDN1m
wz4XUmxBoeT7y/Uvl54ibU0FQdW3aIvAT7ALP779Ao1xZHAkrYe8yCuI01gfdyn9
2jeW2ISE64Ck04AzEhD15aVeJHhVXmhRs26IW+yH7db74GknaomioYrTM3Mx7gVo
RkfS1Igb8cDlk3KvcG2rMlz85jM3OkJftVSOYD6bTvkteZ3GHQvSsrfrhg4jKNal
CGISphNZqFdbp1dAj38zZ4jmO7VB+UcT6QkoYWis++mQbc0AhLoKRlWsCmU/HOom
jsMtU/gUaQiJxd9BMUw44iifCV5OrVadsfolBtmgvgwVmog+CU7X6IG2KFEJGEhD
v7BFCkPpj9uGAVCJYPEcpdI9obyZvrInABfdXHI5OVoWlU4sUE2QtpoG7sKNf1nP
BsM+jdPMYsk5PecM9PjPUfUpbuQ0PvaWkYQ96BTDe0PaT2urz24G3ZdZUR8YMMJS
ZPBYH46T31sHWRDXlqwbsKxG6jRNcSOWMUSl/VPHbX0pXC5mkQRGfUFJXbUx0IlU
KrLVQ4EqQb/ksYX4gzYEvohPlQCphcBhULGL8tEjsBJEBVycRz/l8qa1o41LKkNl
z7UZgXlZyoOVop3tSkr2H8jHfY2ieoLIOEivGlKHtxzPgtS7u8RSbvYhPSIHTtDO
ZA1QVJ3KQWVNRq2TdhYQ4O7bE5uv0/NYwacm9Il3hkyUFeKUXVUz3w7NmdU1D0Q/
ezeAUlQEWC1qQr7Achnd1sZs9mr106YpDKzsV7PKp5IigppgS9Noxgw5fV0ZEEaU
sUBtRVOVaGwelBAkLwK8taG9/mbV6rytoyse0W3zoboYoHu8bKOpdN6JWhMjvE0T
DiVUHbn5D2LxTBL8csy87dcgOcEwyrShFUo8hP7VMTnNFfPmpOt5EUrLpt+Ge4Er
qsNHvFtkHbkDvW6tkLmhyFHdXWNe2l2u4Nyv4KXiyzJ5fSGPxNedkbMr0rU5a1ts
zfMnsXgqYJ76O4f2qjelFcevznpYSsIlWBjE4FlBQtxPZ42TS+gCxY7dfFuTNPQA
GhXPXNAKwRkY8IS+ChjmzuKoFbeYLGE4AC3owMatfiSh0pRBnGnQvoMR4mcltNBc
0KiT4mqzupG82vuOguis0aIYAerzfIUYWfauulaORI8AQDdANmf6T8ptnhArp9Lh
xjT5gB46eomShFwW+5XR2z2vHV7mM8HDtdg7tXm9q+uoF1C7aKgz3tAVRjujCm32
cFzmjIhnYAbkCBFyGRaGPNQ6K7YG4u0Ux1tsIBt3eMWsN+62KFIf7fvrneXhQ0SA
Bct25qSOcuAaMFLN+qtRTnpNR7dmb0dNmrZbTUVHWtiAsg6+VGcklMaP7hFfQ0bZ
RIlcq+HFAR6sm5mni23gmYvQfUoAcucVfKXUWs3P6DVg7HJHHqYeL1fmcCluPjPG
/6QeBr2qZm7p2HUfbedVD5hPFz/qKwlVDMat0IBiHexO3EkUeBtqKeV/fCYSP+fs
hvtaaIF9kYlFHr+NTPt787MhLtftVPy/a472RdnqZ7c77E/OEn69zkW8EgsZICQm
uU6bDiT7oEFqYQievcMf0Mw0U7YGza/jvwKR/GkKxSSDtsnA/dvBV/GoM05Ywomc
B4DIoaS73hg0k9wK3ZzljRdi7l0GnxQm1ZIurwBPV9k1ep4GjTrDI/FWHBtZp1/b
LJfn4x/uRTvv8fwZ/sG5y1C/uMOsLg+E0uulAPWvqkxMrwVb3n6Wfir1dVEeMafU
EbLqBe+BeGBIyu9DqvHPbNHxzOwoxIhWFwuQLa+Pt2UVjwNstbrU4APd2VShgnE3
OPNBiBjWFLqihopjwUUAKrYMUd/y8fzzeq0F7qhz73M5B2futLF5a2+jlnDBRLXK
Gf21ArdD4uNygQQ+Pfy2qx+CnXdKea4O0mNe+1GrH8R9WpAJ/W4X1TS2lO58uiYY
KMcJ6brfA+EFvdVkgJBubCZhV+4snyK0NJCk1ft5aDTG9AgGTZJqg9Z0xQfUb2vp
fBKqfkCkY/hgiruHonNkukUjakI9s1Kr2rHhHY3H5keir1henH2vs5IeCvIE0/Sd
njF+5clcA2UoTy1+qwxWfQK7wj3/NFAlxjTNbKXYRvmsXsF2jJIW5x/j3frEQ8oi
7zOnhV2PPz35cMODn3Blkljpue4ccfrhoaR3cGrM1zYKfqYdgmIFCPkkfHoeXuZG
+3edhiKAdhyBQEXb55DVm7wydfk4FNodvJHtOgVXMNOcSb5dDUGaqo6nHo8zgwoD
UnMwMhcYE/CcERnF3Ir38ICLK2KUvF2XC1mZjVgjtfy+uq/gZQ/QGEQlIzKyjGl9
CIl6TfsPD5vs3MaZDe9bPharmmmnT3eTfxVP2hb5ehQCEXL2ydx9DImvNtUXBso/
rv9bKzc1vvtROY+I7GG+ufREdSI5W1Ufk5uDVjO1YjpFQM1v9/fuHHB/kymVVO1U
o8xmTa2PlCvDzrP727d7fshEZqfPMPVHvfQktB9Qrfe60dH9JV9vrsutewPqkBQs
W71BKv7205DBzZt2ijhFh9RqCWAOirx06kx97yLj58gVnx12iTf5iPhAe5dGcV4L
tJCNlVdjDdlf3MDPcD/frOI/C4XgJx0lCTbPylbB+LiHrNZN5a/DaQxinvrn1BqO
n2ti0GdDOhpTDVPnuGFc7qjGD9Nszjq2sVmBmzoOnuimW8p5pmOEPT5GXt3rx7rC
7sJ60SSXrDRIworDqRtMZQOKeJO40+kNa1ufGRzu+G/VXPMB1lPJNCorHCd99zL/
gt3ZN2SDJY32OQ4Pt56xYUpSPeiCQZZsLsv6x4fgn+zPJgu465tzls4Odntdsm8p
xmlOBP5V+cl3xRk7y8I+YDrs6wt8WxPQvoGv44TolHGbY6pnowrKNU58+eU3BZPu
qRzjwtDycLTz8f5AnyNgtLnBxUSJl6z/mws67K+CXP0ECIeTbvKcotQA10VXCTVo
xGxNPgFt/jIj3fN7mrt0cl8w4SGkDn3nt+ecgzu4W1k9ArfEVRBhzexwfHWERlQd
8Rf7P3lCA19+vCBbOLGHsjVexu7j5JP5GLu4JDG4axuRRnjo/ZOBJhDD+wfUGsP6
D0eUkLjN/zUJ0rdw7dpgpqA+fg8jB2DnolV1vC2LXeAQ+JzsWjbHPDrxETZPLllv
jte8F/RQVmzuSy3ChWy6ZAfIVyk/lZfWmt4pVn6LLLrT0tu9IqgumcKgRp04Y5Uf
1Hpwn8S7IuxbabL3W6v21awqWzOlrAKDaghgBS0n8I1ydvsJpvlTjzsdfcagewch
pLW4oOwd+6cU8JbVuCzKTu7o8nrWZQGjPHBqSMOA23UYLaeTSZZBFmWua+TsZL+H
pFX+E8qHaDnrmKBX/LrS+9vGHJfKTmVEEe9OzCS9tW7/c6j6EkEUYn84uZCZOQvR
zenTtwpBAlaVv9vMutqCUjLR06dRPX5diEtcOCDMOKcXJggqys2AFAJzR0DLLe6o
Pdo6ApLhRoOiPVRBW62einRZVs7HGaz8Vat3/8qkUg+eeJGLpUwZGnXqlE6Bwep2
eA0x6hw1NmyTLvhIIRo9jRX8tdiZVM3P6Z2ne4BwYfZfDOCD8OsdVbp42BbhZ9z5
AjXjWr/kl/j4fKwv17Zn5WbAF9bWeaFVO9nm2qUZGmvhUzcIAD56OgMQpH3e4FWo
UBvKknMfTsYQKS1gHpOdxH1e3ufz0yS/jvNsDiGtKAN9Xdxmw5xLyQGFgefR8sQM
E7pc8UIEFKC0qBZAZEgS3D5YU4e8IvUjMefNhxcO44N1lIvFAyNE1+YNs9S+MJ30
TbBvRKNXD0RqE/CncQKAw8DDdyk9ek5VihRNQuN3q+lYf3jsgOI0/bi3W2QJ3/Ch
efZugpnczZG2p4ldyn4nkmpqw2HCk3L/HpVVUnj0YBTKyIAGshUPkUUlDu14Reuk
xOPEqSFsQ8K/MIx0tIRAdUQL6Iq8lUfunlg/VNFQ2VbTD/VLg2fLcS95tFKtcTuD
V5bqH9Sf8CWUBnMxRx1PUmgAofvHdOFhSpU72nHgKXJAL3LIHyjpAuUHdzEVcYLF
7H/XiDmvi6KgTU49kT+sWzNGXF6cgnoSaUE3pEcje8C97+08P4oIbdsQ2WIyqV1n
kjeZ7aKLAyt41l75SkrNuo48cvXw5dNulzZSTFD9wr04Wiszy1nkoO8HjxxvE3iJ
nWAa/wSKlEqHjUTw1QltwGqCuI+i4ngSHIWeWMl9bQDF5pyifQT+L3nUy/EVBh56
Jcv1pPyfmXs/NDUTTyDlDiwLbNTBGfKHBecyXidr0OC9IqWvBT/PuszskyqvTTDw
vfvyu4pTuvzsJ24wbv2UR9kVfjxv9X5zQv0qFc71XZD7M8LhBcjYPuI+0thd59Ye
iCD3Qz/8DIMPwrl6J8hc74tKVNNq7aVhkyv7U2ZBdgDI7qz4akcToNbDFsbF2o+o
WJlHLiSTS/K3rvgPTGP8zg05wRxAQxXXwc/d0OkjyqzYm3KmbjJ5jn8ewc9oTe1+
H6ht2g/vSkB9g76GLGc8ZHw37V0anIpmUkokClnPQGgjLcN4wdIWfdiO0ivlQBSJ
Gi8PWwpCU9g6VItqMHprGQQP51f27o0XGwYgTugd7OogkWB5C9tw/jZSy/AC9sl2
BdbYFmfNyohqfnmHGAqJ5KTBwTTIdsN7pDDGkaca1l/UEYsu5XdDUpfuTHoPYBEG
9VQgKOI6FK7aXIdRx9S7w56rIExER2YXDKfnxFaLRTR3zkuLAFpURLlG723Lp05W
AI5EXjqr4+fThKtQ8qmsr7sqk1c1WPmLYBR8QcrSXXoYaIzllwimLuX0btta/p0h
NxTnEQjgFOMwOX9H7y6+PB6LmaQG5kjjtdtMoOC8FLj5WFpQXL0bEm0r/qtuYxhq
18lmIGrGU4kEk5J1FoVU0hbOMu7nuZ6tWGxKJn8c0Bj2+EwKDzZpqzwUW7CUyu13
Jxm2YXVoXSuIycKB0NLppe/9ew0eXAqGKjn5ro+1cleTfAxajo6Lp5Kp+CwnTT8/
G0vYj+3dpOd5x+rGZiUIILbuNp84aIS1kxopus/riUYcRjN0NA2FbY0nStNXSnib
3q7mcAwE3KLVEyHwHjKPoLbiRP43t+ZFS15/yrb+V50Lwj8kF1mNE/2W4cDF1Ces
vcV1ZQDpZ3OFVqHs1yUEjfN+CEKp4lhF1noNLyuuX1EKWrX+1dZmkxCxMXsOSgww
2Yp/PEDzgOG53Af8Exde4QIYQlIcjq8TTAGFEEI1kkoQTxFQTU1K5GzvMomdhlPF
rU+s2ORsV2m4v4OHJTF2eObLW+kAIlbGw79Vk4rjy4zxXUTyKg0O2s9F/lPXfhRa
u7egYAXeoFRgXvuadY8R1gU2auIJC09BuVUzIJMcIYrhOLATuetFabokoqO1LLDz
Zk2pPBayx4fAqq3xPJJaKZ92QKpGnZMvQBF/2d+SQnfcggS6p1cv9/iOFi0T+PGO
5PurwyNP+MIUvfD2frEwlnsStrtuC/MiUpcBLbmrljI0bQGNb3JXsEzRqY3VABqs
ntJxveI4pNjGPrAYBiO82zpEoO4Aj0jsrLeJnrsh1bJ6zZK07mYA6nbsQD7q4OqS
+nDlI3NIT7R+CzAuAcKbaBvZVE3dC/hbXk4xmzWTFij0Om1TjbI/X69WHB+rkKKt
uDEAzBYrJQxfTQg9ksJPDdXllYBkX81HLVw3Lvb5OZMczJy809878wsjOiQVABSa
/BmjwhVBiYqRzsS5fTw5Pv4GewF07R+MvAe880IeArprfMoa+xeLatFrC588Tthn
eeMmmlbcy2tLTcBIBqVMosA+LkzJ/VqM7C6tYNKz6vYfRT2PS9g/RhIPysVy/dsn
V3Qbmsi394ldjNPUl7ZkGjgR1mCm7oJAB182A2K68zzt1fOjaEy+LGz2PdGXPyIY
x1CIXHjASJL7YIR1WxOnN2GlQzghqECWb4MEbk8bT0pK6JxNYRNvmyHcaPIZeKON
Rel12JSgN+bZp85qsXnLJRfrVmukrHt31wccdvSHUclL4We9p3VTCYi5R4hN3FA8
vu2X1Ktlm6sOVgCTXyJRQQIBNX/isv7H7ll5Mwv0qn2ysx7GkiJOPSt4LY+FpVb5
H+wwQ0+fLAaFVJBy48L2cR/fz3co9unUdaOVRK5npj3Qu+1/B79baNLhePyBfet+
yQmZAMEE6nCRDIc5/vJ7HbLz4/k/RoWhV9PZpXtA2fVpuiJQEwo64TKHXJISUKDE
ltlKbDfa3reUwILIxjdpcID8xd+mgM4gNmcTTkAPTPALkuK6OZIFec3WppgJkYy3
kwpSsN2TW+FdW3i/vfpjFeubdMNiPM8aX0kB55LwoadNTw6b1oHOO9icK3N7numJ
1xYY4SCoGJWA9X/XwQ8xvtbjas+HejOofKJo6cj8pqNymAoJqksPCkQ4r9VK8oPB
QtCECIC3qIzoC3ahWVgH3trpTLqVi0xDCEA8YjezoOW1hrsOoe0F4c0c+Hv8A0rm
rZGx4Ec38qQ282AJqB4sURFh/rK6xV+CxOkepTrermpu7u2Zr1Tu9kBaREJ/2+I4
uFpBQgDlB/DiOJEPlZhVjL5DZxsQ06olrIlrGKvqLJEiVTe6Fnv+fQZDHXwCoT9o
jSv6QV05yUnSxE4Ft5TzbBrS7IuAoB414H828lSkNbnGxuqOWC9S3QYRLvegiaIw
5Kt9lMvOLfSrFL9DBP9pwfM2B9w05guMq3nE+4FRHDrciz3bVGXxne77QVOZCL7R
XVjfCSf5s93pjqKBt1jiWyCLfE4kExM82N7G7Pbf5PX/Ife87fY4DgStaX99gUai
23nei3vwJSHq8POLi/wPYHjohM7DSywbfx9X47AlmjQOPNqrUOLQwUA54WWXlMcp
rx/FC6PHxYPuNzBy/g2JjWNAPJBX+F80sKsOg6F72j+mmaaCKdnXXiSy/Hy37sOK
EOF9i8Qu3j7DpWwv90qoysWYByTiUqqgr52llmUa+W8zcOyK5WxYxEMZE323X2R4
KP6SPTqBZkTsVzW5PmGvgaisXz39lsU1AI+h5MWKmQMwyP7KIzyQZnn7WydAEipr
OcrVZ557nwxZvoAB5Z1JB3yKip7YE4tBD14UaISZ1hd8WFylCPoh3l69KOkH9qeW
I8g1ns2i6P+RE7QJ2MxwaRNi8HjK/R7DBg2QC4tuIH5R7H50Vufe+xiKh95/B5Qj
uT2BTK0KrSVaYpJN+9KcTopeG6aYGulORAqBrziOO4n8gbbzVZrKylmGGvr7rNAd
mNaDaU4Hk7z/8QuDHsxegCaRZ2IKe0MfJw0b1HRpAFj1gx+4Ecjax9UramRcZWEu
SGoOSj1tEJGCwJ1uKCGABa4HsFI0GT2FpHH0SaPbVO6ey9fVMgPkrAq4UH+8VlLV
1O4LMpZr1qfgbNwYMz/9di9jxFxxTIvyOivEL8OI/IsDOlG6qSOt3oMo/3oFmx/Q
X0DnQA/fxAzIBKhNXs6wMFI15SxN6wYsTByXg7JBvuVOPnJZZICZBuLO+RZR8hVF
FSYxqOm/pUV/eHyEge4+tQ1ZfRKS8jloh1owDZZRg+a1Ctt+GC39YmrhwTQhgLzB
SMm3SH+ITchZAS8kGyHrAdb7tyKKJB3kNG+N8k4liNUrGQNVxMOj0/uOQYXL4q3G
69Cq6DY8b5MP860rnRPPDQ1BoK5MiNvdZy1lYtNu54oXsBGhRWkwWVVNRmeVP3LG
z/mkv17wqrqADdfKcUgPsdBmfmXltfBr9ZUHxsnw3EJQrf3RgnFok7KWJ7HsZ9cw
lMrxtP04Kiqdf+kDk4glMgz6CTgB6upJUVVT3H6IV/NUx9lm47M3ynid1KrUIfL5
rj6nxR66qNkbqgnjKsS+IlYeIDcUCcp8akQ9wUkJ93l2H2gYt6HE5YjVTbX/DcW3
/KggyvqaTU6F9hkq9LOh1E+CADO9oFS9EeS36UzRUmN3poOkSL4i5Xn1maKrM/cx
ekerQ0wSMuF2Ja+8/elbjB63BT/uOw1/PkXy1mlzIlUf7oePjE5pHoNSu6Pszqov
woYdHyWH9/Hd5wu49hDkM31txTzpWS9HxvdpzIYn2Xwq79Md7CMZqZCJ/1IksKTV
2brEq0z+pS3n9T5NQjd2o8C1lECYXI6AURzYIyXk6mOCVmPo9c93L+7NBXQJYN3K
4nuhoem8vT1GhWoFNLrPJ8xGu/AiseQRAgxTYleFLnEkYuXgyuAQI7wbYMSEon3K
tbvoFns0APDuMnDvVmUothp2QxZaaAi9PoelTKfUPuc/Q/oCrZxtuVbLjsTjgJXN
wNMBonEWNm9Z2C4mGOhCcFknJf3nqE9QvGNkDaTsfLSOX6U/DwRkv0dtsSp/526w
Lz8pvfYMwfoTZDBK6K68lgrde1d9fTy61rmOyjYVFNA9CkbtYm8MRVsqH5Qqf6/Q
D7UkgFLYik3lFbMdMHMzbloejdNyKPjsm5GkCXMlJbPTBpSZvkfgL0d+WiJGzRBW
XcmM2xYUXWEDp9daq1o1BU+83BHAaCgixzYfr+gV3EnbhkgbHxauDupsHyd95JWw
oR7mpzmE1ZLeJJa4N4zcgiXF8rWb6enQVtLIp2LuVr4izyOD5sjGTJWbRxjAE1jI
xFDAXEITuEBtDyFVZlhpS6FlkUN7GIaIe+wLzn3PrlFDlYba9FkHl7He7JHIMtUO
XI0aPSuufMwFMtsDSnlTwgsr9qkXomA/zZN5yOG5Pd4ggikGrS7WUSSoMmy1vgyd
2A5ulyyIlq1OUEy3EVt+7xgbk8vxZj4bktnFvxVF0Q9M6ZLYKwOz1tY4ny912qTq
MufBjs4jgUPtQ27ykO6cKx+0Ygb/ERLUXvsJ8tzWo3CCudCxkJ1vP5sO91q8n1e/
7dHD5QG0a/KAfRNt80kGuUEOx5stmc6QJnCO1GCQYYaBhg/tMHzsM52L4plxni8g
htYrXv3jYnCzNsdvzCyHbsUp5MJmRNgEAldfqe7ak3gtg/XnJ6MPHLg5dUqFVQ94
TkWgU6OEDrJ+oMEKNZjCt6Z33Ay1DHLIc9V1GIfPwLjhHF6iUwXez40AEDq9yfKh
BpkNhVyVnp4RNONZgHa/SKpmErUN1ZXDil5rQWyT/ViBuBrAZv4ABKIo2xnaEpZi
ABjxElvc6tJKpn6KsKFkLN3GIpIdatnRw6eVsGD4iLMjtNXnlgOA//zWNwiYluUU
s3JElqwEZQ3PePFTiRcUdxMW3VmTJAlzEV0pGrN5X1c7k+LqY5PwC8z2JffIp3eJ
0rvJ2syg2jBJUzQ7FJHR383QIgxrh/6ROIgwManBQh3lPNovbLyxeUa+yiNPIu6T
QgCKKtcBHAiqBPwYVH36r4kY2lomJ+aMixqBGFzmp8eVQ45+JUmpo6MnbW+Kir42
IPqAxD4xbfkYJXv6Xsc6uTCPdRWBHugBgoKmS1iS8ugUPF0jphYDZCo3EdH77xk3
mPXexcJroyXa/L14/0iRJUwt6abyojUNw0RXWxVB6uUOSC5Ur3amL8F5x4Rfvblj
nBGN1ZlsurkBG/xa/MYdjSsQCYrXG7Oh/i5PPN+8pr5O2EWKadyg3O7AnIHN9AdY
yikJcREwors0w/FQLHrsJM9bG3T9JpQul4DSPzzvuhJv9XTEIN5SBwO5MaNEnKS5
/hexYLaTJDD/+b5dGvKpzRIq1MdCGl+9tUzjuesbrjK3by4A2PZJsWwrhn4OIKEi
719cCr5RnDi7w76qJUKz8/GbEhdkX5nWGE2HGNDwoWUQryfqmLLJEGqdW7/mprbZ
Pek4Y66Zzv63MuDtUF/051+7N6pXRABtGYJYDzQaVNpwsNcrqlpeZhCd4ujU66xk
k4rhcInvQeEyagVWCu6ZvOUbw834T+gZMIv5MdlVJDVlHdyvV4NqOAn6MoGrPEyd
U67TZQUNzxdZ+mvvF5fGX40C+tpWqTmDCHTHO7k0y208lo53hfcblcyt7qcjHOlW
AVxYJnzIKzHGOcEclRP3Jf1ES93FzHZJxSX2x1B0YksUrJLC6IfjSivfXAI8ltp8
12pYANTFua4sZi7CXBxuOawSE5d0U3Lrtv5dkm1GPQZL1l1ncfwilL4AlSm9mhaI
lHs1X6AEKs80P4duavyA3S0rI0Avw+Vn30tjKwEAiWqlUa5NWiEHEtenK0P9E3u/
gfrngTaHJ/SvXkvxspF+ypc9j5jv0r5Z8zsMtxV4viBfZIkk6LS6IgD0+oXXauAG
BsO2cq2WOB3avyEk3mNcUee63Zxb6kGMLYcenjOUyAW9lCxaUDETM/t06u93L7CA
Zf9ZYSN14geQVkZfoQY52yj0YBiD3FXsDbapprTmfK6Wv/WZlPJI6LQPTnD+r1Qd
yTVa9Q3lVHyHZpUvaIS9A5wVpHTHSIRFP8oeqNVbtFC0749MVNMiw/+NayqoISpS
bQz7kJjvJr9u7ZNg7QDZZKUgskKVdIbsWBbQY8gqgWNTJe5hfWEnM/4dobjgSnEg
d4IJFruO7OkYr92LmmMEMjPcf6SF2azfl6SZc6+syW21D3T1oMaL62GQdP4bkGTB
N181yJbQGNb0uYS6jsiUicafMwFAvDMVgWH8K4MfOMoM/odWlO2cjSBZqlom+jDz
1uoUxXAsBWRhnpGO0JbBkoT1ZojcbT1HTlSa80RsaHHPWEd/kEi8ruINNI5+k2xL
5xg1fAF7S9XZaAuzmJ4bAIeOkJlI/Y46IWUmqrR1EV+Xj1fcpXO1rmNqmtNOuu8O
JYzGWAwyFLG9qVVO49/YDtdCxGcgX5fUyAOLO3ern2nkaxOULyfcH2Jqj5cKIimz
izoQViYWZba8BhhXkrXuSE8SyIL4mMkv3gt+4OX7djam9UfF8m5/DK43LYD7FaOs
hJzWgf9qIq6APcXH5DEFvYsC6j6iUFBsHJZcadzPe3Xv5Am+W73gGbsQBzPPewG4
Xvs+gPNkWUQsPRKqXgSltnt1B/hIhDIc63oIxE+YQh0eKzSWjCSNh/7ok/N0W7rO
5YSSTCGcgNkSNVaZdjC+7DxU26WLFMzMr7lVvhgxowuxi2/yPM8+ujIy7ZWDBxpO
8Sq17jNI2CYrSjpZt6ezSbanSqj5Nl59NiYY3S92w3ctfNxigQbWX8sGbaFmeKRr
tnkTqT/qqDR+jv4E9yP3tbONzyeOsSRPbwChCzXXwdvlOJ5k9+snTcGs2HiFcbql
W/+8w49s2fRNO/CZ70c9rEULW6oRLL5I/8Nsf9DXlWluyYn2SRITV0ddm95It6uy
7RidCTo0hv+03UGegOTt4T5ZphROm+A1COMVYnT+onjBZkSuTsTIZg6QG99TCgK4
HVBkaipwUVnhWHqcbAR/gYYjzXnD+ly4C3BExDeGLePaWslPb6Slg2PUaTPuL3qU
XO1+D9Vyho1fS/B+6BPF+5wY2FWLTr3rPwRyYb4IE6843b41HEM/AymwEVlLiH6U
qhBYxTLilky3CqTaic7jHeqttCn5WXgZBce1KKOb9Uc5XEg0sO/EOU5+rf+laiJI
779m/JgbJ7L0pZ0CiPVx4fL7WO4oHrLuZ09DdZfZEM8xDgtRDh5CJ2OAVj1Q+wma
CbED65IdJZJTIASoBJsuT+ZqPWfHdIlpDOf+hGI+iBHvIMRmjJtHA2PShCr0DSmg
LuVbIopgCU0m6EVeNBlgDwV2kaXDFG+4Ly7E8VRBFb1yDHcMjHj5nCxPdaMC131j
/AJxC/SfAyeoSVjMd89K/T1UlPKHilsBqcGSTFYlxGsofFJSODv02K//8KGKOQBr
/3JFELIDSEVAiIO2ie8fmcIWs+grckCptnI//16OXtk2DxxEHhlGkk+RXgnoil2G
TwTLYBa1TMbntXV5q4xRkE1l/p00gPA162aw5hEyftaoWYhcz5STc/EOVS0jpBLl
sx1cODvbo/BWdQ/ZKmwpfG98n0rOpXaUDXMP+MpEqA/4mxgo36uSFmFSoUpS4raF
THt2zfBYjEhuZyPR0GW1LS9KduMDQHbOGjAQ7D7ozAO/WnyH20k3/ms7V4gnPDXQ
Co8WbaShlw0NZQTTi3Vr2s5d2oMnGksPJy/smZ890dIC0jm1EU+AwfR/Zn18HBZ6
2p8Mn6iiGMHvzmYHvSj7fX0wY5/Duckjtd0mEZqvLpdji9t3Jbek9MsIUu8DX737
c3cjTgbycFaWV5aoRy8g3v4M5W/bu0UiKSwgCByuthzlcToMQqks7HD7o/w96Kd+
cq92jZ+ErO0oXXxtreZQOtl5E3uVI0u9iuU2wHS0gsjQzgko1tr0Qe9gTx1xcoYE
+0kn5TQtL0QDP+qHsoNdlNYBOCOPaqFMv9Sd9cNXDg3diFZFvCvRc1qcPQuclFV7
yGmO6AE19FjgVYZGCbD+fsCkssxcuMzY6N1dmkbtSLeMs471vBjsp2oXRL6+u1u/
SEPG/riUO3kADENxLrrgShQVhTR7qoU5I1UGCygHzDY4UMJFjnl2bOSm3uqTKMzN
laYSSqRY9r5ewUFY91QmaSNLPSoK1jyMh0CVfaK06ydP8h3bgZ4L7bGy5C/SVmCL
IiNvbQxpC97k2XgaqZma20Gx7bHKseuyG7PU4PSabMAzV4cOkRcXyixhWqeDKXaf
zPQGq4ECb7QoY978rFQWvBGyOKA8Tcga5nMvb4FoDdhDMdhSaGyR8Ef3sASD5d6w
dQAZlhqoj0fBd9ZrX2OIsLbsyfafgISgFJoE0qVbWln4BeyW6/GNg7brEzAvQf3N
cXM4AOM9yS65HKX8Sg9pS3u3cA9S4yzC7zXeUD1FdW4HRaqmDShZiH+npZE5VUIy
UEweM5bz1hCzkSgpqbzKvky9lrubcY3+YIZW9e6ehl4rPRZvaQQXxihoZb+0ghKO
vrw+VwyqLaw4M0grLryjXvap/PpoRAoc68y0LciRjv4egyZ7FN+HfFsCy0xaT73U
cR9h35SwTM8dZxzFzpy4teHLWAL6KeWixpAyZJSdxH8Hy9lEx9A5aqrGu4ismb6Q
4/ZTWjb7Fx8UrDoylu9Hn/vrT6w31m+GsTcPPQ43jC5OLJ8UeNLcnfJTIMh8oO1D
D7siVY+/SO1I5JIH679MrUI1tT1hD5hczIjrNw25BykiLMbW636DDnAonpISiCE/
zGqMYWWtu12SH6Q1dagihNTL5pdMZPA+U/JOyNk4IbdPjiQXWHX/koCiIg+KjKb0
agBmqRyLBaveH6bLNSBnFTVd6xygxo9VSSBg5Wdz0w3pwWNo1ubzXB+ZeoPb28xl
2UxRTNFPeEfFkDlwE+S70Mlqg5ln2xwgdnCATy8COsuUVJ6s3AS/yM7ImUZyVhUj
4Z79aVmyG69wq2vh6A3f5JBTItaYSugxAU89g7ODSj1nCX6HVB0h2W/UmQtnRmTj
nVAQabvtCt2ZwA423nKjcfYr/5YptC6F7xG1Is3YBSDdC1sIWqUkLGoR9+3vrFq2
MjbQziwU/SabJSVOSvM2j/7bWq6UFoaZuT39ahnX3mjvlRvViK60XJL7Gq67tZoC
BNQ+wcziwJb86rOPNwUKpSQU6p82DdBn5qpWnpfdYyUfyIkllwyaxV8xfn2yQTpn
3P1Snsf6muo87KiD5xwO72o4SJ3DUzPuHiHxJQiOBdxqfHIGeL8Mirj6UGWvCqqc
5J4Nz+1ALBZE43ZNc6RLNE01kmDn/SU1m/7BDQDN3ZZbACAUq5TpKh4Tw268BodY
E+bY6YH4yNbcXpgM9P8JgCOoHmc3QSH1+Suc33j+LbYV5gFCJMcr6Fzs0kSqOwfq
DNedOvLyCgFiWLM1TsbYq4WzKl0C7xW/R/vOsaeWcmoL40Z6EyPBypctfCFqSF37
8IcE/U0gDIbM2HmrSKXq2mbYPBSi54lO90gT4hfDZ0zdLbwJ89ozhwNo9078K1ju
QSN85mBR+O7G/8t7rd5rTCO82alfTJHhPiZjdX66BvtscpggA+8gO6ghW6NV8XIw
T61Zz5utlLirQlfzOSxysZT6ZtyoDtu4MN1cq843f9S33qbF5XihI//BgiOcwoT2
FGaJZCxhwmrso9Yjx4HP8pYJK1m/+d42uvbMJpsGYS169cKVZFJw04TMd83vj5R5
hTw2nDpN2JuUxy+8Ppts2hn5naab0Ol3NoH44mnAUFPwilj0bjvEw40/ttJfxHjC
wjn2pacUhZedL2uMaAfy77Uw/ShLUXCUlruGzpBO2KG+EbE1NoeSAA2mlr/ZYRDI
I7yrhJ2TK/MhgJXspEedtQA6S/6SSs5qMLLU8tzvXsegS0MlBHuuYU245i/QHbIt
fqpQQLWv7YaJ+E3N80x/fl6K/XoqMicy7anVlXs6fJWLNf0adG8j1Qsqy2he33hI
R/b2tMDrTWc89aMjibFgQrI2kcRLN1htK81Nf1s401G7PSZMrT/Pc4yJEfzPfjsU
hsVUqE5IBpWo2XNqQvtqQzyNtdzOyR9eGEKzvvVIbfJSQoy0J9IbsKmmHbggUOYs
Je5n0pUzl7HqmOR6b/Q7l5e8aZPe4WbQ8N9ZGEswNXvsUBNGTybCHPqo78tQTEBb
eoOg+0wl425pxT9GrIKiFEoyCEM4Vo5fHeHNzWPvzt7HQFqHlLBOHD9CDZ76gNV+
2qvCZQedutO1Drba6vCtsuFDjeeZfi5dv0ushi0qCC4jqUyr78sbGqpeHFF3UI61
LP80STb7d152mL7WLEYllMyPANt8qM7bs5OwzFOcgjWQ9lHa/k6kNUmD4rHVeWs4
26T3KpVrT2fVtbvBhFuBadIaEk4TuSCVi5rC0rs73xEG7oqAOrz/JOEiE6MTGi4l
SK0j+xH0cQHpF/J+ZgcbEukG4UaAWgX9FNRW0cFGrkZ4gVJlzvId2qAX3fAau4YD
Bm+z3841ScN2Ckd9c3xdd4bb6GYYHDqM4sBHphQ9LsQ+yl2CxGfaKxs3JIobTjHG
Rbot2To0jGGWWLdYu+sYWWEjF9tNtzrQGoIpCsgAGYejRr3CXNGdWc5aoPvHSUvG
hvpLz+iGz5WVH5kJe3iEdB6nOpdIkG8y7FR0AfJgvL9+hq7CPvYGjM0QDGkadFof
6Xj5c6MCkRumYX7rhNuCdDkpw70r4xFdakbcvCcjMejvGmdtmpRpFQpbnMvd7Fwj
JoEaI9ZA7OonG3OPaGOkSu9mANgtBkuPagG16rjMZI6NKv6qNovdihkVTS3G5NN7
VQmlzuPdQUbUFItEt6irw3lmVVOBFu8Os4XjUE2R3O/rypHKfFl8xExbscURk899
pggCLUfs/TEkxbWJb+r69ZHOEFpTP5Ph5/uIrIilwfEQkn6zPC8JFIAGdrxQcr3Y
AC6FdbOiRG6O7jJ2vZPyxc79gMtN3Du5lroi0xbrLD//JBUkkIOEcfOMLl4AxoRI
52NZ8DTzVEisCRX6Xg5baTjejmpPG7tlyEmjQIKC/iKnvbHuLOb4oM14vKmvHVjR
4HQ7NYGb8UucRvQUbWujbuOhz7yUG0701LoiOlkriREJ9FeNPLyO9LSUIpbH3Cb4
P2RxI0lHit07A8JH3rW2qc0oTgP1zKdpKOXOKqgXxs0UGzrf8RXkCcpOZfvfzR5P
XrFmTQ2wJWymcwlF33T2Yf7P4HyKEbHZThHoXFnutB2b1gf5XTw4yghZVoTq6umE
na+SPRiPGSK6jQJhVFDVg+X8e8bCZTxn9QjqzvKJCYNOg2RahPKWrvnB38szODQ6
tNCL57rQPOie23QIe/uGVjlcyR4tW0B6O3/lnQ8EFQ11xTkHWzP2Sfx3FR5KbfSM
g4m+N1IA9BejRT1U3ihvRIFWD3Tq4iWr/8TB/9e+0bm/JotnbkZ8+KdK/AFk2pbm
1x43f+aF2nUc8MDnh9B/p9jppMXOyTEtAaixhAs4SnhvVbfZoUqMjV+ZQARE3WKz
pm8wrt2VMUAoWhR7H8WtP3qNhd9mo7HO8HDNuQnJWOkVmgTLSJIuxtZ/yvR3z9Em
TO61JYxdX2MQCjk5LCs3g+v/9Bh1FcB2S/SPS/SGb5kTu0owhA8kVQXqWtcfQtMi
gw2rcHa2ePwEJvjSjxlfvEPhX2mb8NVBr/x3r6QNnaX4y4+pfwKm0/T2szTzmg7m
5XcXO3J5mxUcSI4pmBrPxHBUpJ1X4pUVhqWOQ1a90qT5npWRHg45kLA27yB3N8bn
pWxc7sBE+A50fCl0wrSr9YflPcxXyx8dzXxt495yckxf8/T9G+PNMmKBKEz9yzUL
ijAZuO7ofiKXsmhqLwXyl62oooYlOAQ3sKfkYpItHaQ0g9ngU9eQ8gUrQaFEo4zF
m7HdhDf95xkUxd3E9fSzjtdIigWCShlaCfKEhCCXFdIQ4EDswqVb70NQR3vtm56Q
tBhh2byVjPgnS9TE6WwOfv0MpxmG4VMcQtBGZ3XC6BMfFCDURKNEoiPl3I3rb2Ag
WnBZFvPGaxu9GRfHtQxbDMWeoRbI1BFx03Rkh6h40jWr+ivKmi4OwDUJ0U4wkSc7
UJ9zzw+f9NAuneETuD4DbXwc8+7+mJqOhwgRED+DFsBruuylpAKibJgjxk/94uon
FUnk99eSdIsOyRi4JZxJ7ui39am3iRjGFeFKeEWxcg/vjsybOQu+sGIpkZ4OTa2r
YZtE+2nHJjktq0BUtvP+f7xsfC9q04Ga/LLM+fk+38i3ApIIwfg0hagY91ulPU2+
PQy8s+qSeAt8mmMly90nZa0GOfZkb19JBhWv9s4JM0AhAaSUFG/0hYQp88qzO3u7
YTyLOkYCaquQWVc4+IT99G/CrS+bWDB0fu/523GtMGhmxpqEG8ztPAESHPGieL47
5+AKa9/t7GuHkEQ7EHmyiuapHuIqJJAHp1Ni8XJwqflj8gK7bKpdAXamcEgo7cPz
epABoRdeIiRoJGeKi+kDkvTLGeRVRMwScA11W//oepWq4upn26a/YB3hKxVWAeOm
rLou5ejUm+j3o6hUKKG/tAMxoggDkwwQNyxl9KFRj4RQgPBsIzTPCC44Atj3lMLb
A0yjpGnxKf0U3uGU2yGrwUCWGFaqeSpMEzd2aAVkAfidA/ETXx8aC/XpAOz5Hss0
rwOoytvFsojpiFwFNIkF7IL9L5yclUZY4RYDAqZ41h5N23dt+9GM9KwaQAZNipXe
ld7t1x8gtT0GGcl2Ud05blaSxZzkIcB1Rh+W4vmZfAx10nGQ47ox1enHC14BIyEV
XVDpDW72fTeVFVbW835OFTOuHYwuUIpFgFX9+GyIKhP/0uvA8MPfFESgjf1oWHo8
+TwdS/3LCVgLy4Sc+amGwpVNDbbshxxHGdbvhore8HP+9l/RPv4gtE87nE5Mt3tw
RVAgR7RdglUuQ/4DoXJ/QNN0y4LbEPzBLEdvFjQqSVzqO9m5of3YDhSrxNmwWT3G
xtgwFufAqXidX/dJviuGE6R0IPsZvuxLyovPgCFHpLiynq3V1PvZd/biRt8t/NfH
ocrR/bBrcZL7C6q9amPwDLTpWzcKHAViGwWmWoXbwiArWSf5S57fAeoIAgBd05HO
pGde+gKMz1Ln9ycxS0VbhfX4a+TI+6dKJHLLCiSiwjFqN3a8UKzPlS9c8dGSEfzp
wAmmB/wg4jAd8qBvlnatCft2bnVBLxiG37RTHVZ8MnK49FLh5xWzfR4n6XcVs6Zr
RL4DzkYk8RN0OFcgrJP1ZwVQmc00iSR2vsFtCAwHQ/gA49FYkUyj43KEkKnJ2LpX
Z61HUb1dMZqyCUQ9jWLTgVYuXsL//LCgoznMmZgJ3RqBBg/47hN0IsLupX+ZMNG0
Xxuy/LJtTb4Rpfy4KYTbXCClkH0KE1diZVAgYAhB91/rF4YM2oX7yT+RbqJvBS0f
SEZcSuVESa28fj4H9SQABNrKhQ+ba7WGj3/SVba/JEeuKt7p1D29+0DnPw3+0yd6
29dgQQLt8S0aWiu3jXcBKHMhZERkHLOwKesr+KXyGrWN6ZEJ8v1PwdvRRRgW3xRW
wdkJxMvZj3Ioscp0k42M9cjMbOBpa1XrlxlIQoLqeOjD2nnyEjUwBdlAMfjLPWxv
o7yeaDwOzm2NCh2bZ5CbMQLzo54ScyALd49HDPmYHbEpFJwVz3u9Ee7NQmebztu2
rC5hrqDd73cdvWbIGcKEoc7XWtaYunrRT/1/5wtNPXl+nycitmnfYvA3L4Kqo3SQ
KrlEAk/Q4Up1D1UYSuCvXCYaaO0MIWDbbneiuPYGxJ6OnHeYUL0/quoKdyEzwdrW
u1Fw+rabTBkMCx8jgyEgpmg970QXhKOvF9YuzRVx9ir3UI8XlVO+eHIoINrWUjVh
zBObMErly6Yun3vSxxPf53W0V67uwFKe8QNC69+b6Y9NRJJv2qWjxUxGAVcfFhej
CLecWYXWNkFaQxFmicAycelDN/WGAQIROoLrD7if8wZuTtWyGaavugcwP9CK0t4x
iAWwXc1+j4BNGrY0Nrm+vlu/pynAswHzYBvT2i9rGIvg11zvY7wwAc2VNiYvJQAk
KdYCIFo0wr7WHfuEjhtJXe5SY4TmCI1HPXSmSElo//S1KtIfEonmW5AowqEEDXYg
keCyAERb1XaeP5B2kfesic1nrEdSW/pPngWzsADVUdjSb8h/hVoDJbwkLol1iGJn
0XrAhmT3oChZnP4fKmpAKkNZtjpLzKNsmRng6Vg+DY+660+yP/r2Xv4r5UX6Wmlm
jP/jFCkC0418ZOSeNkwuj/qc0eeOoT1JSojPF9Nm0XAXHoo+W/wXPf513TBfPxNB
rkP3JWOKUoF5MBhEtpUAuR+VmdgwxDrBvWyj3Zj+L+gZYJBw3ay0vPPSftF+BbTv
arZ7qXos9czUNpT48wsJUg==
`pragma protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO���lTWl�0������6'�I�3a�819��,�N���QVQ
Nh���v��PR��3�{g�d�yo���%��U�l��jxрx9O���[faL#����wS��-X�^��)�Y�r�g�ޯ���v��P��`�X;��:Y�Aln���~\�ϳxU�(���A_'�N?��
�_��KG+C�ъq������@��d�#"hy�Hd8����|�fϑ�5NB�l>qX؀�x��K곊1���k�-��̉-��|�z���
M[��gi�@!B���^7�?s�+ԲWwo05
;7v��2�ԋ�Ǎ��EmS��ta���U�^����B�@	A8F៯���_�F��ui�+��Θ������C���y��>�A%l�Ԑ���@�v`nv���=���R��f���+'��ؐX9ڑ���dL3��P7f8<�!�'�!w�L�Vs~��OL]�K "�BG���L�"= �j	q��w��y��e�����"a�� �9K��ҫ<�,I���%Ů�́�֢	!���D.��#R�{�,��D��t�]x� �&�_��@���v�y߃�����m�<�d�vh���� ��w��~�5�h�U��1�̏˔�z�@����x�#��>uEhq��Cz��蕶���6��Qi����Q����t2�Źh����P����zM=dPQ�DP��W�)����X������8E3�xP��NZ��l�O��Xa|)������)�^,�v��U��Ĉ�;��*�f��E �{5�B�����'--�ư�l�[��ŵ\�\�V<�}�'q�sgeÝ�����n�;��n5���	��tn+@W��6d�Rp���ҹݘ؝����݉��!���v�ҏ?M�����?(����d[����Pun���_�aǩApAc��������l�������Q\71Rú��1/�#սE���d<�f��űV��,L6�H���+9x�i� B �H}���n����A�A%��<�X���V34ËI���ŏB��d~
ě�, ز������Lu�4u�u��b�����VSI)�H	�Kʃ��SW2�h��T_*Q���-Ό��)�#9b�;�(؜ur�׍�	�� }�>v�F8�ޢgzB�Z�~��z3F��o�
����zƛ���wЋe���������D�]�SE�K�	ȉ�5� EL�Q_R��&-���5�{x�yKI����Y"0�*��/��xQ��H�F�[h�J �Ic����ܹ*�Ws��>y���F�b�Q�O�n�P�@wڸ��}!&��"
���@ׅ�`�o�����y��� ���y�ܑW4��Jg+M���k�45,��Ui��'	d=�)q�G[a�J��v>R��_�5Bv��;D��M��a*�
$n�o}]��9"�����BL1���e���<���V�w��8g<�᭥����U%OdN$�������nU�w�ׯ��
h&���xh�u�3av{9�<�p���:�� }����NoeV�v�_��ebYB�vñ˞�Ns(���<�:;s$�N��< ꢊ`���\�`	��%��t�������Y2@��0���R��+�����8��F{K�e�<����ˏ��Bl ѯo5��.��D��B��*vv��mV�BsD{mg�B�*�'���BO�@�����/8���`�3H��"�M� `�:�m�t�"_�m���Pj9�M����H����$��%�����а4�!k]J���}x�u.�� �s��o"������胫��:	�t*W[�ƍ<
�ST,�$� ulٌ|d���iӦ�".�j�G�����/U>N�ts|��w�,I����0i��T���V�E�җ1�{j�S��1�bh�9�1U;��f��\�'c@�I)܎�+�
/y��)�i�?�˹I��I�ܓ^��!-֫���w�h9�S�d���[�=z��A��F�Ꙧ9ǋ�6 � f=`����w��/��<YХm����	���7�ݕ��˗�.�ۖ�_���C��x�b��V��ϓ�7����3^�)ft^����F��,_���h�)�:��r��9�o�5�%f�s8�56?�q�� zC��o���8!���5]��RVc��Sibe9��U&������w��|~�)4(��h�
=2Οym��<2�$�9�"��X0Is��<+\�|p�3���Cg��~g�_F��=tzۈ�! ���1�߂�ൖ�&J�/�n��ct��<x��L�دؑ�gd���E@z����q�O����G�O3��6���`��@�Ѧ�#%�7���9SM|x�#�~&�F�!A/?Wr� ��`��>V��>�Eq�n�Z\���&�J����_g�u:p��ySՔ�}/���t�4�`�߃}�
���M�ԟl�$�Ϙ{�I��R������� K|4B�%BI�q����J��]�r$��
k�&�� c��3$�[i_2�_c�қ���X
// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:36 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oQm0/zeWa0LCSdgHAW71rPu7lzkqxWK3js4E5I8Zt/f5lJ/zNp3uwnkMk4bb1MXg
S/2L13ZStMHrZN2eRzgyh9eo+wXjQC/+RhAVd8IjbEyBFJ6KAyesHlj7TNT1qvHU
u2T7GhBzSrysK49CC6AFLtJW3y7JlLWGL9HWW/OQJpU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9808)
vmcsTG+PuJkWoxUq37ZsbzRqzOpWXEpgi7ozhkbtSHzTiCIzyNsGp6iAdqtIzyk8
ZS0KhzMjfVkWE4GuZ6fAdYDddVIUIoyyEzPkxXunb/E0HDlB8QheRA5GBWWhKoY2
2uAGrM7XXgCljd5E4Px9Tcl5pQqqpzb/mimhJAaGHBouv65zz7oxH+XXQguvdb0/
OdOEJDbxKUvDGqdTsU9S9XXI8zNI8LitvBxU7VZKt63WxmtrtgwmLglERWvP/yuU
Pcs1t51FNuKAu8embDw1xcbZTiyqRQnJxnvCfVRwig2rOli/nQ5JaMVJsJFySAmJ
QLr0pZLExGkRXCOYrLJlW3dcyQPa5gWvBQDRBV+EvagQ0Ts5qpQAO4XVy+qDMUlK
ruv2E1o5+RxlepkHOipJFurnJu9BJPqlkbDSGYokIvctwkqVoZq+Azx6B/xcjOFw
BWEyVwm3RlJxWBW8TJzYV9NNwzKlDEIgCXBPjSggMc3MPea6szP3EiluijPBNbz5
DFpYNtTuW1YQ8Jl67AAZpyuXq4piu9Z3mj7+45s6Px8WO87NiBY9yGnD3g1FP7lz
nFmYVnlMtnV2zQGq1VoV7Txa/g8hnJxXgxJTlW/jB/pAVQIG+o+Ov80lJEtsEzzQ
Y3dUFIHgZSS/zwNPPESfs3XuvIvjKW+06WzC2uJmR8dmxMSinA01PBckEtz0Lq5J
dCM5pJZAELbLvY+jQ9q2CJlAzKkFzbDIs9wlT4oVvBl4LipAVgmpYt9jTDwaoFqr
KpShKR74u8QfFdkd7/c2tl/D8isY17O2a0czLLGVTJ8gHXko+oojRcalm4lWRKug
ICEnIHl9Um9CWkSTaQVZNN6oDVOaEFUYVAzOh4UTai6S5dIzQLSKMYb9A+p9ld3P
y8ntLK+KHW4OyKO2vJQjvfRAUwfO8MXgpH93W9Fm4hvNp8tBKzZ7btPQ5f7QXqjR
UTsDXzV3kvaXEkcJ0+zm9HOEfaUlaX7f1OKc7nAqEeoddfi0+2e2F5ZGh/r9qWRW
OvjeEWQZf+pRXOU+Z0fuqXEpQ2YjOz7CnC7b7dIcCj6uLp/fpAx46HCK6c/V/Xh/
ZHNwzxSpLCFoeqZtBvbQRlM3K5YSh42XHbi9Nf2tdoggIzyYgUJEHay9H2F3e/Ad
neJEBE/u/cY07h1LfnADPMbLpZucr1ALE25ZLXT3VmfJji+HHIWxAEZFfuEuOok2
/Q6LE1lpgrj06e9Zdl/+35bUjKXLOR8fsQMAzuTtnrasQlCYdm+g5XJk/p+Dg8MV
LSyAXaFlGyK1eDd2wtTRPu61XB8+oAu2t4x2QyZfGXwuhofOPEih3nQMJ3psy+Eg
6/4+FLD/s+Ld2D5cTVzHYwfrCRV06lSqPqcCtmMtIc+igitHHzkW6Ofabub8+qvY
n9X5xstOQmbeLguqE8iiZkxrw1g0xwXP3lGW+pnxDoLr5v5Fho03P/wxY9KTnBcj
xNCaxHEV91Hnjvl7IN7UIQZ9murT7uidQUJc6EVT/EFji0Ply26E1qKRdlKNg/id
s1nzYD1K6IULAGXXzZMQllxJUHibqgcsVjTnlAQ5Mtzy7GA03qqfdXY75tEFgYi4
h7k6aiRxCpK6Vb2ZD88GzyOKyc8szAkBaUTm+TQj7EkWvpnJcW5Cnj849FG1MVeS
cLLUWdcoZtqQZZqvzCdNZJqI3Vcde0j7XsantnReeDyU6916KTOJ66exiEpFe4/u
55FKmC/it3O1Dql4pWRUTVM/1/yWlSgPQghAAxI7uWGZjyGgIKa0MU8vrsN06Jth
fGi85IEQWNtI526BN3dv64TCdlK2ubXaJNJaBkNAwRu7QSVLYnZa9Rpu0Wi0S8OP
mgIoAuFZ5l0jaT1XRqj08A4QQqY5QA9azsGRp+cs3gfyE3WB/OB/vCZN903sILKP
unJYU8bQyzrQsvxoxPxgKLlKQ59SUB3dS2xHe1FoA0fgEuGq4mnSrIZStbIe454Q
5y5hIdFcIIK1SlbVJtVRfKIHQwyTYWsO4R2oRggdgeAY8SeFIgeRu+hmEVoLX65+
re6FYgThmBPQLVdO6h0nq6kZZMQRxcGVKAfLzSzkkuZ3b9lqCOx9pqgLYwuhE8PA
ukYyhu0ImT0v9oSgGC/hzCWMUiHZgDEJ9xX5tq5SgaEUIL/tFjpTsSaT/y3TUNEm
3HqQTP26ZvTG+ybiP+MVG9ovpMSTLcFoChIJtBneM6DHXTCokGVPQ1BXa46O5Y7Q
kI/8lp5SZNnI+LUwa6d++nAphE13RTsPeyh6URTa7pL3xM02iO3N1pXdcaqWEexT
0BTqUKu7KYNXEcSYQsEUSbfB6sgymV2Wnsa8f18wQ0vK+NOaNELk0jzSsPRyDk9/
/w1jakDlYJzhLURaDf0e+aa5vz2L8nnX3NbR1SrL9Tribr1/JMgU7ZpRgjWjkE0E
lBqipyIjpKLjmNOF5Egy+96iHWX5Cf8zLfT24TPE9aT5iQEqFRi/kkrLYSzB89bO
qu1fFP1fClUN0CToGaP8o2H2u6HXjmro1t7j8SnYL5ykQP4F2qTFPsvQWzaQXXTH
HIa+ndHLxIVMlgmoQhhocH/y6jTAoLJrTbh+4elA+mzKCiL+ob2RNl7goIqEij2z
nTHmbaCxnl6KKVylbepFyUenapYdiCk0GfFQqXrXD5AOvyO8JQ1aJRUQfUGr4IUd
kF605gNuECgVG50bW9gPK59M94I/fz3NEs1qT5oKoHhfSC05htMTRIxQRTC6I8ys
Vyx0GIBqsJvZrZsOJqWlM79USZUq3+U5IbtTHWVmvqgLQAjBe0+TY4tvKEJFzSvP
MI/UxkUVIHCtS9snHv9Y5LErLBZdr2b2bH524xjvxg8lP/udBCwXy3HHWseVA3p0
doh4E/Ai6+itEo23Cd7XbXJDSySV5oAXbnhSDy2kkGF4SAsVXHL3DwfwXMatACnD
/hHHkgsQ8E7zjAThuDC1YOo6m9MRgWaSWTnZUzV9bEoHTz/hcjb1Yo0bmM2SlLM4
uzj88hkn9S2Coro6eHNEoovhVr0FjLDV8tkCFZI9M/cUZH51+jH6gAdzCqldk67n
iWsqdaJEzjnHT3r5jFwyp0iTpo+GvNVrVLY0w1D3zh11dg0PM9zgXfCktTi6z1p5
FIo8FWz92GFTANPv4yljhfSA+om311nrF64w4IU6Sr156fyeevKk/N7wZGlyzQro
Vgw7ljxw2qmrW46nLqV9KyTZ4/a0NhALyMMFSB7UIB5vlCiTYtv38YbL2jdkSk2+
1HCdJBzKVSu1N85iojH4SL+pdeOS8xaHV5otbteXCtoWzYp8CEQlKfQWgtgsPATG
pqPrgBZgRK4TmuqzOzu+hcELtzOtfEAybsJtHoAyJdfrcqLW1rrEqkB+TLsCIsRs
lap8/MMbtyUx53lgMQSxOpQrr3bnLquAwCgafX+V3TNY+3SaQfOZLNj9a+HwgNzS
F6P6vi8266W9CWUNRCsJIqIOAwVKe8/TGB49ysOP+xvfRzL+avFSiC1kRb1ydA7q
Y6CouWMHQZmZUP44dpBviLc1i3FIYiZWc1rSR1KksKxeRZko8nC2+kdtxKpHN7U0
2XKDCfkIcgwVWVo6EnE6d1uAMc2nfR8yzqPyVbnsdOD2g8gdwITuVCLHYDpT5v+H
XUBLXhy9CHQ4TMtAGAKJoFtC08gT9b5SCxI/8pgm/JkwPY2v8amcDV4BQqXwLf6E
sWWgH/uqXO/1Kz2dUB6WqRVTiR2KYkbL44WL6kracnQA8UT5eAlk46f9Rb2y7taK
1IhBoOiQS18lH7G3AbqkkJLAJIAxV4l+bRq70UY6/0iROBvH5aRzsjfWKwmeBmvh
fOgaqUXzide4lmLNZFLB+tRGddMJfnglIKmoKOETQurczmiA6n5nTUM7A9liftgE
NxQppRjGpGq4uoJTlf4NUndxLzq8tK/dMvJU2wdCT9YBpyuPgQ1t6IbvxUJ+FyrH
3q3Or4N99broQCK6FPviBzlwnj17tNcYVvS19NGw0QmZuvPyBtjHj2ZaCfL01mad
+x4tyGHcIwYdH5GWPuXKFL3IDFHNcboeVAufavcJsYfqntbq6R2aHUCxZtwF5JNX
KylPtnva3ZkPjzVqFCENNqA1PHwOBsw4eW1wFfBaPrC9lOEvpduuGSSQYza58Ddy
tLqlCNUZE0srwgCUbuZXeEtvRpQonuWKTPv1aLBvop3oYv7h8zB+LPq9H3OXo5OY
n6AYlIyYbvZf8KSmVaFs0ytB1p/2DCeIoYRgNSmkciOOFdDoezwkpMXevisX/giK
+BTzJtZpHJCKAkK/90TLQXx49Elcc6g2l9afnSXe9ysjOqg9RO++La0u4I8wafhx
Falg7SmBRdr5HTNPT4Dk7f5X3vlQs5idA8zpmkkPOm55k6XmABEMMSwgnt2J6wRC
5wAjHSRgI5qW06AHBvv5nV1Gug38MN2fedwG+ZBskObdbyUF5vI9sYMpI5foY0wp
D1Xor+sblbOjrIILhoc0+94wpdW2bYh/DCiJeFTo4Mg8BYaQB6i55ADWxswliPss
eyNVZ7WhZ8N6VsTvglE+kHHHA8ncCMSe8w+mqFBc5lUpC3+UYP1Zrukh4m6QVF49
mM2GxSiYsFeA5LgjAZpR6UtE9Y6gJmYHUAvU8bdsu0P0g1BLJqhbGKDIuKJUASmw
uRVyTkjQlReRd0FKGBJ7ac69Y7Umz9E0VronbewTrBY6ULBl8qDxv2IMyySMUwX9
s0toOcUv3wjgfpzPsihHcd5dLM5itZu6ugCtWZcksR8fh+1egTP+yPEcFtw0+3Rq
KgjlfaL28ntD57eEVs/0X2xuvmYldHC4itR9QtbAE4AhISgJXdnym3bRdZqcpmiv
1wHjj1OxTuFIiXYWHCyqSt2v9CbSQxz1eOsSi83iH0fGqupa8XzvRCk2rjwyUPFf
+v91vn+tYFiXkbRRcFXh8f9tEVq+bqdPFlm8qJEJpVjaQV0TomHclYdgMHfz82up
LsGUs+THeQyT7U18zRqQz1eTMLzZpesLhcGrxDj4sGwDGz1nCy79UyKDyzoUvoqa
HqAs72thGBAQFQSl0ff+QcIXjMIgBfsZkJ1o5rVAek3Avo8RowIVtoyto9mamHJH
gs4Vk1Q2jpKl2yT/H+Kw+kAxs1ditOR/D0D/mcJgKyqJsq6/LwtY9DC3Xqyyz5SA
lmjY8kD7807blgOUzy5wQrDT9JOnAx5UwehC0OKK3qWuG7HnIqJuUOVFl+VozOjF
yIfSvRa4vM7M8qBgM7jMh5Ie1eUoiq8u42wuWMfY3/njv1Nj+OBW0arEm9+dZNhJ
21yiOWJme3kOsx7cn2TM8xY9e1go31q+D684+ROG09yHUIkfoEbSJ6nvAlCKAxf3
2MIjZz/IKOY6T6Fl2BavOo3lOYVSEPQtEite8foB5/1AsEQRF6WTZvrh8b/PwZPE
0XXBIUhXFcxOpI9lFxGLNbmwK8Ow0fJQiEvZXKg0N9XwqPRBWePgwxsTejqFMYvs
ZSFdtN8lbrNhZomR/Us5Do3ZqjNvImNXUruQhFCeC5TkxOdb3Jx4mEOdhITzZQM9
S2S8WVtqgEJuPKvq31eRjMiolwQAT6HnIZvZ2alXZgaGWi1Xktl8Ea9a49iK07rr
S2hQs32dbPuSDiWOhoiklXcCWhjA9bHT6CyzqFYu/aONzYnftL4PgUAdqKtm1oSa
x2h8W9++ITk/klThav4dA5ITeuqNHkupcX3pNOP6U/x0N1PGmASHEkA89z/ufHrh
QDpJnU9dMpYbQXJiBMZWqtOaR/Nmm6KTbpJqpA7e2VAWyGKOtBvKbnRLGW0Yz6kg
t+nLlPJ1vX8cbzZWH8l9eCw0NYBffAl3uZPC/wOiDThbCYpPBV44wS9LFdmhG/t9
jd2QggcRLsTidRwz1UMDdm2XWE/q00uzw4Qc6lTcp5kRo56rBqKRdB10ZJet97KE
Hal3TpHjdhtmfM1wA45ShCWuvixcqJk2HypTaVickiclpi5SxODsnov/dyQbzR2M
UO3928D/s5aZkBGsRj2nBMdmWmmaQmR7lXNx8v2csoziUKICZ/TGEyQV1ipBcaSI
x4MMBBhyxiqTcxayKhBSItZsSiv+/QEzBEIttWx45Fu76JOUNqun+xpji+ky8FF3
RtsvzaNMLBWr8nmn6hhCEeG/sAlW8SlFDkv/QR7Akjl17yI9jOKcGMESRhMUPLPd
1iuq/3fiMYJNTmm4ICkeKV1OY/s+3vb78sh49jZqSNqDN2qN04fDvyQNJ9Q8oHKf
DabOcTe4AyOoYMf1XE/HtpVPgK5onGnI6faouEZbnmtsdry7dGTsvUQevhH2AaDh
CVkOOigvtU6jIC2zIQCR/3mNccmCdHmeWCZSZdF+G7xyIT1ySHx1klSlqcui2xQb
QDHgV9G+pKlDwJ8uI/r8f7eK5h7Df49dnozba3P0S7+w+lUdQDqkMvtFZm4DIBWV
zRq7vO+n0TqV6aKlkkSKLBb5ulC1m5GjTclpLI1koKbpkFHnZBZPTTmK50iYDzb9
hQ9z0OejtJ45ztLjkiZCIIbSVKaxTBIp+gKTjKazufGdQiPcEVbD6nIijQ1m729Q
9qUWKYevPCxDwaV99SD0PL35Jz6IGmRj2yhOLcCH8lQSHHyZXeC8I3/+fWjIBK9r
aofSJyCGp/UmP0pGgKpYM97RR1IHdjulIa6FWisa2WaEac/WWffyig3Z5CWEeG4y
/0/4zcAzIsLO4h3o13dxNJ8KHNN5njv/iHphdoZCokI1iBjJlAGuVHdGETmsujKt
vHX2OnwysMmeN+8X6sZFce8lwlfAKmDbMK08kFBS4l00H4qflnAAyXcCsJyu+PdS
dxk9hvTw0E/TgZg1NSKUSDK+j44nvnMh5JlqEv4yf5s8EqEzp59ukqPlw5wu/aXL
dRZUTi1/CMPKhW1P24kOO766NYpNUAajxZF28fbSa9icKniud6rOjXhuVJvxGMjs
kOjU0fvy/u3tjRF7U3RJLaAn/o0baEyMk0/8Oj8t7zxn+1qlD4WF1a0NOw1n+2Lg
Q4W4AMpWA2JwrdVJavRtrxEBD62PyENO+fcEcj625LcJy/VFvr2TlwI+Uf1ImmyU
haVp6u0ULmcG9K1mUAEbC1+PwZ8r5gX4Q/PBoV6Y1ZEQPwTLedcd3SbqG76SzxzG
TP5hXj/jGNeOeSsOHtRP8RzoniqLHwswu6bVfRLoaEu9SygCSzhHSPBxR+PMHCiA
U8uRqebPjFNHZaGcXtQC7nTNEYlFX/YZ888ZAE2p1AQCHHadTt1qxm7QjJkcKOUB
u6M0jGirs07VcnlezMd7B7qtK2/pHQ8/w85PWgb637RovtT2XmT4V5dvoqB0fZQ4
ZO5CbxMOAvMoRCHhcN37PG6ffUiUfEK2Usql3mU1/049Cy2+xE2BG5loKDHGDzWg
KS9KUdgBDvYAqciLxarkhWxdFdl9jrxCSQJ8ykR/yC85NsA16iexkFlk1o+nH1n5
sU2+hRW04VKMEfWvEFnJDTMqVo5LKIYonMhqBwYBW/BColSEpqL8J7yt/Fwp5kuR
bpAXtXcH5IwvCrhsYRFUPJcOnQlx8Cu27x2fMw2D4MaUW3w8VwlEV5WyADJy0/MA
kubB3NBAt4xUJoOAdwXlYCkb1oA5uLCXKqGPKJlCKfwNF/fVISR+BiU9qHmtCqgQ
Bxw7ylLQEVO2xELT1y3sV5YMilaXQ2Jga/LJBFMVjkAarJ157p0IFln/iEm1SgXG
wRkUZGu+Ql+FTkf2vQHnqm1BwvIexECzkwTQ5OTjJjUO5k7EB11VQ7KHxTBk5zvT
Kkewp+JQ8GF6WDQ/0s6B1jTUsYNcSXltCxXuSvdV6raMTA1UbiwDjwV3hwZDJosX
m2wtm8MmgHbrKM12xvw3zjSedlXe/6Lqmb7P1aOx1deRzrryGm/2sfEN0iUfwqYI
VSPl+A1eUpGX+EJIf2sUUoCcLNKs4XRDEtAxTa1EnY1kdJKd3HdoZuhhgs7ta0QN
f6LcqqYk59F2VM1v5oZaE2NgX7uFUsVQGuP0DBeP+ZnAYvoao602C13IUvzii7wv
zcC2YOEvwoRbx2D2zhQbz6mMqjEYjRzmbbVeFxyqF6lf8FO1Yh0Q9vNcTocZcFtD
DncyfKr717i/g07TI9+C29crcYUE62mnkah6VWhQUSskwW942FB5ZhhK5oUzT+MB
vSwMHCqTOhSOmOAAZ+XoT0dPGBS9pCV1zDxYw9Cf6jx4woUNeV/07Y1gkKemVhC+
N1vCtwZSPZopEqx268MVMxXMp6ZZIg+gCkXpGymCZ00Ifu8cMO7R2+AL2sDCqMCa
NRIQsEPj3b9wJgHu0fureJ/GAe7+wg4/bidYKcHDxB6MnDxxUNqohejpOgD9g/4N
WYixdTH/X+Q7L7Csx5raZkRgUmWsrAuNtKm7I7R7dEgCbPhVxI7XoZf8A8EkkGMk
+/15Rzd2yLmq9dl4469h8gqKDiPssArJJfGjh1NZmMcb/lFJBsyzhmBs1I6fw+hN
M8q0uaNCY3fDZLjWHWG3Ky46ts5o8RGopsUbfdiRic/MMMv1C3vh1A2HGkJtuaUO
S7qVyXt7bWEi52vRJ5feJGx0a0+enp8j7gu2npCzUgH1EPq3qpfRZedLtW28gzsY
HbnvppzLlc4pgNpUbrlisWF4r2+lRvC5+T7U4yGiudhopTAUHDhzY4JxTqugH93L
B4ZToPdVDTJrMJ5xImaJb0JxbUyhI9aE0PhyUHcnjDNrORQ1Zsi+nyDhdGAblDVZ
q3OTWmE5jW+RO/13kErpImDWHF9uf05ZFwRQlDbxAbyx42DRoTwvIWGmjct1/oC2
q1vS2ATmwHKAaCMOaM2DOurEcuUte2yFiI74tpFMXaLufysy614CGN3PMDfL3TSY
epB4qH9hp3o7bkQ8NtCMhqo+wnf9TgFSsmgkKOQRV5ULUA5CGXwceynzVvQiAw4d
Dlso/unFoPeYLVFusoEr3CKoMuCXsdyzoUJP35y4I+fGq46dhgsHBVs4lRbLj/t3
YUcGmBlSbkq6kknWRCcbZiIof7Qp5GwD++4mCxQ3xBS/U4uMZc4/imjgqrcJfB4H
6TAVucLfy9RniYIWXUVWaGx4nX8oo2Uu+fCmkKqFGoGXnT6rv3mOqQnNYGMkWC69
QsB7JEmHw3dthdKoprQbjr4W8NHWXSbM/uFofX2GPfrQXqHQoREaxFQu1/qx8jqu
hfC3WLUB+hP3LdlAjsyL0Eei+7tIQukvDklcVdpY5N+TfKE047nvcwNooDB0gBOO
jCRw8yAoj0zrjOeSmMFfxw/zmKY88ziQOHDhC7FTQZmGQq9nzpSXqTe+2jpLKVg8
NSL9ucx1ZO2wVzp52FipjrFCUzOKTMFHWqXFYgCXQsgIvdL1nyafkm9MowS692NX
jj8pKLKeaVxBrSrZnM+jZO39H+9SFwZab2dHOf2B9w4N/N2aw7RFWjY0spl64yOi
szp7IrM53n+wN1fIXEA5CSd0O+Kgyk5/DUKoV4Wr3q+BS8Gx9qZNulD09UAOCNRR
2va064NQ/GsGGvmQLpUEpt9pTuz7J/izT/DbaT4ALdi4wL3Eb9N6N+XZvOS0bxl4
6NX424oTXhhuH7YR+g9b8ax3MbEEQF4V5p/qElihOPSySthcnKI4IhjqeZB0oWWo
RIqT6tKoAtEoZ9XON42xt1U8+GwHo0Xrc02CX45bRQe2oeLnO3VgQn+Bh9xS+/7w
jYFxtDkjsYR+x5RQRiKyFHn3zpDr9XvbCmq9xaMOVNtZCahnOklhHOYIh9vcnrL6
kYR2CejrY2ziZs82Dp+2TBd82CjozCOsKQ7y7GfrFS0itjKfLM4cVN072lIqgS9J
0gyVewkTDJ+C0rz5CBJpEpvCBFJ7YA92dAnWCsh2olUq6ErTpOYSTCqrxJj6zeZn
dCamidbHr7rRwls8GGYPNhx45zqOA+2dBkB+NaKDtgAZTUTBYmVB81+aTDOsNpLO
jHiEqnR3C/XS1H+te4elm6r8Q75TR2Tzyp7lS/pGKRLXlpjw55pDYVTJM0xNgryJ
JHvO1kxQ/yyk7iJkyQBGiztOozPhZrBco6JlcFA5x4huSckq4+L6jupL8pbj/xmm
HQWnrRl619AU/YqdPPBVl/sqAzDPPFSgzz3Ku8kJbfDWLF8GEFTlzsNChXLPsF6j
ihAX4lTrGsZjOgrCuxV5a9lUZ7M9nV57D0un1EaxZ8sG+IX5bYlZknWsNPBNj2lo
8R9sSDIhAVKachgwmDhy3hf88W7aa4+WZyroR7T1w50hiWfqwKa7YMzvhsLZnyBV
SzGHJSc9Vi5Nl8vcFZSjZmN4WubJovGgO33JLxun4b+rsRb/D8vMyb8JgWvuPcC0
AArLRHa8RBDWMhcyw1Hk6nGxnOE2u2MOY0c43kdPyUSu5e+3kWu0nEjrrCUOXfzl
2gfCiQlBhcLtdIdo7iii2R+XVEskqAvwghwTFxvmlm4Czdrb6VZCs0lLZeRGKvRF
Pq2SMNaInI/YZqHqccg+8IXPpsRL69F18Cnc1U9UMcM7nlD69WdO+yQba0o1NbC5
3zsrxWpUEBZFo2az7e+uV9aDH7UhkQeNp5qKmPC3mc0PcSuh18ifbPMR7zaYHgUe
jV7dParV4PySbd0IRqiWvmAVY+yNexUJL4jG/JM93IIxLg+UsXN6JTyxYA8zXsA4
tp/VnEsJ8OpW3gNkmJCoVaWTfANR6m+5zh3vFNdHvcx227lOGVxo+Rt6CEvdY0vt
OL6w8W6zooHNI9oOgBGkVjXrHytlk0h3bn5hnxP5ufxnmdzBmer/HA7/HkkhgwxN
kl6zXqExKNovzzAJFH84+Sd7aEL/b9wQFIYI0EDvtA9oXqjI2eIl5X1mOBZz0ltC
KdMEJyffj7C5jn/ASzAfrGMbU3mcGn2zoOVINzjufTeqxDl5tRxKKpcyncrWiQ2K
Zt4Bk3f+HRiUqffhkpyYhw8W/SV8oSROUZ9HcQzy5m44JIGcP6DqDiO26xKTDHn/
XEU+TVK2VVqS7OVM76IlEfkblLvQdb7xcR+gKL2MYk+JYbN3oEq5emqEGNa7c95z
dczHXxAurx28qRNDb4IU9InWUKO2a4uESNRcjwxFTXdxCs8NIrfEOWw3uCKJrOsE
4wUUzxOLPnImtAQfW7ZnNLxIZHtpJ38hPMeAZ5pVUGDsr5cVWYNt5Lr6FZ6urfML
jYbexjsBb9vnwgr90zttHKBiey+BAHkIbT1Onbqrr+6DXdZlPidg2WAB7P/zf9hz
pzDdtv/r4weF2G9FXGghjGL6B+hjs61BaRD+kkbB4HRFD2Txrug+YmpjWjXcJjvP
13JFw1hQJKMgEFbBjlXBvjjJaYHuYOolHi5LnA+3JTv7uvmso2o1Frbg0IwvKNzA
vr3AJ+/asQo5LIi0dyqKBpcwtE5zRknp8wkmpeuzf5sOLFn+RQ0nqTcTqRf8NOm2
wF6VU4PBjaLk9gjfpuYlTeGa+WcvkEWsM8mpLrO+3QQxI0gluej1zr2GFaecMzqX
44uNxOraUKd3pXhgducgfsvoFq4/z3ytIctAkaUChmqjzAIuUiXVeBLHQT1CZSXU
90DCczvYc692SMsMBp9zx6aOlxmsWDN0NUdsobxfNYBD2RfEbUvSx1x9pBOlrACz
vmmIYxHOgkg+KuI3ioiBSvhHgptoCCu0sdELRm+4SQ4vqYtlcMr4SA0LV98uG2nh
QlE//dXngejzH8zvCh5Hz8WlQxfZKHxdQQyLp7F1ny8v12VDdwBd7fR5XigFlJIH
Zsm+mRcQYPqM0YeaP65bZl9PoK01DWFHzf3lv6yruiGTkWLQVmzWdEofrbFGm1t7
KnZnE0vGsdZL+wk+J93T4cCYmGoiNADLt5C3rrcjAXdV6EdN7sM47rGSYkSkDZeT
lrCmLgY11pj2tfQ4F3+U7kYhB2I7zM5noOcSOjxyao+zU7AMMZt2y86moLqFl4Ag
+xTm5dzUWcMfekwY08H4GaYB9s+eJHGQXFuEX3KD0erXYr97Am1zH0iV+ZNdxspo
7ZAeByvj3w1bxnZ5LlrSplFt9MnDsMknng/mpwCB5WqeRib2b0gU8Q+uksLsrBvu
w9eTQnREB4elHoM4EzfDCvSnSwb2THDhSLwAP7DBpfqFLSK4RMUIa3YO991LqQ9Y
4a0YFRjEy9ISWMEzry5RLLfWCsdTMRNrHz0o9gj24KKu+QRu1z1hIQwWtZiH3MWJ
jYidNnvvILYsiO7jkfDy3ortI53EMQNl2MKgyNhBbKQE6AXvGqFsQxT+yDjm7h0Q
JbZ8UZ3R1wHwY7oQITOHe+LhfYCw/bbtQIFCe3fLDLoK84JzE/iiIcEbNULQ0q/S
U3wNlQBo+r3ZegdpT+yLSfMYiRsupylu2slEyFVKr9kn7HnL+YnyKBqDfXjOOpXA
mq7uwpsVp5Hel+SM5ewKlGj54vzH30WL1I7U0lG2KGJM68ycFD/qeXvuLAB9Cenl
4Ikj5AnV6676TGxIusF2FzL4+yMfjLzHQ1oy6oqOBWmGCWkhcOZtriyw10EQ80gM
+XQqfkBzmfPTYZmDePsQZojqqoHuVjZQ1xbkTXJbSrQwo4qawrU151wsIC6VlZLn
iy+fA2TrrpP5fv32Mb93hAio/8Fw/MAri2U1mvmwAr0Qcqmzi/o/HTidMJfVwB2D
I7YmvPHXjY9ECTgkEe8F7wYR8p7maudWVt/Vd32joNcFsd0awerxYRtjlf2959Do
3yV74p/dJW1XjcAj9h0DT74kvCH7gZ1fWPkqMedQtV9DJJ6WscvY0ivhjr7sluoF
PifiJa+KB0ilsPDv/sYUylMM+6CNVmbsaqPTXBWj/7GMv017uXfuNFa4+FZJexN0
CI+Z0Hf7WvHFiUB7phhkqgwGgIUf+z9Oiu5uj0x6i3zqQAHMNQ88/iXZEhErJ5F8
ET5DHYATfNIMDH1Vv64kBmu7oyvRusp6MFZo1rXUavbaobJHx2SwOK/DpVpGYqno
0YtyqnRvuMX/rtioP0MNcXcD4psep0ZPUeHpGEtQwnh9CNb+CydUquxa6m+Ma/Fl
b/A64ldHafPwKFair4sIcw==
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:23 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jdvczy/iYSgWitr7zqG12q7N/kDJ3Aoya3hgV3eYAdttquR8KUHOtjTLT05htqvW
7K8JFSNqg+rzeJQwEGPoC1b1HmYmGeeP+pJXpB2AzuSW93lnAEOQIh/NoHrkjrPL
Ku1D+aTWfR500yBDWbibe50azCpg5NWLWDbLAFzDzN8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 89984)
5DIWHp5nL5k/EEkAxy5o4ocyyXsmiilFgAc3ePckAAmOdEJiPV3dqo0i1P8NsN2K
tQ5XKluKCBG1L2lD6dQOnxBYgTN1V0cXnNGKtJJZPN6Tfw9Yena2z0uQzuRkH3t0
lDHT59I3zo6uNkd8LzrQXYswf5pVOgSd2A7/8i0Wrl+yxnzvmNO5onznaxErwG1B
UGO/6pVm3X/4fAckhs0pOCtpDH7g2wmpfUzi+VxcBDfueMRPbxvtoTPA0I31KsyG
pFPoWtzK74B7c5N2ey//9i0zYMqTdCkvt9ALGmhgrjb1u4RKeouo+jOIxvnCb6B/
Zlh6zy24+s5kBRoPjV7OFMNgO2CQifoFEqa84+4IlkB8KL0EVNFH//OgR2A18mmU
jFQd0DK8+TyESW6AiNgXZpqDoqHm6fyoxfotPtrPl2tNloRDtMA+V6Noi50MR3ce
PwJIyGcfVJS3FmqtwloNBL348/a+88bkizINGXVxSUCt70tlX6VnK00o9uW5Y9tp
Vmqz2mJ3L01Uu7BKXjDsLTDk3RWBfZ/x7UAiLHtamwyNubIn35JGKZ+Q3/gFf/Uw
dSidbu9xYodo8YKNWUxLo/IAdLWk0UJCZWipmS7mPW9/op8D2ioGSEnvgAKtVvq7
GJHOGyMouGc5wyAS5ztOAnn+R3y80E6AJOOdy1M8J9Xm8nZ2Ib61mE8pizVuEVFZ
zGtm9weJpK6GIEY6cLuAK3L3Z5nqb4Uv7NJjueCLFiAlc1gylFabfn1b9ONUNXkY
VXgfdpYhc6SgtL+UPn3K0tOvslGRo6lmF3it0fhXpa7Ht+b8q20c9UMAYlmZjPBK
/0eDALJMOjDVrGI78oPCXNK8q/JUbAx1jf3hJICzaN4xfyUn/VAEw1zZR0SxEGcR
znr14RlfUCB7W8eLfkr+BZKGtfxNKdCuz2EHktl3bPrnDcJ72VeGwY1CiPxR60Ua
jW3SZgGRvtSTXljho39TdI74GG/igxYsqE/rm/GAPef0m5tii5Ncn+braTYUnhT6
k3z489RjVrfPk/R6QH87itKoa8zSvwS8oDaUjvob3qtGdmUIU7dovl0Q+FJ00SFZ
1kZv9GQVYPOd6WMoLlfMAWFQ7CY5spzTt1PX8TJRq/wtypbKKZ2uF0mfCnsDka4a
bUIVctkfAwIluzv2UzKwFrNNdTmFyVkQIDtoVsaIDK4lLsNci9wbRml1HRgPkThx
UvXhv3yHgU00HGbvamN9DBk+uyJ4RFKLjFYN5unMAgNC4sYrOu29Lhj81ORIsMZq
ZECGSD+ICOh1kO/hiYGtzQF3VW+R3mz3cnnp/wyQoriDlMMqjvk4w9Uq15kmYYc8
jsczwJFq2Stjxc2HystO+dEaaWFV6VJamfF1mRokZ+aRJoG85BMLRIuGYL0sdivX
1JR8VvxwAmpxikN1aLq2PwF73ZHl2IbK6dZL2W4xYagO0ztpoofbR9qblvatx4Pf
LvJyABILN5bs8Qd9xcBiIjlbM9mtsdEkbKkXfQ8e30FeHU3k1gI+2gbbKjMjRfOI
yKBp1/58oQX0lZce+g4im8i2OvtHMTyvE9NDQ9o83gSVDR6/wlUaNoTubs6Irzur
xW3l5w/es/lXMZ3ruO7bSZV80kDqSv9P1rvpqWiK7s51S6cwnQ1pWgjT4zNzCGqL
JoS3draxvKobgFJjF9wDkDxVKpHxVjyLXqXj2MpfL4L2DQOcTjmhylzO4XLrjjdN
Bvg14YCI0Xj3VWUL7lj3Dxuj9RM2XLVwemgF3wRYD5YQYiE0FG3Gx/VzZMEeSUS0
5ZdNekpKvoNNmInDSx1ChkFAfAMqZqnPX0NN+BJNuqFRLcU8ki0fxKP/xxGYBR93
7b/tirCW0Q7oca5LBFDfMWwCF9P5exkHwJEPhfbMsaONXF+IIEkTvwMAG5bSUZ4p
KjhoEMkBWRwGShK6vkWcHdwWRAsfLAuyyNlL5WTCi8AKdKe0wJ89QyTu7HX/FQ9z
Pwl/i6N0P/+8aDXhAr65+RXi8Qt0f/DkZsCEIxSf8Lpgub9gDFnpP0Eo67UXQBdP
Ty8OM2ajqKnxBxq2MXAVaEO4DhXoLhNjihsN59DL8loWw3TTK2EdOjSpdyQF9630
75i2Zff44PsFEN7dGmFvB40DDpeqJOnU5Q7a27DrMwUjQPToV9xmdZk0lUZyDZzT
IbKEPyK4fbZ35XjTrwlMZia+0IdDMkWTNgRyZbLn2LLHtCy0OgsVl5ahlD/GimBs
VYPpDw1/0AYHlJKv8i1my8z8lWI8c9mMG/3eTzLPPgDzhQR/VD1xU3gF1N/gsmLB
BUYqMCpaS0umKq6WmFuV5VGDDwfenhsdn5Gc3GorvV4kWEwHj9s6TyhyxfCGh+hP
LcP3fRZUXfziwZnYyEo9/f+3IO7ijZh2PbeOlL4Ky8+SN6sL4pL7mDZaVQFKGQ+U
8tXHFfMqKULrmXgBHr/x5OfD2SsOzOfchng5aU0FEkY0vSxjVIG5P+9o0XNoqcs4
7O5SiC90yRNHoT6y4gxhTjXZvfP+QDNa54agY86QxjpFWXS9THdtZhjn6agQPYXe
24x22E8/j74VMH0AptH6Z4rfQb7ewxuQ3S8Kfwth0YBeLS24YpNs5Qv7XfVPWbez
CGs7vFMivqW0xdJ/34lmIm6HPteIdiF9BlgrWMFJBmmolXt9y3aYUbQ/gHkHEmbu
VdMkkbcAkYNBb/ExGNdtelWnFgDRv05bBNLZyg9a2KZNIBqicnHnJVW36gEXNel4
cHcC+xTgCcTvPRlr573CBoDi0byzin1G72qOaOGeYxPKFeV7fWvepUudyJLC++VB
fhuF+hPTyMxpRta17VpbNci7UhN7VyGknxTsumRsTeSayTxwn1emZqy/fy0THiD3
Scno660CW744VmUZePMJS+6ZUpnG3BNNbMCrcivEg3odimuEx2aqMSsaNzVFM09j
EqDMovre18zxleaBGfF+aa/Yagdp2gpCuCHfdyP8Afkpdt9uL9iGSlUtR/9ERHFF
QGW5Q8m5kZdohgX5TlQQkNSsOsEk4mucklwftBraVCy2yzjSJzfvb+aZIhAz4oRY
M8IwLvPHVVHF6pT8MLwrUyz431fPW7t2UbD+0p9py46xghTTe8xo7a/BCcOm6UgS
vhEHCUUwD+/KgibodByjTs7a9aHWY55Q1I2e7IofVkO23ntwFpk0hd2YQAQICbaV
rh5EAnIpgLqtrX1Ghp0qbxyWcQkhHe2ss3YGVglcTVqZvQ9mKTAsEiNsVh41Ahg1
0o50cMnea2amRRuwjl182dX4MLzebo5fM2mkQNk0ymxGbqEO09lWQVZXALtlWEma
evOF0NNbQ8KcKZ/VHvIh31VgDP8ZNRKTOHcSc6WEkuK7f+FgTx78aR0coRuHm1nc
Vpe+S4JMI6LQ6w7tyaOHcgp1JZpVbCCO3Bt9ZHA/MVID1YAJYyxeFdyZX6La72X+
G2zVf19BRT8HAQVtg8OIL2bbdX+FL9GCBCVtBXNK5kiIMDJaCz3yV8Clf9zp2xvt
V9HXny/CSeJ5SrPCIBX8nbGkvzPPQ7TI03j+2a1TpJQGJNSF/Z5hBGMxssNIXHQV
2fvN+L7OJLhPsEAw+A39sfsd99OVfcsTSU7TSfLXcgH1HgRt1rBzRi0YbuN5CswW
4MFSHC+kqFFU9WunRhp+3OopcJRxXTcw9mRjnMWTW/iGVsi2uaG86+2PPGeacZKc
jegVSyI+iXZtWaFl6wXIuK+DHjCDwlggQX4PawlxdmxNwSKvTEAVkw+I0z+JdvNQ
azWEYKbDbeDe+Acu7S3hfPoD4M8nHxzCxL2CQny62NZ9dZPaeFUHG95Dviuz1jjE
r1SzTYuHWWrX0zP4y6hUcBjnkg1k29XNiJqPkUw45/uHr1lTQTRCByn1+3niaOrn
C19yxubI2UvjdgBttVLDUBnp092JwF+Gm3oRjwNRuOEST3ax32+5D1HP6YiQnxR9
ku6ireH0xFa8j4BHG8ExV82DkFwJp8SfC1qw0q4oYTz6t1iWazLOP4LGhI8TYgLa
ijjL1tFB9XxKgWX20AoDPIRn9ayzPWNFzeGYmbeNdKEl5XS1kJKbExLWl4zLB/Zf
A3/qYepMnw4mqfw5yhqHxtTKdVwxG6mrugTGHQmnEtATggIDJUxtGTk+bDNo1Npa
VdKkn8jyxujYjMdXrmoDqkwrNIznW0oLazZXcKcYcjcOdjqupLE3ssAZ4FiaGaM4
bx6qulIxMVtIoKtPfg5+3mgxIrcZJtwJDp+yLpD4Y1zAfpl85CD/5vDhNjp0zaTM
zIFcta0PdyAl2zkuqLdq42CLqzWvt3fkeV7V6rr056X71TQ6KIZyXqquaAFimnwa
+5U6AVBfT2XT0uV9xRTqXDsF4LDVh0QExUmnaLY0MqfWaCCWYTwWxeKD+BSFUmBh
mCUKuxrFuSZQphV+o3fJQhTIt0fob/UhJewpgPoW5UoiPnMN+kpKImLhs4vlvxU0
ZlBn7TDKzzMeAiHP5oWNt0t973UmCOS2pnomtJKO25rLBgX+6binzW93yEUMyurU
5G5iWd+ZKSitZKBFlC0ps1AxWZ6jf75HML8TRTMOcQHw105Oey9snsxOolf2tBmS
YcrjuAyQFon6CeNjxQcoPX9Wa68v2RrSMm3lWLNBMx8N5A9v03kJbuhhIIr8pLkX
lvqD934a5P1/f1abLEW6CmZYDxUy8doi/1gd2uoAKGJOjwkv9AB6lPk925Xo1daL
1A/yzc1LVdmz6ZPCiWL5ETjT1u5lTdDOr84lcLYcdm2gbdmEwQouUybFk1cvN617
E/OveBgRKx7EiYKKbwj9t66xWLgy5f1GOXr6/3q9NJ0nJG/vqvt0I8KTlg05lvRw
AHLdFDiJVZFD4RTvjd3ibZxAwOygEcy8uQttdgs/Y/2D51RsNFLQyQdinOEzMYF3
yiPYNka1xddiSPDYredzkkB4WZhgkVHce/IrheeZZzMFXggRmgU6+1lMFoviXDru
IX6jPHkHsvtaQ9DpWqEm3hqdZ97ekl/m0f9l6m3zcxz30GWSbrrsO1wzIjQq6sTA
6zJCrglh/jdquGefCyvKzlD+GXww6+/Cb1WC87YGmKY4cUlm8+/mj0Ay6dFC0I0W
9SUNZAJsERs0tEmBAJH0vdt3IjTK3gW+jml/q7qg9HENeLCOA5HmExO1EKGZg29x
Z4x1Q3qslvaYZ1BCV9io0mu6z4myr1jfvXh/oX65ty1zUnC27Caj8NueC2UyR0q8
lh/GEKyKNjBtJNcORKxorp7pZKmbVdzzEXQ3HSVnsPyouRZRCepURSniuwm9nIEE
QwRakLPiF8Xr3ki8rkSmi6X1EdFsj5nQE2Rv9TcZqKjXJVCxFMvkDzEs32GwaV8h
7qjB1m9sZsLbMmvZTQvM8ihl1VDoP6bsRhz8W0omSmcSIaZB11nqaFw6Bgz2HJ5l
QVzOTToC8Sj8piIf1l3+n0+EsaBIgqtb2v4A7okc9ZCbNhS1+WOa88S/o0YHE1+O
pxoncPW1ws1HZ/NyzKiyCK4E99QUV95mkUtLkF7NiZPYOzaTvbHm90DuF7qkZzih
0Kbb5JRnyPLB1610jyI/xbUOHWzT2VDHxV9+CEmn9R4985j7uW9opYowjZYFCO/7
SpsKcJFgk0GKYbQu2yoHCBZwHPqOSxL7JS80j0eOQYCR5GL1LK4r8oNmHESWBrvq
0efa2w2z5/AfkQVd02FcSrz6QXrgPfBnu8tZTWKhiQ6Nn6LPq26isM9WVaMA0F3M
hVUKPRDnifa4hR/77D/+TbyF0TGFBFzEghoWW8DKqQ7eConnsUP9YwmIrOasQvyu
TwDyPmWwFkB+Af+HjjMdcu6CDrtT5V5o9mZgb8xlf1zmEapznaf1YsK0D35ppgH+
qATGy/Jvy3j7d4QHuw7C2vU1jOFurJ8Vy3CzE6pIQT+UqqRr9Fo3S/GJrKiZCIUm
GeCf77iwK1ak4slUA28/enhNvJXVtKgevPypyXa11l8pZv2ugecMXAiMMHk2504b
ooZXJ524EclE3eLfUBKDf03mBWVwNTDtfEHksivXWTw63rMm7R3jIFR988Ve9JX4
11lvKp9cR0XL5ACvLljCphELU0T9BWW1eQq6rEutbaAqPpxaWwyPwtchaWMOtIPk
7TVEgDieA1PtG0nmzrcxhhjW6v/xx1Kw+UK/XgYLwA1Db04opdJhCvgnwmrEyYEx
NaXWLl5IOgN4yxfJU+2AuPbcAa8LlWiT3UiSH7sVtaDOFdGMaHDPEiW9r+5aquJa
vi8PmIRaoyUlRIal7Z96KUOMWV49WZ9krKlYGRgflw3AVa2XJ3+d1nU98t6JiR38
Xj7rOCEK1xyku6sKrGuofx0FPX60Eo9nVtn8mz4qnaXN7rZmvzpBuWt82yURXFgx
5y+LKOd2il7Lm54J2rNE6rcoJzTlFuX1nrFv2v+XfLYdw+hd1rto+v8DxIrE4NiB
ZWy8cL+UMPzD02CinYjmN6Kta/38FLFiW9o5qsuQ6AhM0Ovo7EP535RgPwB04qPC
YbV0R/6fDgZDBUWzZ9vOOpJN0xCuDJXB4FkhhElevA1gRlZq+ceHrZcYe1I+ALUf
PEv9/Hd/GEB+bu+Dl/6TIeA3uMfZL6W3p8GfLT5yS2+5xeGSlga7FPfeBHQqijJn
yY+PzszSvQfqR5mICwOqTy+2TdXqZLbwLZIMuLU3pap1EtD7sg084R6FvUFmfpl+
GcSFhpgyWmCYVSWkcFx30A73/YCDE5GOAs4fKvl3B0WsGsbvXIZsCcv0vrhyJ8W/
phyQON8O3ElOOqyxQjdCAjkCsUdiLFjGMjjq/K8dnS1L64aJyrWMOhjg505zsPAH
1OBjg6PFX47VpEpWfsCE1uMi0ob6IQ7+HSXlczvvKUf4pwdhKcVs9JA6kv/n18vc
MOYic8z6e1KeJRm8aONJ3YNTIa48bLujSqV7vzwh+4Sk9q4tJ+jP10fgT+ayGyyR
G24wQGDNfyO0vbKYZddNudK2FpsZR4IXW3rW94iCCD8YIQzzSBKYUb672Md4XuCH
eS+NGB2HXSQLNsO8eOczIFmYFcY143BbNjZARuFmmlsLIEVNu9GitR0GOQ2fH3UN
EFWDY8nSpvayU4ROrwpvLbLQPfVSk4EwdW+6PXjz3SgiEi+uSELKAUQpSu2NW898
vHSl9ACLNGObJBesOi9yqSMSLg1WoSQbNcSUwpPmQCiJV1CWbwk5wKcIjryLSF1Z
33cenRG//pH/+jILO24SWoKC+PPrCdbWZbObZUj0O07UfIaImuSg1mWTUhzAu1+v
6BoLLv/K2R9QS5yZUsh1CaKmS2vgulCE8xUqKPt3hXV4Kl4nfRbndDDXRmcAR0yK
50E6tYvMfYP4Od7lI0DLjfIqj6YvR7bak2tNBTS2bzI4zgtEc4gcdHFE56QjDoKE
8fN8sIfY4WHG6i+gZPS0ZSwZMYSkCJMLBQ6qPat5Ux9msXWpzzQvUqa5yrGitMu2
fpml6A97ABrLWSPVDi72M9yT+qNVXIVidqJjaJkvEgAkr6/3VwjPyYc1NRu8VJ8t
qGgYbgtfv3W3GzFPkTnPB7Zh/iCked6c8U5MqxrKbZQygcwJA8ZqZnequ4zjoo8l
Da5wyevnXxwPhe4yMU4duyu2KpzZLPIkDkn4TrcVgIOhGxV1xO/C0nMKmsSeEMXz
pPFij1xOib4tZ7PyaBFY/pBopZ12JMor7hunPY2vb0jsGFDxyMmAjidhAk740tP5
tH3w03Pl/g2Bs5SwnA7J/L/NyomJ1KbKTP+G8riRDe5iGqtNIggWoz+S22o1NX1P
xbWUT2EQeWuvtr1kg9bUMdav9YDsWTFAmLONfDusyCkTu0HtpQmyDqeWcQBdUkSf
DQYAmzL1Ea1KvXDGqzs1rMa2l2ovkLBhNWaKxwMbVi7KAqV8z5sLa/5Jg4OnB209
n69l+fNMPLRV0QXDHH2HQLAxpuChZITg8ZapFPCUr0sLDsDTSPZ86tdydlKpRj7b
rNazSh3SKLm3UZjuKXuR7qMwcghwavlowrXIJbjzx5M+fG4x1sGfhzX6A5X8Up1W
S025OTgCRxhBBX/hEkJeAV4lufd96NQ1PYHsQ2RhAppaZzU/TX7ECEpxBrz2rPAh
2rPOZtEYmlGAnV/U1EZDqY2gh1eWeyzP9IsC+VMg4LKM3CHSSLXSCRx6WTTFrQJ4
D8iPMEUPcjug9E77w5gmbA/r/LV0ZxkWKHHP8e4XSMSF5qii6CWZkOuhcymirzM6
rqoDYMDH8WpAOUuOENlCaZW1IaZRsNvfrwQjbC6lmCPxVRFHOk1mhl0ov6MwfFi5
GRbLWeEv+8IZRDF/C8KNs9m/yGGGyV66fkWghemZcMAI8zbLm8lBNV8Q+H7ObDfi
VPd3Up8a1UJJn/XlzKCsrZ29jyAt21WiCNMEESxM6d2pQwAmCNh5WpwkZ5wzp4Za
/Ygq8amTlBtWG4FgJkSA+Pk35NqU9qZECn5RRcmY2GI9zecDd6WsWbkGqXFq4p4l
/UPZz0Nb4+v3gdRqGF0SxOSN7wRBDySYvjqN4p2gJoLwseRQzb9ecyma4UehMcDI
XAzcxg8PmjOOmNisegS/n8sGH1E6NMq3Xe6QVosl48K3KY4LTPAKI5ZTg+8YUkrd
IUfoDAF/x2DYpqn7SlN1cBRf8OK6SMNExBVQGod7WeigvxxdL4SmGQRfAkfwURPB
44+7BEvQLITgPbpacZKwy5IBJ3B0WiLrRtzvGcO9baHRlEASkviXyIpqozHHJIan
S6F/6/nb2lC6RVIFW16FUJIFyGMNAutoySTNCm65o+RUR8/3vkTP5RCSRVT1+h8R
oL1kqtiPjRY5rvxjxYQld+dEnUWm2IHUAEY53ZE+hN8HbErmhoSMLEVypdGo1Cer
CPsLikTPNgvePV5RRJjSKNAyWick7hlamSt5M+oVN5zK/ScO83eoQQqLiq7FOp3n
lOifufOihnfsHKgaN26ctYSa9x5BTokgcYp4xJmbChSeC4mAdB4olSwX0FT1Va2m
cuN5aicLJKPvztDrjBf2t/OYRk1vhM6Z432Pszkeuv/IR46PM2zrdTzg35rxaTSx
j+EOCRfdgbOY6nMfl37zdzt7z7c595JWSI9we+jQE+Ko/wOwArENteBoDCOpMMQo
0slMzUrhc81sGbUtAvLD0dVHU7aKBRWaQgeH1/fF030hQ2OAgK9lVMds/BBBEoGC
Z6Z/KmYCCwCafPjJMdTuAJLCSFqYGJwQTGXuGBEaxUvSsrnRjM+JbG/6J//LFm5R
XIUizmuk+RFoMNDXJvoKh7D8Cte9OHUtOmQ3Ya7P21zDsCENzdp5B6iM0Btw9qVF
cxtwMVk2L6xlq1nBsqQMtFdhRo1KJzZJmjnY6M+A/ahClMzHgSXRubFLvJI94wV6
Bge2FqLjlFmqK8E26nHFu6jA9GUWimbx8aqfpxvpnQZZnyb/xVPZ8QahPoLoFsEj
9viX9a7tpNOsJwL5VTEKqJxIsLP4yTvBma7Xp4WAMyX+JVEooM3vgqJsC2ZQl7xN
4AEoUpXaRMUp0bRRxqfOvQVaz2WSsBVKbEoTc5nF0WAH1nHOywXLFZpbhT10HADO
kSHQiR6FMd5hlFCkUxaxVETU7MRmQGUaCBe0axw79cQG2T3TybErpE5iJ+PuDY0t
xbXBMCZbMqQ/FFHEHcqzlgCmXA+26gUr8la35R5zZMvgrvDteR5P/RjW64jsRUua
tnr8Z1oVl+DRdud1l6uUvyJP/wG1sbUtXjIS9+Cqdx2thPZNYr+JsgRWkLb6Bd8h
L/SvABoto9a9BoZlyZXPLwe818jn5t3Znmd7Q4bgJkwQ9fYOn9MIagkesSRtv6c7
DlcerlvuTvSG5pcIUp/5VP8MjlfOn3twnE71h9i1JJ6AVGB8MtvF8x86rocA64Cd
XJ87MyrKBrS32JMR50wbpGX/EdKq3BiZfzTGPE3B/tMagy3i9l84DDZxz1GnrLr2
m8dhWVk+PwadS95XthXJ+3sEtgEdHXvyrIuH2LzTzCLYUazjcEVytNsE43rk2M9Q
9sw6ZAF/d2K5yRQEd68wOZLzTuxIkTB7A7QjxenrqsS+DoQY41aC2nblOhU67nZg
V+7cHA+AwCLthtPRbggNNl/LYU3Kaa3iljSxT+pC3tS7wg3uZwB5q/arVWv/5wFg
sFD1sv/8ouDnPe2VwHGsHE2z8kJae8NdSpbeuIPpHVV52dELyTo4/LW7y9NfObb8
7SB62uzvNba2TqJHWNOf7K/0eVf45Ihg19NvllzhhCEustBDus9ZJ6sU9zZ024CW
v6J7YiIYCi6KbCKy5MCuHst/JwgoUEOVAmcQ5eewu5+zQWSF7YQIJSl/kqQrUqCa
9glNIpMmwCcNiE622B1NQHAyLiS7Zb9arPo6C/IdTetVhNcwzYvv6zLAE3LCrv5E
LsyXQucyLE+ot/1oXFknqGORO5QlhgypmPomzOPxpulu+qqdwSHn0lTD3zsg9KRk
8Xo52HbHYc7tR/RFpAZEukX70ZsDb1tSsOdQBpXd/0LoFIt2mayk3QfUekfZJ34/
Q23Wo0g19zH8lrL8Keq+b8YG+CW7Q+G4FHIbwkJiEZGZFq7DbeXmnKvQILIZpwsh
9T8HpaOuPt+D40gUVL3clR6vmxj5XhSvzhQKUGtImfU1/8ns1zHag8W3UZTV3bNK
JTsdcTWfCjk2a1X6VzWLZy5ZFbXBWyTKVvuH0JSHtAIKfj+z5AWNiXL6ChBMrbZh
N5/MAPUOhITaUYpoOyr8Rq8gwrioWlGPsTawhktZSn3SFEzdL1XNsFcVlFD4D/L2
gGlOHx2dl36gyL4F601efyXq6ZokO0qshz0FIufbvdhYyS57Ri8sRV7GMUh9FUit
7qxHWXY4RYW0bxClhr1Q4ONQyp6zcxUAFw10yrvcqPCqGggFAGjIMn/5uRJ4ncTs
sTuwlPQh9Ywhlhx1YF+eI1bjvodlA2w53n6GjsDu/ga9Mj1WweTMQmQKGlcAcQqo
+Tv3DdvWrxwqx4+BGvuNKRsns/mfShKs21dXROx3MkKU7ESn/vYRATgU40x9WgJy
uazxBpNiGm0u/2+LMS45UxqY/PZ5P8lSdRCl1m1g5wsk1qItlWxlslga+34QsMqp
RBqDTljfKeg8hbzsIs+cuPR1wOwEFxVzQ5D9deyWRTVYIPteRpczuau1W4TIhjDv
RYg28R62z7b85cMe94vTapNuWvC3BstX0zI7HWimxwQIxnLKJU0k/YjklaIA1rWj
NjZXRLs5+4aP8v5fB3Guo9E28d9KFkQ+zHi9+sRNxX0fWt0e8pkLpxRj/WdtpJJk
bA9qcyJFlHLwbi6t1BdGvz21d3hWk+cQ6RDlq155XyjxYkNFh78+njQMCX9/qBlE
Ud2OHNLQR2g8WqYYcvvtiDbIqVlQOnkeKYpglLwB4QCkfFBDeSBTM5uo5nq9rd3u
+JTuwN/p6gCiG3IKO3IIyZ5Oo+S0fmfcj76i481W3gMw9I2Wl8QwtgSjGPY7AIug
tc+UAMUu0r88muHl/r2n2kpJ5oRheiITaHqsAwJu8KttYi3vzVpAsDHwSZE+lB44
7qvoJlvLVYoyq6E+gnYbsZrTtmoXgNF/i+wd95AEwwYM4oHv1qGtGZi+DZYsQwoH
2d/S51QhG97EyB5pnyUZSdSMFDvfkQvSHjQ9qSTjGg/rEVz0Ndu0SC9/+H750Dw2
hB6uwDWEBMkV54f1E+x3cYvd30MWMPuYlR9uREwqPtxNsqBkX7QtqYzVKTB4oLY1
AZ8N+n2/dUXj9PAJ36OSTRVmS1be0dX39inadISdKq9QjxyvM37SQ63YLx4Esg7V
4jKpEOZSa9Gni4ALVsAfN25kld1LIhMrB0xkHgtH9ub/gb8TvI3iuCF7Vr90H/DG
oJBwl4vGnPQ+XD5HZNyflHNF2MQZBYT6fvXO/EoWc53eZvWBCWX60CnyN72JnTAj
V4NuU9iTQ5Vn1snjljx+JiP/l7zSW2+J8In+NdV92QOhOpmf2/ryoZDYhgv4Rt/Y
JKgJxBp70gvQr9Kpx2wvDSZTHOPD4PWGn2lremjDw5te6f3U5EsuWxg1r7/NWXv4
IsFHKgMgvhIpWEt4/yv8bgdfG2cjiBkniDqWrvJBO6fmO7JAKS0KNx0ATsDP4jBN
k4mDJEnEVgHg8sUeyw5oS+hShXtecQLrAfj4tiFyup1Smum6NDWZgyd5HrJ1O+R1
9+QkJiG0806KxKvJdzz84w1MihdfuPtd1UQpcVwKRDFZ4i0SjdFdrjk9Lb1WOWa/
Wru3AuOPkGrRIMOhKPP0KneGwqlGsDGEDxVMtdDCZG1iTE9P92PgvpAAYE2VZZTc
UXl5hxH+RUCgeOP/4rjJrKKLwg3gOSVPMweyupC6nKrabfC8DsSCAyO7b4iNrWjY
+nAugpvKYYnlqgx4eWS7wgiXWS1+ZKjagcvl7igTqNf8gwNRiDJDgvsa58hcfHlR
Y2zvXYSnv+0DMMehQ3trovw4l5st+tu59GMx0DXSMiELr4Vpsn3ztEviNfivPXXH
BaIvoVTdIxUlqcTwuw6esqOYvSCwKHAWmzO0XhUQyMGJ8U3R9uT/4fp26o80BiCw
fkpc9ICnpkwb9m6FnrTEze1tTTGAlnLbGSJTcL4D+na6CHDbv9sCayR6RjC0q/8V
RTup2r2zhYYGf65TG2iF5tUYCca6hL74VZlEJ/dKmIj0G3kuY+Bve+1e/Wo7GDYM
DhFIyeWDd469xVjQrkXRRsjm+CyvxNFAQE3/PrSOJZvxVEsD7pOVvqtpMTUvgmY+
eBdjLl8kuJHdDR2b/H/DDwk31j8V/ywFPHCWmyhXffNBqNXzuisQOAlmRosib0ag
wTF9IEd3iAAejFZi4MHCHVOOLiy2gs2qW1SZk+DlnGosjWlJy3xzgCUp7gabPDpq
doiYVa25GXT4sRQwOj890l2qBhuFdYrArUfPuCIuvg0Cqx8LjuIhlpUZ5onqRXm9
Kvmb8j6jSIewzjqkgVBobXepAKPWhDygen9eMsR4KgosuKjA3p10e9j9Axn0f3Bn
Hcz8jsIZj5cA1fjJ4ttO4eFQLa3NvzUe4dj3NrgAgKqqokdUXKTtKA4tDaKQhx/C
j8MTl6Nwh+TkUoXJSm/VC9tlQAibWF4Isxt5ie3ASNmLpdNaoh4UaHCvbz1d/Od2
gHDp4TWrr7wVbkOYITqq0z+6FpMq2j+bKn5NAFvN5hb34W6fOnJYTNeLJhbX3Avs
KkX7qF6B02GzfKAbO4+qnRCvmDaLlPeHB8S972WJPjeWw8zlRKCLokXTORV2Y/P5
vpAuzYFG5Yfhg6rvl8E3D89Zz1A8nmoCcYyAIlEzS8MF+ik+dukZ69aNEV7yD87c
14Fskxmb6a5DGJduFbh3nOEJkCEufjfbP/s1OduFbBq354Xla1MuRnp8XEtKeAP2
cqRwGECXVtFPdAo+Fuqv6c0wT097VV5IZFdGeUR24D8hhjT6PDTl7bPVYPLpqRCq
S0bLJYY+eRb3mDaI3EdMvh+QJThgAO+lZSVzF92BKh9Iy1BHXfEVh4c2NOeqcQSd
bNhYrZ+pqJKDL/gg3tXG6N/8G5nJeppvMs/Tejhsjs1qtO1nV9cZ+84codoFMkfm
0oelvz3uMH3Pevlizk5n/IayqLxRBdIsjEzpFMaDQyGAHMIxyl+72cUj+Ek11KND
Tz/xqj+AagJuYaIbvstV2i4nI1UaN6YNmOJ8qNUYHs1InCgxKTK+FD5Edne17SCc
M4pee/wQfLsrvkhXap+nRlxi8nMNHCmrwP2LfA3zXb2lTjcNlxMLFh1fNZU80nn7
pBAcNXM85YRiJh6jg1nH9iOolymLxkhYAQ7uIHF/N9uuddKwjROJliLn2kvi97pR
q5I4OfbbV/5qSDHARZz/jImpoTD7utT+jhsFVrkbnvA2IIlJs4ZFl/di8AqmYC0L
Lp95OR5QZSfn8xKDm5VMNUmzlGBYrb6rGOG4WpHWfw8FWUXykVnvnqb1mXJ5WJ4S
FGNp4eHPMsfxlJ5nd2jfh1qlv3cP+jwzRmwj5oruTyIvtvddCOygdkG0MqnDHQ4U
si72lvvP2+ndkBtgmVA6Lg1jgGXypwpsbgqCwwPzrVFrGKG/md00PfMx4o5E8yli
iaZhCGtoMKJf0pqqvfvNXnOtOZdwcX3S16EmGuOg+/lx8tuzGbMjMhVvoHxcqPAB
TJErFHK7Vk34BtFATZNF+16kSyHwEsfV5jrP6PhywNwH1k+uuKWsoBSNc553ofoL
1gBjdAlmK49jmmNduygY0GgOn4aneuC4rVlabwW1vXsaiIUwNzbqWntmtu03i6W3
9Ow70Y72IFJKGQG9DoMfL6jp6wYsN8ou/ncCg/e0viR8D4dy/cPOpF2o+qA2f6EW
3wG4ANT+83EW3IZI1DIivfo2bamjcTFJ/YPK+meV2Hg89K/HswDaIzc+grLHcAKb
U6TeYhNXVO/Ecw6cVqkFjemxuHNvgSSr7u/J2FiZRbu5cLS02NuFCKO8p6drpPdQ
I7RWz5qMqYdYXqnXoMcKJiS63CWrBOlGB7JliywUawwi0XFtWYS/ZI9VFfD0Rb+S
l4GrHsbqXjkYrv4qGNcUTg/2B13HbHtq/mtu2eaSsCrxVd6/cujPrAyvUc5nphKV
+5+t1QyvhYd7eRD7L2ZYoD4IHTwmo+U8uo2KPaAWsgRoTkfEqvisibj0M8/cnJAL
ccRTBQLddkuUI/z0I+dkL/hZFRsJSUAjrw0IuAgnp8wb9zJ80DfeCoosaShgjR3X
JZU+sIOsie0x5Jk7cvkcK5YcZ40BoDaFS4htjfWjkRZtd6wWmhz98h15cEbZBdsp
qRUKbx3lHtFo5ADisUcfq/+q2fb64rPEX8D8LuDP/vi9GeY+uZpGV98mXAG4DlZU
VLudtJllSOWdvBoPuWbyINQ3cOgMe+Ss7IScbKl8UKXXa2rstUoHFEQ64EhA4fdW
sUyaERLgO+89S/3n5KXl/rmXBiN9eH4E34aG0BS70PhaU2oF6/J1Z9xnAsPzk9lg
kL+QGh3DGtf187Ym4eOweL1ldDCuc48W5OBNIM8EmL2HYwrp9LhgPu7w7b+kZdA/
w9IMAmqOVLBvgBbVm/sKO1HjLODp3xTDc0A5aNgIQEPeMJkLflfyHKyRRTvg/g4r
c8PJu501lpaP/j0PtJibM5mNZwI/A5FgoP/03ZfvxDl8waLBYBHR4j1N+cmvjVo6
8fnwRHcYCiiX2CFTbkSxD7K/hhyJf+UCdNQOpHcpOGJCyHPXg8Vg5iKM40UHRIpS
3dwp8me1aeJ7JXqrnl4Oht50v4OWWi5SK4gP4itw/70l0svjjJjN0sdVTptOK87v
nJDjNVColRiqEJXcJ1xGEggEMZ804ilk5/Q440krZ/ti0JxWUNvrpy8PjqxI419o
kMfPZadFJ/tFxhBInOaGjVec6kryb65BUxsLRITrWUR2tpr7Qf4lcpVAvxi4OIQi
At7J6g87ZCyyiz8e2AzXKW/hQFdZsDOHRzRhdRuCXfvuoh8YMxd3I4+EG1qTYw5G
HBEQBMpDRJBLOTSY0vqFD/TuDhU6hXmyBpt/tmS54LEvA0l574yS+r9HqesUUGBG
vTZa+U6xzTn1tZmvkNJ5E9hPyM0u+mqs0EjsgPb9Y4DotAojCEYtsEJOa5rvO6h4
FybfwWW30Ehekwp3VMZWYnI3J0P69+cufQBajQdsYazDOYMIuR4ldIhZsDiaI7a2
WQ7M71vZhjwmLv3zFankfwgHYjTS0VHNywVRh6SUAIBOodXUtsGkTq/+29rLx6dO
PBeUKWRnwCP+YG6O9Z5zH98R0hy7+W/bTuR2vE7RODvCVBsZSKNukq7OZKRaItP6
u9BMygQUQD2wsM08J6e1lx6L8QFglBWNWCiN8Fsmyx242v81GVFsd/9d5N19sny8
bWVwXFoEft66xUPJRx9xwlI/1WUqrG9WLH/9Nrx3iMgh+eEyrvfnj7Gffl5opIlb
4qYMLm2Mtw5D+cQSAC4hxB5ZYXqzNOI6Pfjsroy1uetotRwBsSMogS8USZHHdjFx
9hmn3M1r/xULAurHfmTW6NSQ25yhp657u6BREPf8uRw+n4ke+StALQnbhAOkKi9A
IrW9Fckwlkg977injgtcJTkxW3UWveRiEuQaIHaxPzXxstcwOxR0DeffgXzNhyN/
xeBNKfzYRtmmfvOwEHv8+b6lszh2XIgJ9L26QbsmJ/M3I+iAqn1P7u/DZRLSRFRk
1xP7qqk8ntcMZQV1Ge17DU52CxtZxQZhZFnkC54MUXKC6Aslv+zC4yBsz7sei7AG
F2hShNBle/u4hIfnXmIjkqH5a+wdg6UQ8QAlCJgR8ziStWFqdGcJw9aKu5RnRokO
kkwC3BA/ArDoi01S7Xj8l8ld4lyWwudD2IuQecH/6VsjOFEJHfOSXWl+DlrtIvUE
vfe4jZwSJaDHz/i3YEFkwtqSrntcfrwtmcmYoEs8tFaDNZfSILsL1aXWA/cf18n9
t+TZHlgaIFBWwcBeph0Rsfvocbm9nN8+lZ7IJzhoc8uTTQWp6S4SYCmrDjXCx5HA
c4h85AlybOOacaV3vf3/wurYsRb3NjZdvXqavUbCGRXnu9HpXJ7WedNMxPevUbkO
kmru/C2HUq5SDv1Pefdv6HzsJHL9Wg5Q6gbgCd7/KIQfEc8MYpUBU0FSqGGHnFFG
mesAsK+oP7cXCBzvcIIfdAs4h0GwgwFh4MQhOp/jjQ4Y2ABwxT5tLadPrmBeM2w6
nLjNUuhZlwg7gsZv91dtzkIvCmLrw6EXyknl4sub99wuKe1LiGVMQ+XPBPKOYYa1
cOnRxNVuWO6rzCHXP8Jy2DZpSHXMDOfKF2PHdiNgX4pv/1oja1DJARO6n6SLtMSo
UYU+6BZwxlFaT7cjvtl2dGnLPntSkvcKlIKNbeDFmXzf6/C5W7KJbOx5DPwsvdSt
EJ8qHVUU7cexDiHBSig0tqz68ZaG26WFolQ/KKTeZM2mBcISlB8ofa321Du2rEem
96HRBkumDTeDCVu8SWj7EoTs4druAJKtdoxz11R+LV9k0L08P/k1I+FQn7seBeyC
E5FMkH45x8aOC0HEVHl1fUKjVpvJK8JclBtDeAMsz3cYzpYFz4vSbz0Ep/M74Dtc
2OmSCzNCbLbagTYy0Z6zN87ZUjNP/wWQzq3AQXeUNqSngHTL3wqzP6MAbYiFct6I
DV290y9OENsiWAgJXDOBoEyRP6NWu+6r1xUXt+4o4GCOKNIDryZs9c9d7/JPeSQU
HxYKXPHtMWLQ7OBo7Cs3ZpM5DZPZUCx7nZxmJME6gYbUMiPkVqDtIq+1BGrFSIbL
kcawl+rXRgfn+3kUkn0HDDsqrp3XvJ8HFGa6x9T7apxR8IO7YbE4ECDboM70PARN
TMJdVZGF6EOQ6Gn+RZw6Xl8lAHm/QjhEzR2ctJBXV3n5Uh0yZ8zgnSfZ22jCTBs4
Lbiv7hNTrG433hHVSPqFwgNmvPexRjDEt5f5ldlfkHR3v3SGCaTXLlan7mDY/Y/P
vo2nftScqReMYB6oeANhFgetjo3+QrDX7r1INsGGAQ/M6w4Fs0b5LIsrI06DMwK0
Uy5Rl/AveKt38oc+7NzhabtOS1w0hg+YCIyhYG6wN21Y4LZZOwTcCNQ87+QYGg6z
K1wrnfp0R0YrS2KOEwQSwOwGeZu7lj9w/RFGg/Gg4lXkLxc8XhzEdPj0Yan/oJvF
6J1qb2dTQ+6rBB3yiTOtd7aWscAaXwASVg7jP1zS1CKQxWb/BUzsey8D/ep4DJU8
iTZR+1w2T6xOQzLVUuUNSp/H9HvH9onSZDFWejdlFX8Dl32EP/EjyZouE+co3zm1
I0iVE0OafrTucirK/MVoxj8QQTYiCviL3gLqCe8fqpsjLJNm73ALhabAQeGNo0uP
Qg2inFz9Sui3PWVxUNGs+S5g+nv7bc0pVLbsmFWnwIRfAMC7Duhutuh/Q3NCGIY/
BwIxPizk0aUkDTn4oh3am44g7xXw/G68irJYS+zQGiFZNSUWG3U9di4UzkTy7KaI
MZ/HzBcnzY35QQ96Nk3TKtSfrSMnWYgULzJYRXkQIrcJ8qt7v7g64lPMo3Mudqbs
S/y68Gmz6viuTTIVNmGRoYnrKVQAP9AAk5rQUVxzzcDcGTm72udufLCz+k7u/afe
aPDcJdoBIiheBShm/uaWkGPDHehmSpzUpQHz2oay+2vaeTiyp5QZe+8birqL/7QQ
WQTaI74PwsF8UmSO/c/iNMXhvICdw+YoPF+aVEXqCvha2fUJ1VfM+aUWegu+s/KR
OjGihbz7pXJDIWEtAdUo5pLfVnTtgqdHWmMWjAdNe98EaZbkR/MqCvrDO1T5N3AR
JNf51pcWnV6jk02LFh7N9q0lRan6tvsJIPh0yzwcLBa1D+rVZILTK8bWHbrp9MFZ
qOeaS/v7FSq2NfRuE8F13hBdGv4RmP2vZPjGI/kzeV3v68RHP9JUvJgFI5x0xxx9
5q62M8lwvA4Tnb4c04N/wDlDcawtSFj/s8ADfuBHzB3q0ujP+wxHC6FD+gQ2RMYs
E41/1xAehxr7eBb+FJDBUAUIhKe7qhxX9oA6Hdp2Lg1xD1ilcrDUnw4q+g3ImNJf
kuLvy6Rkv3RAEblkbphypEFz2qRdO3AdysDf0DbOiu01P15pDWOShtn164PkJ94Y
vpwB+jpEhwXXs83PZajpy/+mcbRc3bQXhVNHjEx5ROY7dbN+wyaBLbiF74rjJ261
aHCDHjc+7afXITRQuT+6nHmm96OJEldYiAXQbv2w+NbMtcfryEg3XTNEI/deH4In
eef8HIPVmMjRWKmNKnn2ZILl7W7CXoyUK6Wh9xZO2EoW0Hk03VwnvctIVk0QUqP8
AbcMVnjF2rjQ13VSn48WPAGBLZ4CjN9Hkd1gorwwGr5+4e3PZ9G5pNUnnEldkBxc
Ey26rAuXUg0q5WZRY3o+Z+qWZge3tBXKV59rpElDG9iF2jJay8/+JDg/PJGRt88w
UXm24QO52uMR1uqjUlmJ6RiV8w5cxOB2sOBZ5NRcy3uPnAGXyvpZH3EAsTvFbzE4
rTtfNAwI+XYzI9XDLRFa/WYtO717vw5q9eP5+jHKNmoo8vFp6rhWf8YLafK0vH1u
qZPzN9jusbJJ3WDPxsc2qZdYAQff1hRKrEZvmnTM5m7K+h4mXV3v6+diWhueaTtq
Ig6C35zYWN8ZJKvBKYzSsPpZeWbOeCRtWRTgDpFJnvH7y7v32G29FYm+X+10QsAS
NQpbmMoGXmcFXZCzvnfJ46m3LEPGlxvhrTYUrc5rPOU5WYxqcXHvI9w9rU142jA4
ALnSMM0FVpDM4jvaI9na7irVCasDFIMuAB0J9NUzz3PChKb2Zjb3BrVItRZE19gJ
Cz0n/wfNuo7EwGOKbfmbl/rHdWcPEUHVMlwTf2KImumNhh51lcnOLVb2e8tFV9X5
W5goRFHt1iGgeIK7ioQTbxs37Z/gaY0jgDztlXahs2VOIBWKttNB40Lw6YWcWQ2h
AzJkUR/6V0hqCMk+lasO8A3xlNIkRd9c7dSenLuzyT0/vHKP7KUr61Naofh8cURZ
vehAAO5/XVsye+jp3V5L66pHNTflyBuWqSsXRkbOwoHXXhxMG0th6C7taSdjNBbY
vMPjI8WHbCgmQnCwlC1EKk6GfnrEc4cVr2ujg2hJ8uEmjBXn2uDMhBgHVCZs42vk
EGVB29xZgiJC5v110fr1Mm1YiBYCueTvpDLF2SYQT1M0YxJGYaSFVcRZB2aC/bsR
jAMZixMWC3LzF0YnwBcMoT4VSa7GDkx2+JKfwm1ZSj4GzDyXVkSc2KT+i8TLE7Dx
rAuCmX/lm+Cg5IQmgS+IxXIikqtaZKSpTd6ftkglFM+fq5KEh2gyinLQr9Lay+Z/
rWjENaJ0pJzMXSfbT5viks2k6jLxh+QhhLynObPXZqloubypBU7xGki0kao1BUKx
6ND6Ilm9izqIoUC79EZTU9njv61KGsi4IYYiTY26dqDbRTCkeYsRZj01cBW2ARFY
eJmecpxN1mx576PHF0eOuhpUKjTV1KV4YQcNM9DQs1asEAZH7rlmkhLoyO+Plg3y
TdeVccGo6WfF2mbFU9mU4nl5pEv8PccQa6wW3f1KYkd9eqxJmKW1BBlAF4YjnHtP
viXLaItwNBmE5AeBG00zZzL78W7huP5UeA1VQ0WlgXbGOOz+qKG6DWDLgwkm2cu4
1/w7afmSKXmLIEOmFKIKh4j0k8s6Ubkx/koMEv5PV7wJTMixCk/gA2tN6mMMinec
QKm8BII7zYsKHkSPiqiqum4pSpe2jev2Y9hdgTmWE2j29mIciCUDIP9GucWeLt4m
AB+O2YXeZwDqI+/cCpP5jXewWcMzovcLN487RBeCN4TcaqBYA0m4DfKOI2elX5vf
d/auNf+qqTFcIW4IFTzSYDwZUHnm+CMZgepjinGvKmt/TfT2JTL9K2xovTj2XmmU
fPfoig6QsEKpOKXhSqy1GDpjrtIXCTxPJ2zb7QIDB+CM6YH2Slr5IsWQ+fU2sAbT
d81+i4Gd+lDIrhGvF7a4+ne5YIKWQd/g9isksbpyRih0zWm9zPDA+72O31taYVST
977d6yhCi2o3FRlTucCVWgVmqS2+4g32Etn2+MySk4kyNV8of1kr5qTdNkFhd5ek
1aBpJeESANvWAbnycXkOj9U5Rw3q7otnMX9KyBeWmc0zptY7c4/fLyBTIbRbTlN3
rb00P81igwXNhkb2/WSzcEe4WDj8GTqlbE8MhVwKXhsSskkiveA+rx7F6vUBi4eg
YG62LconIR3YTfbb8wdvM4tAMjblvoaoH+yPXC/tmfML2OUbhXjZMfosWuCtjp9+
ALb8uOWK5tU/CeLOKMaMmTa1yLzJN27G4eMkE2yiL0IMKBcRlq8rKsyZJBg9wxQw
IF87bO4Qp/3MTnN4LfzHHwEp2iqM/oWCYhCN5jd36tUJfjb6Fg2qF3W5P70Xp6E7
23fUngwCmtcaegLXUiw01kokuWR2WnNLl1t46p6qxdapUb3v0EH141YexH8861Sr
cLInNLOxlQ1kUG1EqB1bg08DwR3iJNVpR64aIfJbVugNRizADZN/3NkqRom0MOt+
ReWJhzwUQyY9RtfenDcWJrD5GnoMYag1w9idcXp02+SFwz5a+y1XTbfcH69OvwuV
ZE+jN2/vJlvhK+Mkzk1NdzTiKyrkT/q6WSGr1IUhx+sBIL8Rx0igc+89JMpdgL+K
rw2y6ZLvZgTy1KgdxJtHhcfDFeV8j9Cjr13g7aRhKuaYbDlpbl6Hxnf4o/CPPgXj
xycX446sKpcLox18qsXxuzWW7kS6va3BcXhtJLSB57qMJwTMYeVKBRB5wYpghChR
ESgX5MZMQkBlOuGiuwqO6DMIFoegw9Zuglwp4ZoDgG0yQs4CUQ3Z1XH5TqfE3LHY
l6I8NktHCGVVDCKerj14RMghrCh3+aNFVTQAwX7dX32f8cZPKpAAQ/ceuiVkmwbh
XpWh4p+tyPkWx98/mbxznY2EfZXYDnrQXch8AVOfsKkRXCHQKCtQzc1TvsYKmyiV
5ZbeFnU5+WavlH2JBstrbaG//WpCKT35K/RWBpTkwWRRk1MPQGEAboBw2gqxBCDs
rZ2OpqyrtC5Ug3f2uBIRrd+ugKmnnVFB+BdAM9ETW+xLP7QlNCKBRVZdKYSjTLdi
IIm0wdWvxjiPvbwDXX0WVmefkTgIInsR+TTeIhEuJgysAMA+zMAkXZlPbU0+MLtv
2Ruf3GUKE4pkh9S0/l2KO3ITcG+SSTEYk/6vMmVN5RzjlrDXQAemmaH05bOYCe1r
Sc7moSwWvpidy38TIqeyXiCRr2BGQKZm4yORywr3DYcUV2Orvl09HPQaBv9mNLYY
30jtCeF8MP0eL7AggzqRRGOh+Z5yKKYcy86u2dROYXeT6vw441UwSamCjzY39sxP
Y+5YCpiiS85BSdbcuEb/g4R8WK0Y8/Fq8z/FYpf/FAuTmFyqpfWMz7CDs05M1CwU
8UL6wc5utzN+9yQ30Azs95OXSl/Ggs+OuN7wbPJoCX9xT8mI9F5wOl3cjWM+PCE9
Rf2+KlEOWKbhrR084Rd5jswbIWeplrC31y95Dwr5vif457iCCZlmqWsI9K32wber
aiF3u7D+v+mQltHlKeFsKD5Htt2G40NSbbolJgaufAXBbMpX+/lcOmWc+qBFPXXR
xQFZCsmSfX/gICGgvDgwAt5N5C8Zj7hBuT/1TycmY6pwm2Ql8OhurZcsCDJgQ6Dh
UaiZ8p5w071dJHzGYw6MxMKIQastZggJ7LuAbakTtgmF7e/l0s1J3YKwj/8dkRNf
T5EvDRGNqRtxYhhqfB2CdXEmfe9HGxqf4Rnes7IKywYTvbqNYb/2rINN3FgLTsur
iP7GCgfqqC0Nnzs19gx4pakIV3JSqPHKKPFo8Gsu1Gsa9lwAFdb9ajluiEBFdU/a
BsvlvgECWcz7mkuJsD4PtTRoVZweUfoB9loZXBG0srzp2Zt2vcfOgrq0k0X5HjrO
tgPzsH7MxqyfM9osEy/1q+K+Xnevau65Waer1N7Lq8voG0znwV04cYR2BrHlLDEE
Dk3FCUjiwWGExvIMCGnc3klsmh1etBRWm5Jiik8CrMB+xB2YEfrpi6XZL8UoSUPC
yAotsrzdRd8GueDK3PDSZHm5FDj+Jp39p+Sz7v7PNBcXCWOn6hChRrZck/b2NefH
WOBMu0WpN4HRawQ5CH3GX6pY8zvALgTzdNgAkLIqh/nFETScAPCtR999PSsL7MsM
2L6sCFIAuYkJ81Yy4wiz6U77ccTI6n9HaaCVcctB4a9pnYfGgDtYg+yHInqDwUPT
Xq4p0x/V4SPxqHgr7+0eK52kR7LZMcjdIDkhkSkGC5HXEP3naRWLaFEwtjvfQWWk
BJU8Dqkx6YH8TzMYVzbj0eBiU81e/okMd8Mg+PY/2tEBQyedwhYKRmemfSx1aV+n
xsWci+npjTaaZMNEiopKUTOd50BKX0OwFIkKI23R3esfu9c7mdmqrVJlceNwkpOx
x+NIlSGa5BXMRmPVRoiuey4TLi9irI60bZ0y+nVTPN/dVYrYkBd9OX+iPlswayPf
dJZfYOvOHozjO1yGf5DVoZuzVKPE8kI0IhbSRq4Wkw3JZykg/Lnd7PRjTMcBoqYc
08rGgNKJa/7GQJXwbWuw9KnJpDN7NpUBHsNxUJKt2+Zb+Mu2ZpdXE196T8deujta
Ns5k4Z3retl9AC0ss5CS17JOq6E36jpvEkdt2jkZEbxQSGW+z1Xa3gEMWHAOK7LN
SGLYETAyyfFLm79BR0dySf2Lj8P8ZsGI4uNOdQTyKF/vO9azNXSyx5yhwhXEQ6uP
8HG6PAFz3okPIv2dFeZe/8AwwW4OB1ZN9dNrRwPxcbJaAbdd8tB0YverxTme+Bmg
/5m4mcqFhI8cgqucUdIMDmXSU3r4VexYKHdgFTH7so0wgoRHVjxlA9oC60t+zufH
CgFd3el+81QnG0ITBRSxBOG9CGl4k0Fal+/R3R/itgSHl9csLdkwmo8z7b8ZFHkH
O/jV+vlJzOHYFfwO6AuTPCf1yUX7GHP7tqDw/yiQhuGewxUb6uAHEJWW3YglLyd/
NpAy79/2BRK9BJLetitWJ1wU15H5ibrxfLrEq0Ivshwdan2A8SrIZ2RKjpetCX71
CdgFrHvsqXcTOBsGgjaNaZcr+Kp1bZUpXkmBtWzgk9lOQBa0pOD5fFdxVgSLcb9f
2pfIcCDnjgGIA/+sZGG78dESYIdf+8eQF0dmrSVVsYFO4gYQF9Y2FWLvd2q1sD9X
Ku23gad5/86mYjizTxKLvRNlnQcDWDSawKQwt5kOhpw3LiEKOiwXh+ZdwUNCpEwd
vET4w3kUUv8NUci/7CFPJ6Npgyo4a5isLdDrW/3liBYkmocevMvNKeFS5x8NlDHw
Pjktt5E49zcMzDnkdevA64elmReQ9YSh8QYVFMXbABvACDlYsIYYq+AeZWAwOBC2
kAqwACKbNqKuUo2dQ4rhvAPAoPkBBOSGEArT6RhnCAP2EixeAMs7FK1NX3q+Q5sz
ooh30FE70t8F8M3EADuby/MBNNS/ya/DQ1Z9iMhvsL6S3I2XPUpyXlqFABuzePBT
UjjGtZT7z2xA8/kuKbbQpKyk6ncUkBSB084i5rPOA12KHGmMgHue+YQsPFypimOs
ExkEwOD8Tst48W4/yHvNaQwBEx3IsuoJvnJ+dDpkQiq+KjX1mafLh1wicjSkqV9W
+saeHEq4QjBgGRF0AfqnnkHUmiQJBEyZ8r64SHD3OJbmCTOPDoVRxSy8+AL6DS15
sEWs340wuQSc093pf6fHmSmwFh1YoRkGmSouzwrEiQR8hZSEjaYoiw6//dQq/qq+
X22Naac9Neh7gYaq4Jq5uOyuGlfIjakcl0DmJ11yePyOZtyTf1JYp70qZD74oze3
THCs3CUq1RasQ3/waoHhVLY7I3mG7SqS+6G+T5Jqa15R5ouF2IQZknTPRmDg5bBs
0zRYYCnWSvmn1PdecBVfZ60TkJBeKhYXSCAHMWYNjLjLvUsDkTREs6NSEQSlvDPO
1PSdtRif1KH/Un0Tjm99vKIda0K4M1wMZ4S3VOa27BDv9tttS/w/19EaQmy/C/fY
QFrPmeJ2mMdl8xzn9+8naxcXIeF1ITLlwu1c/wuSPpKbd1JbOstLHpPcwl6MSusW
y7hlNCo/1f5LSKLgQxAwHbdOP/RqGDpPD26hv5wFvwEd2abM/da6JMTutDOdautd
ha2TFK26GnQ7Zo2n5tTuY99lbXwwq0EJshtJe1V36hIjrQ5BFJYW8weQsoyMIeQw
dgyZ2H93QVdy5jK9QBzxdtcTSIpWAOHp2sF0nKUF1CNnbV3zk/WahaxjlddBs3qK
9LtRJyFxw9K+f5/IuyJSEAR0GnM+Pjo4fd8PPCGzKqUMVmQIQq+9r4cjkeR7e+1D
BILH3gqP2aNAbkDr7sn9myQyJtNiUXjWwP4WUYmGzRUN/zKeTg8wMEs+wXrv5v45
/jIk7qt7YfW4rpopKn7ObIPMPFgrEBjJCsuSlfN4gtrSAY1/bR3IrR6lfsHRbm12
Oyppj/fsv6hkuSRTvoOfEqlLmnkBswxAnIM3K3OkXxuwpBRB396LEuEtfQk4ZBev
IeoxXUB7iQ38k8b9f5pl2lsObIN0vQthSRsnh7LWrnrxNnWn0Fxmvux30eujh1Wj
IEqNeS1W04SzURzzf/dYbtQW1uuAe/+Za+FLYE+XXtYGTDlM5qg0lZdD3EnDqcsq
AVVouuWDlSJCUWfzAS1hV3Uf03IbPQi0N0q8iumGJSticUJeYkwqssP1ZvtoqB8G
QHnOewvj6qz1LuTZSCIXicbk6SQ1KtB0PYKqqdvIE34VwILtg+NvzDrp0dyr5xcH
94r01bFvBrlMsf/NX3889tqCl8bf/AZIvkyEIMcuSEh0C0ZqINTQn1sN86Oe//3j
deQsyU1i/jVExuwhM6xymYY1Iv6K56OnvWQ9+IDmkhPlPBvx6wPBjwffRhc9Thrl
lsOPOQCdytKno40bivooe0jgOuYpK2F9re6i9+44EnbHtAmd2z0f2KaGD2nG0J5l
O/fhqS/bEkbREp86yUpEOGo0fzn/XS3iEN2Q4Ba6lyuxgE7CItIFct6Sn7S9lzbv
+1MJflI5NYj/zf013g5/SqAt9DNI9HpboRr/eNj5R41t5Wh6uq7z35dbL8V6ir3Q
ecQr7S5TwKd59gSz6kIxSgnIilJNCAOz6DSglxmq+BR1xvRNb3ovspWevMj0rjQM
4qcsgx6B7K4MrtVT7BH5vaHLlyP/4djUlTnIg4/IzrIWsDMHUTblfo4oljw/6McG
ZHpNQmzONXfbAV1WMeHqkFOW3dflPjAT/VDJMAFAMED9KO3r92dQWJ7k7nX49r/h
bXbMgvVBrykE9zzT6n5RNu2nC9ecXT5mS2uODleRApv+ixQ4vILNF2+xqsu83h27
003bRjlYr4Q/bZTVrmGzL/vpplNWZOdvc8EdxbGH/8Lu/CdPs40UIhQ1z8xfa+OE
etwRDPb2Uqg1B2yzOMMkeGuN6hkr/C0o8SMsGQteA4+u5Qus59ZP6QEqZzdAVgva
tZ7k0xYTR3U3yxBmFG2a6VLAtJIvZzss0syuqBm9bxoOgw+Vi0HTP0FCcwambvIG
XVqxIn0P6Pzs6YSdZtRnecgncsL8b+La2b9+s/AZ92QrY89p78eMk6vurnSFSE3F
rMw/kMOrRnXL/uApCsL/SyK2b/HTfBKgicZm1ZIvfm1pNgD6by9Umlj9EAPJhqui
msbNyfIOe6qcNpCx6Z45jJhhxl5Fec0Qpi9I1UaZYk16FWH/uEBWSup+140BEJjU
ZeKtXNs/qoCPzxwsaCgxfMgnKK1Tbrht2oCcLe2fZ4HZt6HNRwP8yZNvlaoP++BV
EFduqh6QyViyLPaiUqs6m0qm/0ox8U8OQisE8PqW5cH7M/lP9+6VBz+zTKpZiseO
oFJWUELiWt1M82rjVsjJGWF7gi3ztphOmsKhbxEDFzWvLKQ22cieg16XcPxrmIv6
KJkrdqMUd7ny3KSHosOpUYsQIYEcM/OJW5IeuI7r5g2oGrWZmFX2p5T8mU59NB+4
oFELYTCc5G1ZquiI9cVwfIyziVEKS0d7p8Keo/QslMK4Te29NXR+CkpqTlr5JCkB
kbYsPjzJTOwxslUbJaxOfsWhVySS62DNGMZ986v7RnyXlL3xKuPivPTW458MCjE5
dKOt1mO8c6a44dSbN0OFXqmWogpgYzBVwauzv2ZMfnnDi+BTD7stdsaKF+2MAQ4H
tt2r/ZqzRsYOFCXm7vYziN2h9Iyv9q2lFqoXzqXeiHJGrJYmSh3IPA+hzuck7C9S
K4ZK78RhygKgm2MiMv3ibJ9X+sWJhwSNyXAUNXS2h9bRxUbvGv/DrwQ1J2VLLeeB
OJV0Ks4FWqSNReqaI+1bM9H/pzMiLyPA/vQgO6aZYcR5/NcYHqSelWhnH1yT53nf
QFGkE1lVeu/ts3Is4naZ8oaShY9DvfetyAaMu/1Xv4pYTj1HA0YIPP5xCbct12zo
cTHAVp8r4ogaCMRlgpkZupQk+9uIa2TC2YnN8Vlzd/XjqljAOyW/PoZLiCHVUo85
Yh+fzHmLIi3ZlgLIBdlJ6iqotilIzeC0wS5nHbNCA76QPlzYRf5rzWh4RUazxM4G
CmnlkdSQ987+hocfmmHjOU6fLpp7mP6NsqSN47gK+csLhsA3yAWteiBaIWOoHyuw
hGm9ZrOgRWvfByfni/0L6Hu1bF3jeqnfEhh7rncnnoD5sUEqEf3ZHH/kTrrpC+CB
LWTW1KZInKi9++abnU35LH3NLbEP3Pt5wvPA5VAG8E+AVw6kAYL8wfWFctaAecaH
pniObTWqgINP19sgY5fcmM0UOTciTG1YLGfuVKqjbzG2Egx16hMEM0RWPF9qDJJ3
KsQDsWlIBJpD9iMwvff+ZaaEQ4yWWCV6qAHh0cDvux3azoQjJnyDMGiKAMTIwbhy
MIQ3s3mfVQ4HWOmIR/bBTwpeb5OGyL5Np7sdLG/nquhUcsFxvznKbleRxGtaqkXR
VDwTIwnfSFpM8Y7UuxaWPiG1sRqC0IVLTfC2xk+NUYM5W+yKXJ+HkpTz1ZUQE/1X
wzONAnuaTk1cA22b+8QnGaz6jVTbw214SQbQGkFk9owS/xogGOCuCEBw95uqN9d0
G52seJExDWlm6gcMB3gqNUqrCS3iZtOm1Ocf0MxPpzbmv5qlM1mw1cFLF6VbX/na
ULVUTWuJDjWRZMPQsgaXGyOCQbokMBSgff8g5Elm1KupDBRx5V41MS88h2bpUx1R
K5xu6psZb8Ab1N8zT7HoZx5C1crS5r3BUyza+Qk9YsqS8/8XBTGg7ZlkhiW2Dl06
watfT4CHyohZBDw/jWfhC0UuLArSjEBE5FRuXDMEG4xE4H4YQ27EnnGjB+pnZoGd
T1i+4LUMShurQSskDe4leUQGjzNhpaX8VjHDh54F9RBhouSqCXfHn8WqEdUBR400
KSYMc1dVIry9id30DH8KPnPBI3U/2WmxK9yQyQ8iTPq9qk9jGyoiP4apNyWOZioB
1oYg640h1w41Ipk1nqRQyh4gaNkTa3TEJwuHcG+d+dKSnhsvQtVI4ObGNru5G//v
bethhAffoG/w8Mda5MR8jtN3IHiM1DQ0Cadv5mpzWiZbqV7Tdh5nXZKq9oncSV6Z
mtFNAsSyQJcigczmgo8pbknzUyJqYwSGvVxh4eeCmkA32TjDK3xsjEQnELQGIwRa
kj/k7DkpeULgc2vlyo5guppz8UWXWjHPmLlfqUsxeV69mh5zzjPtcRq8xL9h8ZuW
am6uTF4FuA3s2Ccn5U9hivxqGDNGHXTbGyBnfrP/LfDo4J83lU3uZqW7w5ch+6td
CsjtxMwB9cyj0TZTdLgLVvJjYRtiW06Shpg7OR79gcEz+yjxrpXmtjyEH3NuPHwj
CeNNio3moqX0ZznEAB4KeUqv1VYqeAJux3PR7URiajJH+axakLwbJMcc34VVZe2t
C2i//jS2ho2UXmQLz4AXF8WwyGFUe2CMjh2MtvG7ryJcfBCsO9TbfL2QRJLhIzSa
J0rEFWFEZJFcHun1eFxa8cNKX2pLr3OH+dsX6Cabfb9qHtFJPVtSVlcXdhSgcQ1E
Be2vtPqGiVggWBXavnnWZnC9sBEShvOUkHZl6+V1WkfQK0tx0DUW//7MmTZZTtgT
GCnLc0tDkW6uWLxsjZXPLxEoKEpqib7XQuxs/+m6OGEbomvXNuodrXhIrQUkFIWI
z420ryejltZsKk23BIjBzkModSvwF2augHXsbddOiEjK0IS7WTTK99mlICXeZp/6
J8Pxa7XxZpfd9WrGQ0N7xCN6TYM7Rdgf01GuIrIp2vHHC+A4APxHxiCzivZcpaQG
MRKELsyG9lBktooqDX/iITAAyagQNsjM0mQiFJZymVRlwCAyXeIFsZdxk4quDgej
bl+R91CsCg/s5+IyTaqba36KVn5YD8DaDiXa763UgqrpNO4+oe4Q6G/Meytixmdc
iSzNbre2Y3F1ZO6QL9F5n/9T4sCRzIk30wYk382rXm2L5lRBwWfPFZH7LsqnmlX5
t5YMZe2pzs+s45vncg6/NVpKpyFUGpBEgb/9Yz5YeKXgkre1CiEA2rMo1SzwjnDu
07jvWp3DYzZSAG++6jFKa4N6lO+SzQ1ip3NXXwCsqRLVObULbabbF1ZYybOGPxVB
OAnGe9sRuA6j6VvMni5jm4Jg0p5b/uOF/zFER4j0m1IzWnD0rt45t9c8tq2Thdqn
xAezsjZZEA7F2IPw9m3YDORNsjEgaJ4PnvskXwrV+TRk0knIsEq3bNviK7T7qX/H
+OqnQGNF1tRx4h305Xov5me07PRN9W22de92AC6lPzPYTXts5M4Qm5YnELjo45Ik
nD+BR6XVr/7fB08jEdxj9qYHCjgGayWE8xsyshBgXEB6PlIvLjml9GN+ZBB4Cm0w
F1yvonsYpkxfkAXsWPqX75NoZHNRIMhkTfoBaN18kR52xd7vySZkvhqrPW4mnruO
FiktIC85ITLwI2fEBUKCBwC+WPuLOoNnangOB20r7D2iOO3AEjGZtBD2PBkKDPUV
Mm3Xg+klYunbeRAlw7jBWHV8YVbdgCfgHXBIMka3kIVPAa8U/ua2DDmPJr2sH2jS
/dapx3hpUq//jMlap3RpL56bWTP8VI8QsdOiDFDJWPXcn+CdA5I5t8mfXPSCzGO3
MJWVNy7eJRXPZ/AUiawve/zQ0bZ7QSR47HjSy6W180oHbd+QwjlFZt9aL71nEuq8
p8eSTQUuXUFX2tKzKDVCQAt/7NHDwf6zecFZtD+rN1nOF487jG7VwpkkfAaR8OQP
oXBTBcOYmY4j/ErmpN62Hx8hZoERY6jbPa2XiErhSShfLBATaO12MS+wT4uPKtfH
BqtMx+R9I9BPkqZQFlcXKfuzcas7/ARhUfwma6TOl8CiqQekT8jMT7hv+S/r8cwo
dB+lgFV6ob8OhftfiWfBchNV9gtc0lQ0Io6wTKHXK3Fo+u1H45CZkGg9ScZSkgjX
g4w2nNhQKBJzi8hvR3pdLTkGq8W712RykPLzA7jz0iGIEeSawQirAPez8e7Kr5SV
LLNB50Y+5/q87vxkDKpJoChM8Gi+H4uEGEDhi1PWiUSl5WGVc+Y0ce06ZUOYSNnB
hkotgq/E6/+whnVdgo9Hx3lfDIHPFb3lTfzmx+hw2mxpQsakrqIM8L/QwmLAZIjN
7SLLiHtjwfCUMnX/TUilLWn/2+yOXrg3YCIZcPozs7ROgSGVENx6Czl7cI71QBIw
IsLFxCCbx6Ur0Iq/c3iN2U3VsSZdxjFCpKA6Zdj7hcf0U1w6MEZSJ+hotasyB2OV
3nH6AqS+WUQtrrN1m/4DyuSHSY0n2bSnQ5lO3Ixx+47ElqdI2qKkWe2chXyRCtRE
9vYpBWLZFeShPU6wSm6bUX1picq2QfED/78HDx5uLwmYqlY0R6p/uyyovQ1QtVIA
6h2zuZnqLnWoxbEaau91mbbBOKNQSe+SQArpEGYS0NFZ4UApVqNsi68r5Eh0pImj
hqBRfmc3n8cSoOB0D62F0cjH56DNgncQsldxHC5PPo88DFLgOvBsBqvIho7v9RgX
sNWkWHyhP5u2EaA5SugbYOu3EQ8emTeDeDYWcSJmvqbvOlLv0bm7TH+K5lRWpjRF
Fs1UBQQGQaON/7JPKRnLqVItJA/ffk0Qu/9MD+c6Wh8x88BEz1ivXq+WUw23c/Ej
dVqU/oemk8geiv+uKT2h4bCMQ6Sp1eWCYebGe/PfGnv92JLvDzEaIapmdZsueMxA
AqI6X80obiLjDWZ1B1jE4Dvonr0j2GtC18g5077N15N9R3TTKmMaIVioQOxg8R1e
qIJ0erkhpxsSahozNIw9K7LlwY82HJIVxwknJU5j1aO2dc9YMm/ChibiYBS4r7xr
3w1HqreQHWcSC/h/ToINxdACb2bhXV1ilQhapjltSjufgaYU3NYz+bi3woZmc7Pb
A0xBWBJ/Du0sg0Wk+/gZn/LZTGqM//K6fSpEXiod43BF9t6FN7rxb9G9UMffqris
ONM2r5Fcb/xRsOKkiuxAo+H5JsDVMIzAvNpKIIgvkYi8etdekBtvdoD4eLpH0tso
VvgLU825YVH4glfv4PqOYyVdbasypNHBMKkBWHJ+S/23iI6u0jUm6dn8vuNFzE9J
V6jU+KzD90wvsFdrRxyyjDcdI5He+Mkx+gRbcy4kPPVv7582TvyK60GHcxmbbLO4
s11ue11m0NjHuJ68jas0o2KPODYjJY5IFtZj4PMV79RdTv8B9skfTHgpJH//1AM/
4GAYj2uJyQI7M7hrwNyY2fv8T6K3j6iM/WbLztFfDZYz8Q5YITuMoyIkKBbJI6OU
Doh6W8HaqPF9c9zxGVGKwfu1R0IM/ZrFt9CgIo0laRjxkIoai1YnwpoOstfYun20
X4KKngc73b6ypdfarYOSnNzFmeZiggvm6oT6Cws91f08WgjRzUiTqMT7ThyrRQdY
9m1/FrayXUjp1/CUY3ddVxJP/YJratERP2m2EYpsbKMX6hZMbn8oyfhXo8iqp5IH
1rmJlKcqgr4AnIoVsC5OCyvyrGPWl0RdZcGx9HOBcqhHLfzKdl7fYR/faHh3/O73
vajW1RDkE7d8L8u0mrnQcVKXefJZVWI2WjHn73E4tsXM3mIW+KxSD3rP/f03tS7Q
aOa5iVmQuzidt0QZiYT4a6fT8KxP01HhhMS883p1VPQhAUJ66aZYYpxEndyIcPio
xF8ICZkzoiKGgUuM++VfFaBgvZhMPKyOd6jqYpp9UeA0023/cnaIbs+4dkFwkj7N
3kto3kKcul50Kby1FDeY8BKf2zpSTKwP2UjBvwKGaN+HRkGw1UPZsHxW+AQ5TiW+
1oZ9u2n0sI6fyPSHlKBmcvJub6aijb8W8LgaAX8i8nTJVDDjzSFGPeYfL1DSVK7z
hC7Z/P/6ARGxXyFmut8Z3FIB2Ub8+JE7GoGDXEnVdDtVZUsyoE5RNMy56K5/bGLF
EiyT18t6sGnn1scjGT2PeLWXJsWR+z3j9CQzUx2+Gera9te+fm6zemUkYykNyYWB
6I3OsnhrRFWbmuVONUaiF8sP1toKLaSbSeFTB7bHW3jGCSZddOdMhZavl25WbgxM
PfJ4Z4mPXePbjRyeLdm5LAxJI9is4rz+Ju8Tusmt9B/CrTW6kp8c+j7MkLsW7XmX
TJQXZDQIGkhCItmScmy7wvRj2jo1VJb1j9z6BdpGdyZtgaY4mmxxnuNHJrIYnYQe
01J3gjIqxusYwZ7/UiTz/8UFx+EdnMB3HH8lp4RcCRWS5B66+WliC33jaxllkt8M
chMxPkTfLrhlWhKKDEHaPJBOOkrSOGbUapLIa9mJR6EVUlTI7pM4CHs7oShiBH/3
x0RXxn0Glzhnpt7JD65YUfX7kcYplBP9hQs9ws4CrSM25pFjfer8YqOmL69pHKHB
xgUzhZ8Ca8CUQZHCLvHZIGfjuBwL/QyQhkamS81CbPHmSJbsO1bIdvdxMRVBzIZM
ShW8i2eVjVS3ohdYYuIo/21RzpU3UimOips+cdr69xq/+MiaxVir3uM49sTQP/tM
DG2M0n+9r+JbjlN5PwAck35KnK1TW4CUbR9mJf6uqKGRxnoyCJV0jC0EfsXJu+ZX
nINspCKBLvsu1cxtBjK7k3FIF/Oe5A1pab4p54UmKDw2qstrGy7At6O1KBudySzM
TIOM6F1u9W7g4Y+ec8ZQXIavZKQwOJBFkxCsouLdh1/lp0m65CZG2bcE842Hn8+S
4tSrNjnuwkZMXM5/Imv5RktbBH8F1hvHN6FZZQF4ZxpgSUnij3jhZwRAYJ3czzGU
9qWRLYVgBmqJhcMMly3f4zwLgmoiWfx0vZx6hftz3VAJ7NMofsFPRPCAh/9FpVHB
tNoQrbVB7/wS59l3DuYe2l2+vvdwyDrssq19jdqVXKHP049N01O/ZYUpJs/HeTTu
Dgs+Bp6E70IMunQEHru6oJ8X3FkM4P6lGvMb+z7p5ZCmO23cFrOUvbR2BEO1Y1dq
Q7OodDBkwmjQTgSctTFzFveymZjZmdUp8yt8ZMnKHiaeVUd2OVTDc5YG7ak3e6oo
BUNzrfiqoR8daiTDG2d8WC5qOOGx8cTIUtYbfU5PWR6ELW+ObKrL2SYiBEkg2Pog
Y6wd3QAUicpK4Cb0L0+iI7DOo7sFYG9UyL7MoJuSZs2fmNLuFyQ6hXJYiW6Tf6E6
TpmQya8YaU1KD4vy7X9zXgmV0slVsw84ZoMqJm8xpMgDxhclPleffWdYPvKqRMVw
p6UsHQbIxp5Sz14JoEtvEjNLgIZWP5VeDwGXbkr8Gt0qRV8NKZpwY8GRTZYMV78m
oEaiAl+hVRp+ZRSpydZto3dWgx4Y2poYnZP4tPhZYm0B2U3skWJ6vpmeOeEEUBcl
LyisJIIYUpCbLKE0EF4/6v0Z5qEVKaGQx8addT32dSymUmgW0XRwgRsm4pezwi4P
ruH1SR9l3D6dqUE6A2D+eHk5lt4xl3pUHXGg+PbYQ5eUYFscPorADqQ3WJgMBDrp
GjXUO9F+nERCLnXPq1ZnrxfH418tEl01jVrmpcSNonT0pQfcGslz3DWEaQBdjPhi
vtQvKF4vY2Ps0xyZO6KfV1xaf6JIP2HVRiuwM8tGrvkVIczJ6Rpje6pZx3z8KPld
A6JM2ggyPoWIQsRO320pbEHh/PBgedDslm6F0QIe+wpXCYpH/j91K3PSxY2YjbXc
Z7TVjNlIv/dv9Rx63ITyQXrUoU7PLVDLxSFN4OG+9WVneEjMXyoeg3F5wdX8u+hf
7ph0zLtNgCTAzbFNk5UqqdB8rAZrzSfznSxZYquTCn/XTRvXixHPr11jc/tbaoVg
6nfV5w0S+aYVZnDHDEjsAXwhNj01mo7pT529nndWBSCygt+LREoTctekSYiPk4xd
i0znTxwUJkOro0H0ln4Qhz4PaiQb+ivJ653Zk/Vb7kV/OLKSHRLGZcYtH6TMimEI
50EmqSoFAU+03DZtFm8P9JbRE46oyWRRqpRO+6lpRfAygzURLXUOcTr5YSxwmksd
Yf1j2IFjTRtkweFxnsQ0djzSHwLBId1g7MrqcbzXsY/iGouVbomu1rXn5BAncDj5
7kc/HZQMvclAwySZkpZNzdGtscEsZ5fapo/ajcJPkNcQAt3Q9sqlK0xoHl0ozxyC
/5nxTlWfMOtyL6B5IuttHeFteN7R/m9A8YhFVjVW4LRgsX7libKLT/LQY8gr9vB7
a8zQmlVEPWylPrLIeFD05HS478tW+/mMvrjva3ypVrFcyYFu1PXQ6+b7Q0k7EiQg
1/yCpntzvtmTjD/n2zoKFo35CiQrQodKWLPeem4LVoNf4a24SEbjk4+KPobcUE8Y
0V19QmNrXSrxCguqhcJgm8iiGLnWa3rYYvIlI4rVizGHelhxKxB8kgiZ2P57oX9B
2TwIWJFUeoRXZgPRwPc6il6z6pZSsyBoHrsUd3ENhmrbIQEToxshsLjfNUAv28ig
g01eeDZ7qGnBC+aUxwX7KvwqCOg8NzBUmr7fxEcSv8mBkpcVOOprQ2aVTEDtVD6g
3lSz0o7PrKFVyiknUEJf/q94O01XKIRuzzcQ6m/DKuYJLJHWHjE24knz+z/FcPMH
YKK/dV5c5hmUZSc4atl9Z8M0dx/HqQz3FRKNVHh5vPQaEMP9Zy7TtBbxvhnPT34T
mKZdI8T3xrYfm+nabSDupM8HZ7wjv0d0CWJR4WejJ39edzOwssScfRJ/XyFSsvl0
fBUmjovfz/28h4gRkMkpfayA9OSuFN+qKvY09iXDL68YazLhbRY8dKDZhdz8rhZr
9EXpnNeK/sxbBuBfakFg4/XGZAMMflYBl7+6Hl/nReEvIta7sVMhk5scR8YFbm0e
p8uoz48/KFGi8/BXylpUtc7cvEe1lGvhwoBd1PKktfMawxYMSPcM9xWBXU6LanFK
9i4Tg4R57WoiirrbNHyEsLgbD2y2kgHyZhLHvYixAC4PB5hKh5W8aCgG/twArgpt
BPBi46jX0tDlldEMB0z77F6sFIsFwfBfGD1RkMFwf74sh+1Vg2d6dyUpXvHrHseN
WtCeY1OLelb8TMglkAdeda5fmJZXbepCH1XEf28fKOAwU+Vp4oCzcV44hMXLPt8X
nrhMUwSj0ssTUU/LY7HNMRZegNeHCsigfgSDdHrY/RN298jwzSiLinHbyHbHSA+Q
B4PDpK5xrdajjIgv5pnJFHxsB9zAgEVbuk21RH13ex9MZARsetZLndO7b3YGN5GM
OLYx616Hz/spnQY8lgy1gHkC36/uadOkJ9aKfIrib26iyY8ZaQ6EA4pL5R7Os3SZ
N2dJv13tIfkYF4p4VuhnPAMByANR2VNq4wMiLvTaJvIsswERsNhFTub0gJjJVUHt
Qn9QqmDAgUSzIus/Qj9JxeA/Yj++ad5iUoSjP+UDQTIG7ygr4xTtv77Yq4KHhDq1
Gdz1KGXdEhPeFF2S/IMUw6pWEJ7kcc44DjHIEGcdDINqcM5+scjBvf+hk2zaxjF+
cU7RYPBQAQ28lwR4ogffZmq/c0H9nPoIReXI+IP2wHrF9LtrqnGu40iqLmAS4K4S
pa9tILT+6J+99J0N5/qF+2+VgeS7rpSfJAnaMtKj5Mb14eaZkfDLEiV2i71/UhfA
+S7ajabrmoUgefL2SzZVGuJx++fWd+gjNkK0UcJAAVHq6UbE4HflBhqxPaC8CSq1
n+y1oWCfzPLM4W0lzsOOl+JGa7Oi6Ywmjl36MuPtUuHK+JXX4tm42/npG95Kvfu5
Not99FZ5Y/ro1vNlbvpLxnPwPOEcbJHB8GzuZWibqBjNLLM308s3sv5d7ud0cA0j
UHrt8Lux5LnaSvxjnPoAuZMKxPkbFjuOjw1FOJ4okQMMkjv5a82NlIO18jyVPj0h
OlERG5EZped91+UHrk9YUTUZX0J2QP+l9OlScET3/QUwsGhdydpxFNsK60LCrlaV
6T9yr2S8DHG5qEhYTBLkYNTa8DrRetE3taxZyW9Hq5B8A3bxalHFJOzjzUUIwbLu
T9QJ/KR+wDvlG5pOq+M+XArXtz1JUg+u7Fes2j81pIBVSsKoyeyK10lyv9eWVOLH
JEvH6vl9zbDeBqCrKjDCqDvZIrXxhyQ/fJlWNFF1YHMbMaKSWTbXuGBrO2HRuP/U
kV1cbueQz8KhfCRu1O5njzBBFx6qeVN7KtHoH02Fv1P/YQ7o0KfKYk9RDlqUlhH4
8h6PW+54PrV/dmNzOSf08E8w03Zpc6VzVe1kc08whtsFZl9dnmKxRtwpmcfdz38u
7seuPU3XvpbRPwT/gG6hWuO1giTPNlLfnt9yXwWgFllyJqLt5SW7jWoHwzFWt6ho
1Vi713aFf8aMfVyIdRqeQfobXUu4Fumtt1ocE5o+EjWLgkNXGkOggicru3oPo6EL
wtsJhHf5vNErKvWNzaXn04ReU5LnUwmFEAIyW67i/zVTB3HNTZ2Yw0FJYXjHf4vb
7/PDm4CL9u/FkaatN+bq7YzB+/KqrKvIwKOLhyfkFWmEHF62007DyBZFOsUjZ0HX
qogU2Cq72IXArROgAsMx10vnd9DIbXF0hHotB+wJXSy9uW2xCMazjOHE9Pd17Lxm
eek2RbiaJkYDunNoSoP7IoUTu6nsg5yN4PUuizSGhkpXBxIi7HfRb1K0qzqrMFKM
Rqe/cGvPpXFKTg3pA3wNyg2viIhsluwVrH+rVojt7vUqYEwja8wc/r9joVcoABhi
LCzoxj8mMyNBVqoVLPlbdPM7XyffBs1Nk1pYdgAnuuOdcbThKAKLLZDUg0aHQOko
ScAwo64OqV8lnCFWS2wXcb66/cPhgZviSY/SaisSjT+wltWsxvxJGi5P8KEVdziQ
kGItaSx5J3A+Yps5tQ/auNAdnNOomFnSttPaByIv6qkdTFUcy/wwZRzsZdAx5g1s
rxDNMGWBO4/PEO4/YJghD7RoHyTOGW7CTIYc15zaklbsO0iU6lm7R23JsM7Z3Zrb
vuGysc+2+E+gPU9KwVlr5Kzrba2ly7h/Ms369B39iUJ+JIK4RcuK1vTs1xNjjqme
LWra1/VVa8woYW0WfrwaO4wv56CTcBQGIi2NPAIUgDyYbZQoFrjwZOU42W5803K+
OuObeL8/7xBi5AOqdIpJKMiLqo1BaLrCN+pJperunmSN7iG+uItjpT8DY0u8lJW1
NRlK9Nzg6yKFgAoAk5K5Hr1sNe9wOlZiZXyhYm5ywxyQS6QS17xKHrjKgpfEKDvB
wONxdDKQdH7IHoqKqjgx99Oj5gp7NcSVSG1O3FcHPkkGehKylS8603+469RudYhk
bxweOwfQ9nJ2VqvuGKfiKulr/3gBRdK166meJAI4qqYVeIjlywGmNGdpm7sdgjlO
E9XeZZJbHG9XJ2s5s4Bo7mR5J1ep+y4qd/AGygaWV3gxM3BpbWvuYWascXY7DQm5
bulL1/OUKvGL+O64j31GFOlqj/V2TmN0JSAe1sXcd97r13vSHfwZfozqUjUk2ER9
nIDPzj/GyPTLrhJXKkfJA7fqxb1wpN57QCj+AZbHVyXYUDGp7Ij4TautPI4xk+TL
HVSxzSkB4fgtSG+HRT//CsjXnhcpimR4Vf//VZ85OK9GeO9iHglZmDd34+MnSjF7
8lLUjG6C1ymcgkFD7NP3naZGtt8GJQLMKqOkOmGgpfgePThhk0+AJfX4iZ9wv9cf
bE16V8AsTymSil0+uO+V4p0bmgJP9jS3QTYOWFUZMFKO8OZC0tEuzFOaD9urDXD4
Qv0lbs4BHvOKnKOEIe1TYNTMmbqs7hU/I4hsF1VOU+lFD1ehR73hgcYa+EJ8VYgG
2qawj5EBnTOMrSzBvxjpPb9DNs5/hh/QZjg+frU1wc+5S7LWBQ077fPGAY1G4JQ5
fGtVGq2KeLGp/hb5SpVRXncycQGXXPvNZfDN5QntW8mEA4gg7moZgM2a6hZgBRRi
oI5pqIbY3/deA4Y//MVXwR0I69VLF43Vgjy7IKlWOGolP+XhAdxZZ0ptB0eJo/fL
B+n/ejh14JhYQygvSY8CodxOwcDKuPS2oaKMwoUKD/6i0rXhkRqNalZV4NzXdjvU
C0633c9AsM8/zFBODBVvERY5EMQhDzCUciFO0bSdSqNGvEBGEbk0AtYKh252cjq1
eYjhDAZtpAHuzkY0sc2y3mD8f3TFqIfyJFtcohsIypwq1oqXqUgrh44ze961I3Fc
25xYO4Reh87thG/z7G6joGMB9zCJi4Jk8fJKgeQfcsdlO2GxaU95MbAxsk4Ng69y
QcmN9bhbL/WvvFnTWj4GFDkL3XFj3w9kZ1vmw/rXANKYClesLiL/EqPzcKctCj2A
0JNbQBlnbzyn9CLG460U7oQ+5LV723FT50Vdk5AnFKQT+p3/7xxj7Pqj1CpfXPDM
ej0n5Dvc3vsxZIgDuQo9vnf1tg+QtL7/Fuoj1Ap/HJR/ifBq/UqzqCS3ejADMLcL
FmUDlU6JvLEgX7l7FIfbkqvRLzeB9V8HBmYCwCh6iAjoWaXo23rM2PygI/IlE8YI
litQE35FDKzNHq9gJWG6/44dahwVQ+HZ248v+PXkZMqTvWxMUCkwzgKswp2uzcPt
ckywdH+jRYPcO/g50uzfrC4m+8lew0YxEmHUXrSo4BUKS9dVtud2B7cv2y81h1JV
7yzEvmvoEUYjdIpzawjZlHo6lqeEmlDMdyJ/E5hSGCOj5Ny6VEQDMMV9NyC6CQnR
D4YHVk8SUpD2EUGATzPMWhz76RsDIVa+wumCFiwZQOvthWrHlL8gi2c+dcfIPq7z
OtZpGVzeWs7tkeZ/74j7jDv6g6C8+6ZwIXFfhhWtgE61XIfSiAdg+9VmyH6od8K/
PAo7l16X5KrqPUKyLcXeNn3DgC95p13j7g9xtDz76Sh7+8mBEppWor7VwqMT5edh
uW0xoPHawZJqIv5YD3lPhOotaGxZJDc1bttdmEmoEre7prDca0yZVjwhxPuZQJFM
tgHTYS6cU6gqd6Pv/9Be2YapTCPb5SJzvrvuokSBTogF0FZDyb5Mu/UmOuoG5a4z
XlRu432M27qv5+RXTdxVlU3veMwbFENlmBd3YYkfFOZxuicodVz0heYg4OSY4aOM
CS3vJBCPB/Z/GtHV8/pfOkfTc+zIUQ7NrbMLCnmd/Dt7HK4QU1KhpevSpWJWAhKH
RC/WcAOCV6va1sUMZt2cjkXBvRKK9g28LVZymkV79e7LCpmQoVxO2KtTHBSo4dcm
djjvGT3k0py13Z3BAx0OUVyfG5pDmpvK2C2Ayn8+59yV1np1VbJDr/M/pDBI6ajd
BR45acghXDK05FBhXtrx39Dg6M+b5O6tPoPfi6YgO+JgfC8rvi4LsRVmqigTOqKz
T0G0WadBzQWvka8GBZecAwtNG1pagDRPiqbhjm4uJ/9JL1/vmPspVoMQC6FnwlJt
6haTfJJReUxQhaa4oF8QcVhwUoozl0wh9vciGldmoq4XptIL0CVOeM4cVuwerPI5
BThH1dm5eVLLlP/5vevo1U7eiwtYVkmHQduLvA+yK3s+BcsmT7zO6Ldz0Gs5Eldq
6a7Ab2/ekTKpxcSFp2sysdSUhrgk2t/4q+LLIhCXhpvi5dNjjJzJSnVNPcnaLdAV
3RtqXnZXcMK3+RCbrni4YOyUgy1Yd/9o7GwC0KEKevbv/e5+oSU/OSk7QOFlst4d
UnkMFF3xdSK4Zy1e4AVfPOnPwxHCr8pFx6W88RkEiXS/KnlkDi1izmHMEuN5CVW8
DJQYUHth9ZXVE4m4FFYkq+/DruMXaLQLcr05oOxHEsGmxdK/22TNGmu9x0nv3WS2
1fQXT/+pV0jSprfMknUqMzycBDTuXvZdCFKU7ZnPHq3hajx/l9OnjHOAHEqjjbmG
CgDEcpgDZGZrqmbrl22Fkd/v7uKqMtgwAhcHG6zDRYinLFEdVGo+BCQDJpHJuSDW
0TpO1vGMCHg0/nTO9S7KUBx0FO/ndHp0RWzZwOaBrXyUGE9RQc1UHYh44W2N2mNx
0rJ9wLGn2IL2cV1dHFkLOjL7Du+wKO7fuYVD/sKFrJVOmvWMem7404OQev6zxS14
2UEpYGszL6Hg/yWpCxyf7l1fe1NTGmeYDsuCf+IrmsK7p5ty7xVNc7I0IF4S4no/
Ik3t1/aDs7d8giHddvrlDUNz527vOtDzVGXFo8YrqYW8bt5vt1oxWdbSoZHHgZW7
Z1LJfe9MuSwkz78N1vurqbIVwrxEqghakk3JQOeZIsYm+XiA+YJKFXkPZbxubs5x
X2mhNmdD4X+uQskQ9DkKSUFkDo9nlTiF9+lpU6119Tx37mxk1ZCL25xPV6WdnP+e
RueBKo4B4ASvRgGxxlDWxLykqAr3pWgVvUbKWVAZY/Pnbog7aX9mOG0dLDwF+iDO
wtSuXGXtHNWZH1M4xbMZw0sh7/udQiE7SwVnfUz+9j7Q4bOcSMBCFIPpcHsumXWI
EIsXR1XNeBEmRTmJ0q9cj879ML/ntOOmXgUm/CbUfhdXaI2aSxAM6e6Qc6fVZIlf
0kox64dix1jwZWInaH4uhOZufCYDFU55hCyGyyt8faGsc9KXXTXySDZwFKwAA38F
1ersXSC6OJG49+XTAYfQrlvnQWObTS/iDUjXWIrMY8HZncak+WjHUu3souEOrD+Z
K/oluApiRGVcyz8KRRjgtwydHhi+rQXqM23kv1zKAU6VplZCCGpnKezeM6o5RrvH
WMQuwXighQkSpK/8eSEFgbG8HsVvE0ltD0mFWNO45AYfZ+ynk4akeA6bdXG9tlam
PAAegGq/8l3Lo5rl1OagpySYV3QEtzvIkI4gZDbLdg3GjAMhYfqbJ6N/NCapxfPB
IXvCmh2Xgh+QXeyyVla+ARAwPN8qfSMP9ZeDcLZYmiQz5VJcQlvV5BlBXtWyjPeN
TBrIupegGCIVQCKHtfiXWdoGjVKbxuQm/5SzPqMOIg+Mr005iRh7aXf7pYRw2rHi
lV+MrIRfz8yZ31xNOaZUcmPX97vyGVMw4jKCd9thts/P9NKcaqffXkYPvBdNwnfF
WS3nKVb86E6mcKnoTroLZbSr2mGI58ZDSmOuqK3Hfiu37Yub2TLTCL7+MAaLN2JA
7AvoxRWl2EMzc47CKCM+37xUctFpGZcz/UwNgfkhcJ++zuIviDB0bnMPtgv4ZWs4
1iAmb2jGzGC5CYI+Pkx+Xb6KY5tDhBXWRB+3/qfngqYIAcTyCeqt68mldixrqKaz
p7PDto8Yoonn94+QBzKajAnqbxBRVPaSYKA3VIg5YE70W8ZUtb3MFsdTtT4ZRcWS
Bew/oWL3TzUnLGKKE5kOh1VZRWA4VWrExUbKniNUGwaDQot+NlFbqKuDs7VhDNZX
4gtAOi7UZu5OGSMXgqbJxLA9NB5oTsLtueJ45BEC5TpaTQCGL5YU7+lx/1MDJjlz
u50qzXtPJPORLwZ1Sttsttyzd1D7YxIcrW3UsMY/dJYatLCIuJCcuWtOd/ItuFD6
tZMdyF6S4s0oulVKESE0HDnLZI/koHw+lDHQKatm3k+SRa7zoFVcy5oc8c779/Pz
9KsZ/Ra5ud2uA+XuW1rJF2CRgKI/PshXvTYg8E178EwB+WKZfSRh8Hzhs5q/iOif
JCWL4lK18dvg4Lmqeiz3UHGFzZrwMRrDECqLreXGKZtEr7wFicLddE3BTeiOopmX
3wg8e1GICkbufQUY3YzQGUT1t+1nVtg6/xqB5FXP3SN6eu6+3hbINIj9xCfjHkGH
dLMIRDrD5P95h20TMFDMClylPXBoYcpWaHvE01n0TzdA6jmdVt7qxMgOd9af5D7l
5X031IuvxTQkKvrzFrP1lqLtGoVBnCQh45W+S8YkAydjqnUK8II5URe+8iO+geCv
cElrgCpSr7wMuejv2Ge0CSnaeb/4ljsTMt/Ex1b/TOYzpBBvDVkugX4WBglgBFH1
I72Kc3JVPTiArFYepnZXbjcSa4KK6GYxhLZWXQzjYGwKfOBq2SvCK+8pjUlRH/5T
EGkN/5iT/ewOh+8PL7bSly/jCaY7jacK8vzH2LuIqWxRRbgt+ZQMdiD/r2pXWEOZ
+Onag+3tLa+YXpQshwW/R6K/ycgo6c52uRVPArgH4YHcTo+t/REMOpj3qCTlNXrA
CO1X6ZRgCSb71uYh6hDmPichGrMqU0zynE88xfs1sjQDDljOA/05qp2p4EMbFvmG
Qod3kZD9UpoyY/F0g2Ce38BN+zDCqXAo68rl53JzPkTNqLSfuM5oSIZ1BrObCIVQ
BHcFPKcc8snM3IL/Bn5M0yN41VksCc9NXg25HPDW7rp34+NejrfAWbBuPSGYzISp
Y448dJGsGI8VhbgQyaPOIuudCxlJCGq/qkoWBFPwPGwOI8mix/1i4gxO85LlywpD
hlXNOwB3n9/CoAiEzA+F6bs7Pw58gPWtcUtrREtXJhfcOsIodc8CGPCQs+pga6Lj
LvQVzDPIspElmS1Ul5bLXcB0a5vqyv8IHUpSj8xf4KkgNKtOP/YroTSs7mRlx5cR
y9R3yKb3ZlwFlDhSRvozkQosfV/ytpraHBn2V0+OUoxdBaG9i94DjzFF2qMAYZPv
Rat78exI0a+muEUbOS86aSyO7tEitVnSUlnUDTQeN3vYU8ywwucfNc9xlnUJpK3G
TBLOf68xqheRx7yFSPpkIYPtO31gePzd/1xKQyHkLpdpSPlmCLYOig/rJQx1B7st
hNx0IuN3F1xeibyjnqNQvSPHqKC/cMCYqj28OgB5EmQSgYEeRnBF4jzmGPWP/yuI
s07+HOvj6zRPGGEbJIsNASTaW8XL5bgOTdZPB2VdDE8Oole9MNGk+zmpXfBlwt5a
fOrAx5/YXgqgRYh47A+fNIRkl+adQZ3M+TTLuy/eLbzmnG4yk4q5gEqv8aYFqTxY
OVr4RjP4GT8ETjLOnG17pHTgBNXL4jZuc3gbryYNigO26klY7G/8yZWQaK/GgM6e
ubYqgTE+dPZHmztjDm2VcHTn7jSnrMPlAwBoooq9P7GVkKpDWKylQaUo84HaXzbN
oeUjBhTIIMdSBV54Z6/maX+Zk1I0t8aJuEayIYmYk0pgUxrQHYcaDzNnPMhnnL/q
UiOFWU2/UflHeKDRyXPvK5tvQHidnQ+kFGjmtjpZD44X7Pki+j/vj3skhu9VZnww
v5z2EoZ1Nb2MarRhPjcPFNAsGxj/sUigJVd+bHr5J6KJqkS5Ml6wr/YRqm5jATvz
WTuZwoldvCdgClfYbIma9fZPmbPzf3T4h/O1W4RcntpV1l4+tJORIPN8JTi8SOZI
DC2rtEtLi4zizjqxDv/0dPkdyFvJI7LJZRj4AYsbDxTFqvVQNQF8MLqEkIa9g2do
sWpYtTb0tLFO9YQ1HUzwOs/uBBK//e+dnp/3+Qbcb6bA6Ax7pFhmWJ4NwRTFPLiZ
iwBwypTjowmKOLi8+AYGE3ii1/4DN8ZVuyW4OznAqwU8urH5v3GvdkZFmxHfilrt
2nHCufPKZ0ulp0Avm7PV3mlVxasi9S5VJZsBoqirlp/8NA/oQW2WZQgNpDdi+Zup
WzQDxfNja1saVEpiNmvHsQTXi3S/kl8XxaUTnRIkgLSsgM3ZKaqWPOJmxOCABsJs
qZKNTm0A6Bd3f48v4N7vG1If1eTx7ZnKJ39AR2BDvvcCnYfCp4GrU3RpxkUdZzkC
aq7ZQlNRkhUbXTZQyQBZCHrErE1TMbF/vCa6MDkWZWXgCTBqkGRvNIMHE+I/7J9f
4eZdl1H0SCp5pCejytWAia31lbR+1bnQ8v71z5VOPEkXxK//k3PTNlR7qS9Ue2Gr
04HtvSPc8TJHS3SRJJK92uTeT2vXV0tguLnG4FfBjKB6YiXHJNehPZOUGfq30vmh
egoXPiTxGVNMsegqkYqsO5Cins4IwsTpMYbD6HbKVIpMEfCPv6aismmAvc1l8Z6q
I6u5k3Mnlx50qBoMs7p/IZo8O29CY8hWGky0jzoY78FAjLnYYNuwBogiwWGexYrW
HALD1ThcQoPEj7n3xRcQK4WG4X36a3zQLUAGpWJ2Y4e0M9/vlyy2ThaS+m+vA/qR
oB5e5ARaHCWKiQOARKOV9eKph4PpdgceSRralTu1waZSZ4AmDKSuC+wx7ETbMGVf
jLjQ783nVP1CZXAhj6Z89AuUi7gjucvbWm3Zb6FXP03SQTDom2pJX99c9AGX6Wuk
xoRzzX9sB2oq/IVRxaPIGP4ld8DDINet4unODwfViI/nDWpaT2iEGMePFX2JYY/e
sqgS603uXixawjYcNSry1PJzm7YLf1TLrES9QfpGS0pYVuT5r3jI0AgLnGgy1arR
TEASshWUdyvWKpztKj+JIMm2LE+kSI/enKzxTe880uR1wxhsIDcBX8t+BonLkvl1
bFNerJ4PmSc4BqXTG/7KeJ3T0icptCVDWJHAvyB1wrj0NphYWVTHCxDAVbhFfmX6
RO0vRQ8g1iZ/fIT5anQrRRu3qvHr0tujv6t44rFZznGUB9f16MeuoWrP9ndAS9Rw
GcPq3Cv2taUJh93hRjMm8WQPYj+0R235HA8rwKYsF2qSpIhs8X7/hhQNlPefi116
NqQnnuVe91Hv/Zu9XIAINverDHn7M3eqTvtgXCNpoecNRGvatIKm22JGmI0TsHAn
sHcK1EQCq/KYWJp/zEiUUmVcHEW+uR8O3XvdNEHnpTJZocTueu34iWas1CETxzDt
wkECSv7qBwWOOP2PCFKt7BjeDjK7HDcvraVi5qjMcTdQIzS3jFbJaqxbeqCLHrag
pYEtngOlDDuN5ll2BCIIfxNpnnsSJvRoUPCiFBZqoCwQiPCBCaVF7jeiukhiYc1P
iaK52/G6vLPQx43iFZAfq7+MP8IgcFx5aQ6K+PRQ6hW/3RVncjTD5zurwyseeCR/
kHJNai68TUHW7XRDeN7388OddZQ2oSuzQR8tpaMlqAur4kPqJCdNdQzZ78QyRSr8
HcKhzp8XQiZg8F3p30PfrPHx2Hs8AHeLKxS6AEzo3BtWuTckBv8GxTFkW0wmFcL4
lgbWQlpWlTeZy+skT7QREqiFsiNoHBV3zNAGKBKP3+TZ6LC7JeYgfHn1y+Oekp6l
FTlmRLBYZOSuA7VcfCRHCE5LlOrps1mvbmY/w/5onIAMxn+LRNqjnB5cv4dqaniu
tJWMrAGHGA1asPR9oy8zPU4fjCDUuEeA0bzEDurpMQOBbdrhoXsqu3oiNmiAZuh0
rNA0azTJ7l/HgjbYiHNuf67yRpWk2duXa87Ki1ozsj2jlIS3O9G6s/AwvFMgdO06
WH9zqHbK3jKhNHY19ftJtDciqxpohFH3AVld9UVZDKRZR1bVyC7bMau1W+ESGA4G
I+4uiatwrFr/daZJLj6c6Zg/vq3Z1A8d4wyjSMjkFqYOKwjR7oxQEAOviJBqTPjL
ZMsRiLb5TlsDo/f5JrYdaBbiePe21fRRfPcks+BuhkMT8XMShX3RzDCeFdaezKuJ
eMSxhQEA6LxsZZGNclDg9dt9PNA/CYb6jje89431u+DWw7IUvZWvYcuir1Rxvl10
qVFRHYV33IRlCr0ehJPZtUNNFcsj9th7gTCuy5NNq+qguULEO2zwnlpqRtJqiTRG
NLAI3hlnZBfyuDczWMikzmmLUAs3H05qJRaZPo7jQn3lolXKl+W2CM6ReOcy+KH+
JTlP+PmFaGSKQnBMdpZE0nJCieEiKLt+cnnEgyzAJuf/FPclR2x0LD14GE0s7wTV
XVw2iEuukgi0b5cVtyhzKdNQ0j6153kH7NQ7a7PQl27WnhRBozqCiCHh+O07mV94
ungl+cxRumuzRgYtvV4qHUhxDpPV7+4t/FvlHW/zI10zJwUfMT8V97Ao02BdT1+s
K4KVUL6Eg6u/NWvFT+qL9iU0X+wa/f1tSc27ksKM/JuCu/uH+OPbwZsz14hnt4Ge
vTL9MiMuUhFyVtYWLNhmKkGQBWgucgZsufBVOta2hl0J0yVpAPwjX6Ca+xjYoNCJ
fwKATD1A5zMfg/crnByKjS5QdS2znOMxJ4jQ5YzvLkES6/3M1rXMYC9XUESnH/j0
vjQsCw0p8CYiYVpdFFgsqU4G/tlGZBJobsisd1nt0rIefjAy9hA/D3dHR79KVcnk
VTCMEzfi967/JWYtsopJt/hm4N/R2Xm/Ky+QqJb8sH4MhG+VUsmblIwdEqE0hdYx
oCdvSTuZuEcBDmk8QiAuwU23aNptIuDegMeEaCKolHUiNiuYNIeiC6ThFGaovPEB
OdLCNlgsBRuw8JIyW72OcKGOsjd/6CMeWObiRCbjrDQtqcn2NS8dQKEr1+mu2rlk
zwxZpcwci2vEUwlNIATo6a6VF4GOE38Mio8tvz4ySIcEBJV3tXUXb29oM1EQflIQ
n9z4PtZduXjIL73zFKrVE2pPzbS/EscrFxKA50Fo/siUPQZfe+cdA8hdgGYKg8C9
aPIJm7aH9Srx6YHUznZwnod+TIp9dy5tFO9BFySs58vdv4Trd2TiZRiF8XzoXdbq
SRiqqih2uT7EJDwLHAyTXkMcHwFfuINcicGW1xB4mJZGfcM6hqqd9Xf4D1SUX3wr
cSU56ivzduke5Y6SMaNwQYCrginWloSCemZIkNfkFuifi0RlFPCQwlye7e83kP2z
o5DwX18SSKPaFO9JWwCq2HEnEwWkFi+Sg8NZth5Sjqj5N+GwpXn7+s8gREtSV03h
Vi8KbFy0S6X9jYAnMLUPNebultHBk8KeHWvh8M9R2brEHIyRMX6iQYgrXIpniwIk
v5IvLz7JClkUGusLvmj3NA/ni3gBPJz6qFXOFZVg5+6zLYvn42Nu8rjl6dvqgkhD
I1N8cATBqpNmbXuFXLR6bx16E4SqDrUQfpvFa5BXcBbMPfmW01hgcI/uqxOQDQPn
MfgFJhTH4Y9dvRr5DSF4xp8osB9kOANf1ZSu9BlmUCYJQuFT8S+ZzKfy1FDPq3UK
EmndvpavnYpZQj/MVO9UBAfkMHX4nGk9fCYf8yqDRv+gfOniNI/W1MGMMesbdrj6
dHvGGHPhlbe686+yDn/du+lNNJXAH4XgzJvm2k+BrWjoMrKyNlUESbzVVRCA65k/
BsdtuaFTT6ArDAs4fxJVWwebSfuUjtkM38Uvo1uslys2iMKSGTxKNSE08FCMYb54
5Fu8YWLTMp/z0kdcYd640EgMrEcSGHbZpifQNJ8O7GmzHC8F+kd2tm8xXmK8ZE/V
rE1j2+uoQKvr36RkYaPxBo8HhWkEoV/8Dy6dx9r0esfOFtuYs7i+PhYmEQp8xWr+
TitllM0Vn1pSG9+uevqiwaPXGqR9GGo/AQGjZO2pd57GHbZG3aavEBv8qe5zCoIC
psvfEb7EmPXTig9PwBUv4Nl1cQoQt00mY7YOtR7fWAZCvRUMl/1f2nQMmE1XJD9W
U9qun0PFw76WP14CGwgzAdUxnYNtPMr9dXDwIQUlzLUHYXVGHfTucwXRn8i/5vHT
pNWy9U/oz7XLlV7XNp9zCPuH4TlgzLAZqxpvYw8gnS1/C8O6jz3eB7ykS1HhVaye
oDMKUFjmytCSx50RPv1UIch4HX+07smAkaK3dccThW8173phZxxmB2L5UureWM2f
a0V+aUbIcHgXZEodXZiL8H9lwCQgdmP/E5skphTU3CtGcbXfTBF/Bql84DnyCOMZ
P12x6YiiYmYAkusZN1EcEKfxQcDaveV+SfrjcZXcng7nlaYL8y1AKN6jVTumpzvU
ePspF07JcTAjU6J4/GZzqcTntgTNhf8/NOu/XF1Tll3mcIpGSwsiqp+/3PG26Fs9
UHBOR+cxy2xBiew7wiZc+CHWOfRTA6e5ueyypcKiOehHM0Vdvw4PRKsI4LBbGD+D
c3GdwQiNwaQIe0v1uKfadjp4fzgK9+LOovv82PaSlO1+0b+5EQdyu2Ii7syzfYug
67LX23dgxX+hkwVFrPoiNLj9gI+OsABHyJhC5nh2vxlXMd9pBb/0WvWeA5aDZVX+
9Aht6rV73GzPKbUAfVphbCtcrB+3WyuAN/aQLLfGgsuYt3YNCu/o2Y42xVBSKn/i
wCm/IMmWLm2NzgoMGCgCcTsmKEpopYjD96+iDsvumBikuST9YIAqOQjBgtkdntZp
kXTzaVVQ1FPWG6H4oRdNHokI/Gm00z9Cc12Vex34TMmI4bkoyrB72ovJFdKIfEXj
0Q1ECj1bkY4dsrKKLDPmf7FOX5oPZIZxhTCy8D+3SRNXb5eg4o7kaSREypG6OHCH
Z9+kJIZrT8cyegSz29Oshygdw5iSpW6nE3L+qwX9EYwb8Um8PxZ7xFiGHQgoxcZj
EOibBdq7Y9HOTecb9wJc3HKkT34zillZauE9xjnXcwpXOBaokSiiGnnjVD87azs2
1x3TmFrg31qdChPyjGhfMpHA5bKRve+72b/fS0dOG96fCEVV1KslyLS6OT5fyCZi
WHVe3eXROJi8xP86TwRNpjwaU5bmrZ8lnhrt3y8d8S9/73/YJyvgC+mxlr531/Rq
4O98es/hmQtMuHiIgCt2lHEfzSrdv7U7es+/K9laCE3345VBEvdgXTzWJDjlzMAT
XGxojW2vQhJckniBUTz6sT+3KqmWyCIiLoL3iAJC7fZx+WqveZ77TypZL8NR2LYE
orkfCQeUW0ams9cqgWuF/YNT4lbB/FN/DP8Voy8ineTu6COGuZvEUXlChHgygnJy
GQYB1gj+TxPNsWd5AqvFZt2ghWCbspr5rbg785uRliuKMPenBDcQccuqdQAfTv3/
Imk4HE5x4Z+jtpXWLFD5oKOY3zhOy4SaKXaMIqfE6LzeCsWF4Ube2IqRq5gFjbZ4
+9cHDDaVCjfWl5djiqgH2aBuP83AUvQ0Ytqm+tGWjp3rSc9jjL33ZTO9c7fJFnt7
M83w0oL26xqsG+ZRZowzU7pZIsudcuCaV12oVRe+ZvTbeBZGRch1uimb1XdgF1tz
mLptkOFZKAyzR2tPNjKFmWQRC8JcbyamGrylk2MCHCrecCUrtRwS3cTYiSudUBYl
YyjuREF3U4dBMqAy4rfRp64chexpdE6P+9DLF8e9D9vB/wt35WvzPW6g9NERtvmH
QxWAWraEcHFN5PRrl0BL5GuFzaJYdGJVpOsz4XAwnedajb/bJOKDa7KgkHZemgHM
B8AuLKZHxq3xsXz6CU0rr7T0sqH1DRf5aN0Y/byaIg9fOeWDkdIWA1LRg9o671CV
iCSTcp/NvCil/D0nzPmdIVUYwr+tXEzI4X2VsHmRbaTFMzCoaidvyBPNzXBpbGIj
WYvJr02Z52BgD5rwn5Dr2dKoGwPmWBFGFQc2akHGTsmfLxldMTGBSgYZ+vk73sDD
h14vKjj4Bd3msZ25BOKGHAbxSCZDHC5QO24NdwO2EmgDXa4AQJndHwAd0gx5MdZ5
/2kTH5Yu/XELmS8BRcYxX9mXb8XCKsj7pOoGB/Ye9PWwXLof2bQ2vfAzrFxTd43l
Rr+TIP1jMHIkbQNLpe62T9ZCRHsACCYz6T+ouki3e3MQppOkfSKnvabKVRQZUYSJ
3Lwzk4I1P2FZQESNhIJAYwH47hyQ014tsQzrBhm4Yo01qASERJmM65akWVTIxFV7
i4VZisjkREUsFgndyHtynvPPua+DpVUfRg2lY/7z6qWc7/535yoOrqfukA1KMKfF
VEBmCTNPD6qixt0IVLJvPZwataz4QySHMGYvYn7X/sw4sT6E4SF7hvAgUchny2XL
W2/YeNN2Movwj0He6J0k+r4zMtKx/J8/b9uiVuOev9epvGYewiJk/lMc4nCUp4jP
7I80vTt3sBA2OsJ8/2CYYM57pE9MqMg8hG0Wyv1OTjZhJN0AGMU12oujbdtC8SsW
xvyjMxRgr7BsFqUJlfmuH/yC8Pah9dC+ZcCNHCgAoxU4o8UIE8SCpEmPqOl6stYK
kbpmNVn2KPtFs8qOqvXX+n8eZ8d9Yvecr/XNj73rYEKLOh6wGdLKxEko1Zrs0mjb
exIc1hIB0fqgK7g5/z4VHc1ddfjsMDo4X8bJK9J3GyKWpXbDuvyM+CDevUN4PlIz
EzWJYKDh1/06zzRGbrWD51qp9HYAMqZibUYQ8YIhAgmrhhbABAnPFrxz0HFMuCEO
fffZeuppvE+rThEiFxR+qwyO/llACSIL4+UZcdq+8lxdQTRNLt5iw4YPBfmKaefJ
Ry89bNYW3ZNbRb15GEVyh2I/KhmGbZU16kxJjL+DQYfUjhOU2rZLzj8Lw3dhYGZX
62UUQXbbwm5HjNtfutij9IiDsvxtzoeZ5m4FP2LUUwO52vOfgQxFSNWI2cEN1Dhg
AHApilH1SWAXEWZaRmN46AFABweZLV6FgBp/Yz70Wya6xZYjRcpZzPvsvDS5CmcR
7W4yr9K5EMtxK9/iUjrqb6oB8WLJJTGRw0AtHefLbTOq/h0dn/xUSHYZfcP9/2gq
ZoTx+c3HK/JOUu3EA3WyX6jRWyQSbNXbwvlZmFLZIoEAJcHL+gQlBdcSn5E2hx6c
ST1z3cZuXd/Qf8JyoyBHNgpQCo6h+7PGSgGl1L9Pn+mtcjzyYkcZjXlZPvQjG2b/
S9WqpNmdQo0iMBxooDj+bnaVwi27rXDDOYJ3L/xOYD8kko7PCAie06V3sO+j8q7l
C+xPiHIK7LYxgDHGgBAt2mJRnETZdtkkbXhV+Y1t8uBwrhWM6vCwCLekBvjc3PMC
k7uKeCCBvaG3ihOCeiWy240FC2XYHdzLui/5+0iM94qr66D2c066qkcGU2CW1dEr
/p2aHrlLzTjg5XuKuUJL8QyjNz4IvUantmCxjb7UAQQs6tW7v8BhpMzfjSievixf
gfSG+Dwc3C0tUNn0kRt93eZMaDukVjr1uVeVjvYWWK1YeI0ktk9fw61hjsOdacuO
A20N9fGoHxmNcXg4CfeRJN2ys/Zz6yEDXkYvIWv4nHj5/wPeIhkIe1u0vNtjtSdm
L4d4cWAJBJLYvwn4//2AEgifEwGuIPzSrVc8MhAFHF17mTCvv91hohPXsN/fRtfQ
Pq4p/V99JvDhZc4yAW8VgXFlRt6wuysqd3LOIbQQTpzWj3EJ/fapKo4ap1J4WjRx
DwX+O7aNxmr6NAMOVKlPpOIQU8lzOmAbaFiJlZePdjretEUytG/7cRgfV8OQU6iA
93sIcwtlyZu6C2IXTXFJ8bVH4L684msAt/yZEe/9sTdE8iIYtaEXPVgcfmno9xQO
iVpoDFM+1fnhTEhWRLOF1YBVxt9QwH2UyRT8+8fHmj5Gy30djnBOFfJcXixx8os0
vvyTBP68CEFHlNw+dgk1ksUljc6FFN/+5rA6e3myCezFvN9zKYDo0RqsDVWYtPLA
XwYQl81ukm35Hyr19/jUwNqRWTZJAkH73C6naH2dPV6yfQ7A3hotXE5jsCNGPSSx
x/bFzdHjFlKOpcjSFfzjJ9+GqfWiebOswXCTl3MdHHUc3yb7tx0cgLL681g+aeXL
uDhqmTHV2i3UCbbGeIRliwUtId+5DkyK1eKekNevkxJedJsDxE91uv+Dk4/qusLb
otQyPlFxz2MY1N0Ae8dXiSwAYeYQQVcsW0U4JDo6D7N/hRPzg9j9NHTAndavFqDa
WYmGotir5XIvK17cqz2pPzFVwEaB7ueCOFJq7GclzQBmkFtLlGwe1i6TqXdmhzhs
qDDPMiFKzyia1R+BIZYZFvoyqG2S9KlY5N545jyC+Uox4EhQ7sBZvHtpXR07weIs
dFQeiO/xfQVsbqQzrb0RGoknTQ42kmIjetNPKR/iIPX4jM9UmSo+VjnirMRiwWPo
xo5RMDRdstR5fsMtYn302PInyfFnWE65vdU6Qve2zLLyakhoZIrdjITb9fAjkSqi
4h77+TNY6+8wGqoOZVqB5AMYrNxaRv96AqNWxi6Y/fCZjzo+dsDgMwEvyvyMqbnq
fanT7gJCsoUgu0igdtrj4awumBE/iyXqEIMtw/jbMr2VzDvztiCoVHaGK8ID/AZI
zPo4JGoSeekmC5pLWo4ersSZHbUHRK8xi59ZUM5ddlRr9QTAlc9q/Ti1ciuYvvLd
6l9Im4/ocN0+m01D86fkHDuVm/tQEAR8uy78fDJTxVs2YMQQtlsb0GJ3Loe8eoEC
42YRo7SxBSw7wcV/ygYmmmxjc7V+n+UuezUZ5wAB6pZ3tTK7LonPchwR/6ocsSnG
NnOxECz3WuXa11hd954FqeHAMg98iRf6S9pZHgQyIEG7c9AeU35x1rTtQG5YpP86
DFVKl7P4ah+SzpC61w+8QrArm0Ph6pXdMkK6cVNVgCHWgOZbdQJLwIPpJ3cW5ez4
fJrry/QNSx3V36wlQ7W+d7hTjxlNG25oR3apmkasTL7CCz+ENWPNK2hfLCyzDMcB
LfDrh1tv6sbMWGBrlp9+ne5y82ZSld8zsU+S9He8VHS9xAL1AiOWyyKrjTkGExvx
taXdXyPbdEYXsJ5ujx7q+ooTB6U+REolBDU8H3Vwi63l4NM6WVcKDB2RRmlqGQap
U1ppEtSGbo4h0JwpFDz8daBWftfwFrjvOOT0cq0hwiNFMUYvtr+4Y4IyLqK6j6FW
40giuZCXFdSkCI3ACCyIivJFb7Htou3lPqOdJHIl558giaidh7hwmRdDMJ+s0Ffn
Z+S9imPLonicsVSryjQ69qoPXaKDNxfkKczJ1UxlVvlKW6g8R1tsBU8z/QpZ0bkw
B2pcXjF6KN3fmEO0jq+FtAOLDUWEY3XXS3dlgQ4bT7UFAiXvVhb5LyZrb5bizYox
PEMTExcdXITPfGDLaXYjUsfw/2kKxRwBB+cLo8Ul1NaUlDLnWyW/52y+I4OCEtBA
rSSMxKlmJFPW42WNlgEDcLnB3EHWP8AI9dUCbKxAdatL2vehLBQ1qHbh+1u2k7Xl
Ou7FEna3bKBeWWC74Qd6fBWmhmSCsjNUvSJZP4oMyUPh26ifHz4Kh0SvIZv6mKNA
2tWAX1qboYuhp06q6+rxhdi5RT6HUELG/XX1HeLLJGwkunsSJITEbaJLoF2FzNha
2Wsmy0e2Z2eOp5Hx9duwWeQLWnbRd0c6Ww7n924f7BfCWLeaHxkezisALLcUOMHj
ohREoj4oWvgOrQgLIYjIcRXHyLC6uqPPX/DD4bEjnlYGzNa60kPfTLTxgs0cpqH2
8gzuTnzi/t1ZsfBmcGdhIUu5vmMXY+S77Z26ltWNl9dkwGm+dffQiQlsrTjpR+ss
qKiEivK5iyZfTZKPyb5ywR5n+6ZYynPYkn+Ex/OFASp/96AmjXN2l3+cemlOPYw3
/EmEnuHLdcslacSbDUwJHjCug2+iKAVyO3pR+ejDwiPcTv0q3/yrnAmWvOPP53v1
iBzPwoXAKWl00lAntUgxOS+a4wkU99ueOOlOqDnQLAM2CqupEQbL4O4uiSGo3Slx
i/qtj7ite5I8p236OsJ9xiklhZxbNauJA6PfgMAWxEUIxhVNzm4ikHvkOksiRun+
hlKS8KVjPsymS38n9woJHEB95S5JxC2PUdaUvm/IM/J5FV0c+bIs0JF7GjL//9hp
eRBaXGdbDzneBlZTIRgF8rWTLAsKHjOEA1T6aoKFyuqJZIfxhbSLHqrnRJhwlCq8
pxaZmz1MjzJsjrBQpH3KNeqLHDfRc7BmO5XOOMe54GuiHenivpy9DHZ5fWiWWxBs
k7kSrtq6HS21DDwJOLorK6VsoRPRXXgn8E5RnAdxTJXyzO8W1FEFb/UrahD4/XE5
ZL4W58n6Yf8UkpXNuFwD+KPZqa6eLqb8Wo0uTjriURdcmO9LgkRtCzi10w7ItqIM
IuSnjtbtgMiBAwBNlJ/BpJcdJ7R1Ult/QC2Ti+gUixLeeyI3ohRSQtX9OnLsosfj
+Hc2kp025BzvWUcIwvhVNwvZtK96LaxO4JApPvCImzxd02GuSY+uf3ZljOMBF74N
/90UW5IDcv7o0J2onZ9qmTDvMweE7xxd4Enyihind96kg5RAAxOdQivbXDiwYwLV
Jr3h9Bx2gzJm83LaT7iFL2g7H79VrfBSQkMUiZ26hLyycj9W0OTl9MY3e3xVlpjP
DhDOyxtHFgdSk9KFX45L+T1w0GYqtNrTWqKsAFPrOgYFngpoxhGmbNyv1mnTwE6i
Ju55zdoLCSFGfzTLFCifO5SEGCa7TNYOUMIOy/o3iixvusQCLLWx6j2AhlfrO7Nh
IipzBTkV/WpUb49nnQ9K7Nu8JKQQKRBEQuk4nOMQKfVhZqPw2Ohylpyzn7xQ+Ioq
D5JufSnMI6w3pVsigavwCzHmU3U3IMXMCPDFliL1RPZ+nHHVNoCkOq6zP7wXjFp7
lu5D+TBW9CVrobwOdU3S46lix2Jikpr8ytqwKxFphuno53H7VWi1AnR8BrbxXl7/
kDVJb/zEl3zThAL+1EstAVwB9qNgwcSHQHh0YCLJYfFkHQOyczLNj9WLUGaYe50o
vuoYMBz8XZkrhxqrZUNoPTtLxFxnbaLAPjuwaaxfaylCf6TqMWRIEPxEquqIvXy8
RxfBLzipJwUg2tCIjc+JYL4zr5GWXy3GpzXqxdilLmGYgmYVdj6GUcdMTrnW0wr9
dtweIcYYjSWs8esGRese1jFFkstFvdug7wFrksbP2+EsOGTeVb7RbZjGRlISajBR
s0rIuZTnGC6hX/7PMyWUEpS/PZAxK1HpzwWPisHgXdb+pkuohJgU3UqsM3qvee0z
IPNlsOpG1QtD0GMZqePZBMwe1GknM9IUG2JPBOH+RVb43XHgMWVgZO2K/2Uxi+jK
kYt2im10IhxT23tZl3B1WD0P/jWDyntQs92+XwIabgih5ZtDkNqwL4MUpYVFDef2
7rMITHlkqW8aKiCLfbjwEnjudexdllHV2BVpQUbWc/NBnPxtdW6ESBYIbub7EE/B
Zq41Py6d8GTUY54iyC3TkJponGkTb+XOmrM6bYRK0yM8XYgKvXghrFWaCiLN9Ogb
Wp8pHGGb0iE5QCO1B8ryIRphZ+qy+u3OlQfCdx49gAYpUWDq6UYZXDvy2ZvX31s+
HLgHusolrJxn6pslzdeDPkrYzXjylT9/hqlGHBMMyZxVrBMjIzxHd823gxn4M/G9
AqFqFU+ou7ho7rbdJgiouR+N/OCWFcLjIpkDc3KLR8FaKG9TXkXj0VRT7ifc+vRU
RTUbHTj63W/BckYxGEgXW9v30hVd2y6o6voSqrAvnO2veKI+UYlpVa5GZa3Vp2+U
6axODKz5mWiPAnvtnAEJaX4hpTr3cLwplUXTyHQ89721Sf6S8tKpp+g8muEortXc
Nr8bLzUqhR8/2ma573RPHzgxF5FgIo1nQGI1ZUT0MHLzDWkrmk0e2pgkMR3xZMji
H/IS121ijFSe5denJmWUSAREBJFvlYBZV9K5zNYcvL6wdEq++7omTIPi7TFeBaV0
gUd2cfxNFeIQIgU/H/kMSmxbiN9/LplsWmM5qG8hv/ARcW3di8eo1XRkZUVjPO9G
XrhjU/cSeGzTY0IE2XJDS+fm6Bp14YvOR4LhiZ87GVZVWLqvqDq+1x2BaDIxz5Dj
XvSHK62tsWooZWm4UHOfkIrPXw/ZEqPm9SmNgkS4qu+7zX52d5qNGHpdRF7KEeU3
33tGX317k74M0kc+JdvRIit3e1h/Mf5Nz4xmLwo+H3Gh0WUcZcWgz04RIFW2cdpS
WTsVTKEV3UBLL85G31IH1Gs27xTMGInkSJJdg/HFB7mn+T5pyMP5bXdIWYJRVFwh
/3CPDgryHLMKPaOjznpGjN6HKGbepv9rIQ91a/86tGTNnWIkzS/98R22qy168jvc
9+Mt78yXsDEpElWJDyE40yFau18PQ8Zrc6W+LP0i6BFjmei07hmplLoC3NXryIGy
bwjqpWJrQPy8psJQWYuUxhvw3CUVvALhxyZRuhRpEcSNfJu07AyrY44DhqOQW2g4
3YQbERXVskhsHQlf/af9tvY3ZcaNgmC0NEVaFO+E/m9K8kwhB8yKb7eCsokz8H9F
NJ76XrcvMemYo6ww9jPYAi7dYZvbBZu7CN+0dBBRzWUG2XWI8ye4u9BsE80FiPzI
V6spWWVWcxWp/bIqhhAOfK3H9a+xlrVGVMnSihnM3ZA5xJMwnRB15qYIzlyrjazb
ixuT6xyib2YA1hT6fFJDGDwrIoUNk6yOyX7aG1/q/Dfz4LS7QrBuTQnkwNXak9UI
fONu2dLVGOHWFAx5LqeAm1JbIcbX3R90Tld+1UJj0FmT+LRU8VADkukMIv35hTyl
gyqr8At2iInWmJpQ+vu/5I1L5GtbfjT9SwVDAMyytZKLfpT5IxXnJEUSq6wNg7tn
tFr8h0lzW6EqY3XliL8ayzIEbbmYA7lyD+ndJF60wqtptzcUCPM1C0Y6Mb0Gv2yN
CR/FlTi5uH05gU+YdBmY1WmGJcczEeutYlsrLG0I36IskSQLWnA9xaXGk3g46RFS
jFhxY0431Qhv6mOnWWJm6Il+eYrAQLapRx8uiULNwu1i2/smTXxeOIqil00y06qT
TC/epeads4XNEzGXVNjmh8OQ1WFTGKG5sbwToFWuAQBwvYMLH9DgfdMZQUXD2MTO
QE+FxmJ7b7TopsGfC69n8oYp5X76Mh+Ud7oMz6as2ofZbrKoPl0ZM6XQMaMp3w+j
7QaOFwVhYIRpqkAw5whxUI5G7Qy0pEgBoAnWQtsQtP+u1Fx5ojH/EcbFyw956+y+
KEEsoZ0RNJLRIZKtFtlQ4kjADTRFPg+HhYFjSJr3PUN8qHgxqIszFxWxMHnkH3iK
WVNzdfHLHS/quUkguBvtJ55PFKxe669oMSVCXjRNc3GqBFUGnO2wm24seNU3I05X
Ir5wXCu8gsg4RZ/+zuHGFtrV7GPCJy/PcYV6OnHVCNbkkqe9eOpQaH9UGWaA7Fy4
Y7KScRZnH+f7AVvAQ8Ee+dEcWMh4Dm/uc8gRFzyycTeGVt8h/wmRM1LjHYLPDNcx
dnkQhp4BsZ16sWigOcUAM7HziWPyhdw56Vtsjrd5UzY6AnYR9cH31UlQ4Z+GTsLn
2BiOTzb9pqTVwt6Tjrl7fhPgkg8ZxXeDryzIgWqvkgV2HozWvhCnJONxNBCU5LnZ
koDjmwz0fvz8toxkTvOEwpFnea7WWhdJzfOH6YxQobYfi5cqXD0j52sY8LJ08iEt
TvxMtIEqVO1HZV0IRrEZcnAMto9+1Xtqqv1laMG42xbHn3Ea64cUaFiqNapyXQDW
AzK0/CG7BUdXIkNUxP19Gk6hQJRU0ak3IkJHaIuSEUs38/xemKffiQjYl8N+yhLw
Lvy6O1B8rdGSWIW0eKjvUXKnjt0W2LqCPB01i+HgZMLFg3JcPWX4j7a8lOwEBQxY
t7S3s0LF8EVuUUEcDEfvDgBpvkRSw9o9Vo6H++4jas9OQBPy+y4HFnWUmKpHQhcG
qawHfT6uNTg6DJsC5ImzBRx2OUh09u9ftvOiVCDYRtzoXDRDfscNTenLI2lAi6FI
N8432PFxNJ9+trhlTs3XPaQLN9f+Ll+9dU19uM/Eznm4Aw0n/nyonXe5GLisw9Jg
cvliKHSC4cVuWdBs223MHOACpciYMg9M13bgt4flvF0TiTN2NKfVTo34ssH0n+M3
r/TlyMi8cEuhIrCrjVHc+tveWKcpFQVx/aC3WEBji5OW0UQeMIj1maImNTsjQsFV
eyUTxFkxhNddHiFD4+pX0o52owCAoMwQiUR/okFHL+DdtV9EXyQch+UQJeQTlEkw
rDHLd42wZEzYZ9m3FtR/Z9wWs/dqRkzR8YQixkNfsKaeaSCum+yuy2a7ZMB4YSIV
5VybhVXwgs2BPeq1kkujfVAIuwZ6F+gxdhnR5aJj1uVUUcwn5LubYmaNzr1VMt8N
dtfrlOIrcAOSSDH6YxSm1v9yBm5sL+dygDhGN8WcUcKSvd7ZWoOZBW7nUT5Z4lVt
osTw5KnIIHl2kkVUfjKVdmH1pEgF3Crker2kdDgrE+qIVF3tuOKCYy6Kg3tP0V3X
QYl2ej5MKb0sDT4hY8k3/hy1IH7nf2+akxUcWMtUQ0e/3lzrQYVkC5dcla0Nh0V6
+RIYfIZKzqQENmcTwQbP9DKQuj1g8aelQpJzte24R6yA/kApwTDwhSmVc+/Rm3Fu
ag/ar1tkB5sYpNum76NDUIOeIbjQMkthr4q390B4le0YTNKzMBbCGGP2dAtg65+Y
eQqCdyX3mh/ypBL/UJ7qM2feEsrpAoHVztk72BshuIoq7OLvzaxy5TTCUg+DY2ND
dMaaQUnbtmfGywoISFNEs6XKiqkd+RU02KDVGpq+B8D8cqyViMAC6gH2XQUz/EQh
ajuUPvTEE9XXS/nVyRcKmd5WvVuFFw7SHtBw2JJehkTEW0yrKd3Ik/PpJLNbg8MH
iZKFALBGRtyzC/Q+7g8pyxNegmrm0zRaxIKP/ftJAw919OCLNKQ5yLF0zrIKxaU0
MhtbDLWc0QjNHHPH80ZBcz98k0NG677FreMbLyUONkVz1+FIXCTyBcKPfoYJ8fLy
5XMKKKRyd6KnhKJ5iDnpaik1irA6CThPAQ2nLw5DuMwI/9dEVp4wEObG6iiXqmU5
8S8dO3RFNYbbBU8Ll8R8t2nkcUKWOxrijzVNxXIh06KVw+/mtaIRPg7W3ehSUSRG
nvIsiX/vMw8dG3cT2F72HzOM0057pqS73mklWnJsuxhEZl/gnKXHqXaQZXz8Ciea
unhMpHlt6u/gfBDoxWVPGuBrUjw2lTaJ+213UXLqaSLCTu40vkLr7RIYs9YQ+umJ
JIuEIzARn9wogoBy/c4AnoiswtQ765R1FX5qU7NlA39AOVrtCmFANE9qt33tOCej
jk70I4Rk08pxtCuu3NRJNLR/QbcxNRX/UCqOda7R9JPZ6s9uDYUxiPk3dUkGODpj
ou2IcFpXw+6kosWnwzJg9l3KHMabmj7SNcB+Nq0SPKwDgjKLDKkY6sLKNO90TVTw
pEpXGqIPc1KhyIfnB48qlsBOzGg1+7xfGLqAujXM/1+xfa7ll9L9dKkgImcNlhpX
E6OOhnlPXop38lhFeCbtFNHnpiuHm+MUP2ZLrgBX9YASsZxFvpWHeHeji3H/I18v
NAqt+mreXarU6XcxJQiiZ+p+nohP/3liVwMlhq6H/Y2VO1a8p2RU67ZDW/g1zr5i
K8Bm2sXbnX5paQ2X9W7kHOFOKucOlWSrMxr8u2uEFx2qKPrKWQCgjCJFF+l9ltPe
oLR3MOlhpHWcyy0x4ooq/Dsu1PVSu088uj0MK5gmqLmQ+38BszpZkOGhiHF7Y3iX
mrwu9YubmZFdPGvcHurv9BSkBi9uBvDPsqVlCTBnW9ocyBsWua4JI155jW4NEz8D
CTSx1L0LE38hFL2UfFPicaLGfhh/OvtKWVC2rt5yhz8TSP8WNx5N63FAo6b8r8I8
FB73LfYNGp2Bli9gS8cwK0SXit/owaVQq3Fzo2KMhnNI9om7QpHDzWa75p2iOnhe
s2EuktfnXE14UPpgpdzXeEzt+0UQ7EKw3Uh/FYgkzCimBKfNa9rJRTLKxUkzcjXP
QVJ5FXKBuAP7A09FaUQoWGKw4WAdA1mYbld3SXImD+mGeTYP5vXgDIVWf3Tg+Igj
6AhuRymV90k1oK2zE2967MR/sWfnN3cEntoZ0noShfrI8r6rdJskaPcQqmlv3WYL
vwmdMbnADtzgGcRYf80Gb5FEFO+FmyksmHMJmbanchb33yGlZMJCWN2MIKvpVs4c
xV06tNmCo0VttdStyVWGdw9ElA1iUYP9JY/uEvPf9wtbQScGjM8FWum+Jbv5nozO
uwa8uSQ01ra5/Q03c/PKRjbO07eNup2EwUzrhSmmxiYDvWSFq3cWGUtLX03PuFYO
fizibEJus6c0SKvpSEJ685ROTEraYel9ffq0SvNqBh6cNehm3GSOZs6ugUowe1Dl
pwpG806e7iG9yIP/y6/X9paXL/0Xh5ebP0fhhLiLBT6bFQnvJ1L6XOUhQtcji18P
NQlV1gz5U/TDzKnR5+SqeWj55Xt3ImxbZOUaAWtkLFT7Gb2aXqGbY6F+gt8CFy69
1fBdlR8IsNHyBjUoMnmxjUX2wIlP0y1LW9OOKCgy8prejni8Jq2xdtccVmzqv9r7
6j9tjL0x22ht6Ddeh2P1YYKExkev25t1ff8ocai0MUVv0bUGv3dbrOJ4WWqBngAu
F+cAoXpe6OaMJFcDpvMth3y5sdHRZ9pEgUNjDIzturMzeFtybQWK3zEoRm5LpZNe
nSMPreM0HopNZQn85lF1tuHzkxT8AK0IrcbwG/InNEY6wPSR9LKnFgGH2cDZrrZw
3BcMpfoKCUJ/hButJ8UxvF/1MewoMowlr9BGR6Z9jead/Sng5TNWCnZHyeUkb6y8
LVErKxX+Tf7F31lDoiKdVBT727H/l6LFzCl0wgmgpz/JKMvqfxm/25sI8NEDk3dK
MdrCgzbakQAw62j3KS9+Eq+Q3HoCTfTct2GSIKoHw0R2EGG20SoJF3tB950iQRMz
Y5lUvPuXYAm6EZduqh6eKT9rnxkpw13xP5Q08Jiy/mHCsM1vQKAa3nYSP9fN6tJP
+vT/Bl6/n3SJkS/z6t3jdHkQrElgXpTt8kAW/vZJT4fn816V1x5BP56C77yhaKlJ
xo9XSMgmY1MUyx+N2req4X4ecZlnzG7ALpT/GTliiFhTkSU9maITM1kQVOlfRb6N
8Zdu6T+368QDPDYkSMStuYYtGQnKUJUy6sjDIAJ5Ivr5ByNc9lkKMMLSTkU2CnSH
Xvb+82EXiyOv+f+Ieqa2QpF/Xc7QoB+9XG3EjD2e1/ABd5WR8hRGJ/NvT5hr30em
WhTX1Yv9OFc9Sk4pobuW6iyl97xjqpNZGYm7WzBJK3tpy28xsJvGg146FZv+73jA
aHhXZjF4Lj9tN1OVAz64l29M76a0Mh1uDyaTzyjJaUw9pVUKLXx+qr+vHpvdgu1m
9ZfGNfYiNdgfVWIvm+rPcLr7Af2U+1bAO+B9gwVIusWftOv9FchKZxd2S8obkDn6
+dj7WxzWYaiY5ijJHJDBK6d6j0A4CF/zB6ViW7aBvh2Px46bNQdM023naHDXOYkT
9SWKbqOhag5tBvt+iyLuZmHeEFjqkTGCwDlpWU1ueQBeX2EOKN4bCOno/Lzxrxso
qNabVMe9yvHAnWSP/7ePjk6c6QNO3HoaBmOQ5EeLmn8ZYdNZILZL+7e91CPm60qT
yynV/CleFkT0uq3lEgvxtrKO5QbBvj5AI8fVseJbVbQg/hu3+FRzrmV9PXF9RFNG
o9AaIE3vVdz8uaQZjrrjBT3QYuTcrdvQmTFAc1yVw6Mmv/ikhbnVgKuAJDHtmEgO
7eopclaYkbJBJbCz/Yw2CY4bFkUWk9/boOeUlsPucD5sHJko9uFyK7MD210nq1WT
pcPKk2ILwmlnTjiNa5NFsL+W3KgFcsvL2sZj7NvMOcWvGuFN58pCLwa4QZQedRYr
xUlYSNCz62ZtPs20Go4kwtWav7mQhWCO2Fs7ZybTt4tg2hUkm65FkGGg8Kx0VZ1j
tfz9zAdB2e9t3VMLZvnGJvBOoUEk6Mso0n/oATqlvNZXSxr6NrgHaF1synqdJERI
Q7U7Dk+Umxhrwa1TdIjcHCBVgbp09guBFDolo1+g4ckQXcUdqHgRd23TlFk8HPF6
38EOy+lbrIoKEEkjZYeeeXhF/RpXwQh0vy8hO9v3RHKTn4hzYUcFw8UzFwDh4yld
5ajUkEL5YblEcxYlP8r1uJnLc6n7e6BejwvVJ0gjqfM6/8de5biMk1E2o8eD5/iz
UnyRbE8HHruTaBkMUrvimI2ndHDoL+MeUOCpIMGa2HmrmA8084CqgXSB57ywOJf3
kFrZVNrvMgiJeAd0K1kK+u9ako0mZMpFcGHK/vQrRmv6CxtismXGDYzhj6LiIs6U
StqtXPBAFLXCCApg2ZNcvmOoaXC3A4IR72G/Smg+71mOa2UV4fwtPpD3mwMN5mXi
3VHs6xIDU28sp/g7Jn8d523PjzEpUDbbZWRNoR4iy+wNG/ZQM6oMVC7wNkZ3RnP3
DajRFH0tOOEhL8ibVONNe7GH8CmkFPBDwD6OeNP6uKfekY+ho5xSa6KOTKgl46WC
rByPFmEWkQNFgcy2w0jy3JF1Dc0DYMuLW79BAz+i95lqLF6ksT9LVvadg5SAlox6
L2lMG5wjl0k6iPBtWAcDBWoNfgzDDQI7Qx5lZJKDdEzv7Pa+Y6Xh+dZ5QyvgegaF
fl1yBXSy/mF2RU0wL5BDQt+qPy4o5OigCJoX2d6b8tWB2BdMBYWX2WvaiMb+xmJg
vRJpoYbJb+62N4xoF85fLTqlnGeqABzGUCKU0LEYef1x3X8x512ltjQ8h/Ai6TsT
2bCuBPTXD1TDikHsJeRXhmnj3d4CjGGSLRjZBdhqeIzoZqzOPUCRGpbZ3yM0TOWR
9fyyippZjDwXu5wnVORNfJAmBT+78nXefFKPst9q2D5EVZ0FSvbdvi8Pv672Rujy
/h/nb4ji7arH959mhp+dmMmHZMvL3yuqY3GQZle3674kLpziphk2RWDYqrE3nw9b
UYxDFxUQk7ksEqrKgPlYOA4G0uxgxrXLhCV8jGw4SxnVEJdXlITL8kD3waE+/X27
+oDUe0QdiNl5dTe/l263vuJFxw7BakjyddZ4mNOVHfmvC3+7Re3HELkjGaIZpdpD
rrJqL9G5Htgw3dUy81Giby11bp/tF7O7k3RR5bn8/71veUYGG43AiRAdDunGTm+j
+4t6pmR1yy2uHyngUTNovGKowCp4yo+rSvMpDqJxpAG248B1FoRoz+f9XTgYvjDH
aCRO6i0l2OVfbBkl68IWyfiF8bE/zibjlBI2q3zkClaiqyEJiMIm5P/q2omVxMAl
oY4hcOmkWtPqPn83hOlQgPl5gabSC2NFDujHN4998yglleMy3CqvMepl4G1Kp1T8
vjmkAUo2pfIMS/V5VA1kRvBSWUTtwOsQlVrExAY5o0XjPn+PwKf8DAbS8hZuNB1d
j0yPTA8PGdnohnEgyDP7oBavucjIO5xkKWmW13WisgZ2XoonjRXAv+yhGwzoh4bu
1VR2OmtJbtTAZvA3ZF/sjS9yrWZC+dQOI61uTmOQ+IO5pI8L1QIvmW4/AAuEwUO/
kAKsFYNlw5S+g2zjJkrZvxEHpiiFw+WSxIfNnpxurqmuD5ZteXEyIdnR2VBqQONa
tTxw6/Dd1LHoHZ0SetI04CuV6HJygWj3+ludty18w1gbYrkSJej1UBoIDmbKPjOo
HX/qFQxjK2SYmCUrN68MMq/hzOXfA0WU+7R5ZLTtVQAP4g8KJTX0gWKC/ekYZ7k+
qEO88OGGfeGbmJsWoWjTmgvsa33LPhPKnn63bGYBJfXenO8M+Z+Ok5lUuzpZWnHu
D35/T89QMgnCeuwEDYwA7y/wWSHRGYODd58zAf2/gkWVEx/P6irWJpVeTWusYpQp
uExjGtwevEmerTz+kpF2iktk2JbqwYH81Lx4SLDa9/uMoXqFq1x9vVO64DwavX9O
pXQGj+yBRh2xGeVdPI8CHnEz9zHYybgob52DRLXVCmhctMX0rkpTpfWjlTfYUgqJ
fa1ejp3z5UshW28Dc/ZQy6yKrdD1gW8GE6rsbW1yF+U2+C2VwmDeLdiy8QiEvPFh
3wocp+mVkk9O/ogZX2ePddJ0qq7h2+fjmYlwOOJm+hCgzFIYbP5u2aYP8/4HR0ni
KZ74avbiAWFhbecdcPz761L+mgtsYeKQp3Numq9P+DGm/CZA/WqrvNliWmTCypsp
al82Zo2uIBLsZbunrXCu/23Q8TJ6m9epmswGKLab8Pbdk36+u9vbBiRY2LkNXa0Y
OZYcz7RgBxZgYFdZHk04zMj0ovcqPu4jOa9mD1/tPcL1ClFtkA6PrYtDaKTrSWq4
Wh5kTwlZSLhLA8PrpsVbauNkRqvfsz/jTKb3OhDQgEs1ldoqWAiuyeSDMVp3R4wj
H9tiMUTNP8RmAR7DGtQIM+aKENrQCbTksxp87+Z27xYFV+A6/g2yZ7zQ+s41XCY8
nG8xlNLj8JwVIaTBZVGelEdBXsIErvjZVa5BcwX7cIXCMHSSVeBpACXJnlfuwSGC
TM4q2+KLpg3BXEbN/giy0jLVlbAUWofrB4F2vLto09kn0DKzVuhlTGUBnUfV3AQk
Tl2YlIV4NVf05F4qwHeRVWpAaUMgIzEzafgIIlikRRIzN8OSxr5W6OiplG4Rnopp
5ae+J6zpmek5FSVxHaDbK1YDiwqM//RU8OoZHYkkoosvSpQOlmAZW6mfFnH1nRq2
S5AZFNoRoFCovTuzdiULjGaGcTfQoJdxaF7ZXQc+Fm8mydEsepe3gX0fWeC8uqEn
uveN9GEtN/4KXdUL0ZTzo8hqM/j7z70K4vUAp7HnNTm3CR7tPqlW5E8pTr/auyKb
Yk6t67us6RbaKfentos6J/gg5o1jXw+bDHHaG/r8L87okeVcYlQQvP8israrQsto
xcwo/PuGFpwGV4yVIpiP4avbMPqXF9bF3rqdCA3ZZagHU8ohBWI6vySxeN3HCMw/
YRUgqBXFeYl5WSa4pKQS5PD6z+SpAgHfJ44OYmaar0kRK9iMOIyuCPqLx9LHibS7
UmeoRtgB5vzRj7DrQgnVonRBbg1L7gAKghBBskmJ/36KkaQAx6Ic5sMn09mwfyLf
kEzRaVHZN2Muj1eD1aPyeEvhbW774plSWGhpr1ShcLf+twEbKVGWSEjNbwz9eMs+
7Zt/UXnhdiEe7n6zySIJ9jg6GqzPWhcvHVHY4cT/54XuBKf31fD58K+cDJ1Bt2N0
rmWXMoIlweNWjOL8+fKwz9/GtiObR8lfW6qMijh/7lI/M/V34/NejG9b4YRzXfQu
IpINRDVTpmz8nk3wVgHroDcesRsX2SaMzZN079hWqh2+3qgkg6/q93OL1Zd0z77y
Z69322V1PjKpPpMoF6zw2cTwFcLoXlwxV29hSqu+rwmsfxNQr56vn6lydzXF046e
WWcBjpJZ4GihR43ceI1FVeulrTxA/QtDZfs4R/ov2sfCmVx/C4raOwb1VIMCpJDq
a3OHyTMQfknm2ddpkVeJhp7RpzU36OhHe6qZJOXsQfNEC34nw0HHftYuOtPO0gJc
AGt8dI8EpyF1FwGWancpfTHWeUtboBCSUB+wTOojuGcg1C4NkvedKRJ1lTTVIN2N
Y400TZAfWREmGgctDzmkijgPDxO4zLjZtdVbcp0M5kFnTQLPOMRb8tWmr4XQQNZK
sXZWh6AT/2v7TTpGb9PM6LOe2AZQLmzqj1PGRBAfgtq/5aHsKTYcZunc9rUK2XU/
HuCJcjQHD7z77U8d7HlqF1ZJji/ol8W+HjHvuu7q6Dl5Aelen7XDPriVHYelv1Uk
kTkRGW6sfA+METixoRXJRrl7L/AOmYZ14Vg2Y659NPrYlean3/kDnuLOKBz3Xln0
pp/cXXSaSlgRNTDMtuy8vEmIPGxjBleuzboucLbdDSa1ZfgGkz6cCkh3c/0t4B/h
TUv+TvtqEYz/p4qWG0LTi3Xq1Uw5sjSTfIB23JFse8JOMnMicH3b+OLOeM06SJ17
PVSIrGzfdKsu9df0HmZ0Dg9HoSo6YqhzP4dyQoIC/jOvS53qsLh/rfts4EOJunWu
0nOMdf3Rp1r3Q40rbZVZ7Mcc715NifoMA4pgZYVP/2yEuC/6Vd7P/X6jkKGwGZkb
3WMv6kRfXc5YrWsMJLgN0p9DOgRx5kjYg+eYBFMJS43N4Xl/TBl65KpJbcsfQQJs
Q0swO7FwMALNNcSIg4n6NrcInj0RqzQMO7igfA1/++PxU/ya9Mq8iYdkcRlYIRse
DReZ2iurvCOgC4w0ZrZnNLfKmLUD31Drr0iQyzOZAPP0Zwy49omGS9WKhkjI5dWt
8dMMq7LxdgWARAwQ81DaxP/nT4K5XonVIcdgoUnVfBbKnuSNTOz60NE4pstAK0mc
7fsN4s+Aa9YguIJNgOPIPFWe2RL8P1/S7F+65vDL7as05tt4XAlSchYgnVi6MQbs
pEPUo1SqVF/Ou3iZAtqDy/NBN9Web/dzj0/YIjyX+gWN9O/OKfzjkavqBzwveiU+
pjdueovfndmbZLsCFeM+MQTXXvi0zGX5GAfcoAGjtxmXDWMfhyjog2nydcAI55DB
03NfZAODYbwrwazGI3yQ8sSf+S//SFu8TGuaok/gHBJlpC2rCPCRf5U5mrmvvEYj
AippOLMJ0t/kgKhIGhko90iPUroPMiK8NUmgl3ra3x6UyskNoqJ9Raxl1JtGvnQN
f8FEr8c+9KnJb3Co2fRPfZ1DhfhtpuI8Z7dnK2n7IkCN1DYl4K1zccohjXmdb67d
kKHT88354/7pCqG6m2NdcEuV4Bv+ogD5gkUEoz0I6aOy8tqMl8yZIJZufH0ttj9S
ZNbASvEpcWKDagehbZnn++fdTeGDNi7mGd2qaI2OiHs0cSElvdWArdQsOcrs95Tu
poLDlVAT4/KxOwpyZaHGHhrGgmZqLqbISnc31CpKLVwlCaRc0RS6Xtgzc8s6zV7Q
WLqpXtJZ6rcYIXWlwpwcyLZq8OhFivUYNeJ2y/LPy94zCyQBbXnBZ6MkCo2nIn7B
ekbngcOB1CicPDr+fX73226YLVX4iOLP4U6Qt+/905xUIz94hM+pxLRuNofhlAc2
tCzc4bRjSf+BABwv7X9yiTQ7QUvGtxkzghRrVb7UsZHxpkV/4uPYKacweHvoudNS
uXcZ7KN++kHr7qPDRpVgbTRWjeR+znuQP+/TOgA0nm+2crbgBfnA0qAXEsJZT/N7
wX0/1idOgAi3jFzTFIGQqbilkcKsSp7+hpD5UzHn0JIDm+1SITY2jnzOwwqNEUEX
z2xX6gRtw4m9n9fa3Mw7tkx2uHHiopItbhrs/A7eJ9Ygmh/uD+gik67kGGXkq9U0
uBsre2kt1GY5unIyqLbxU7J5MFC99ayewrBKCGIfOXsAXMKmY/19s/nI/ES+nakn
SEAoU2AeGvsUNAtFgBQ/wyeMgFx8skTM3zcteU21xF/5unY/okQ5M5UsVmm1/4pC
JyfUs10wzKNRyU+Cc+TaGs96Z67zJ/4Nf6NVbuGA9kSfMkiKvAvyLnIpZnMeA23X
a2+aeUY625Ks5nANrV68xWu07d8XYb5JgFoi+bqOdaGz+RbRJT/d4U2H8pdi8sYs
Z2phH2IKqxRGAvknXI7WkP1NHsEArfx2uGAumz43s3vYcHxMbp+JMT7IUme/JS66
c0pUkGAWRZLt+M7P1nl5a12qL6vEVi9l0a2Dcx5pvK+xGTIX3FHsJ5S4V5nbDKhN
nEcLBKht5SfoCGapJCOkZrPlUbd4SiAEnpA9mAMB98kL+w4nuhxPPwmkLsjSls9N
it7ETAMIGuMVxChedT5p7hxul+G9sI14+M61po3a2TlWR/Wheu3OT1MEjKri75hh
8UbPN5eFDJyIL/uODY7gt0olsbawvCblPmZwtXvXJ/kq6SdBnXqsu1fQXGx1uQZd
3TGufgExYXFlVUNlDmLvupWlSgMgWQc6oEknhFhsruZxIkqVFjtVj67dUDFhJrBJ
IBiwgk8Qcz2YsiiyOMhp7ImCz7vRw/qKHypPo7NwBQyvmoORF9yj2XC8Cz0o0JkY
U+m01n5ZQBsR0gTtIkwSw7e5Nf8cWkU2b2+Z5c5Lk3YLVcUdj3K3MK4cIwtgtwAO
7MExpQq8gmInrn6QwSmMzf0HAurB+xiB9lLL/MWkmtzWF4bUqRN0PKsKSrXB560j
8EmzFzySYNRb6ZP067KjVwPr9/+yz0c/IwI+OH40xaIle898fYaAhODC3dvwZMd6
bZgrSlYQ8ojqVwZGmTX0NJdwDRht7vOz6JH25KHJ/MnGbs37F3uO+fYZwElUZsRU
xcoREALzGcFVdUP/YdyR4xvuncn9T3ZxINfm7402oRkuSayhrEEX1CVqeQUdN3VR
Q5HSQJJ8PCsRNepsMrbkJqiJnKXVTJWp0tB6vKp0jhbNIFbPBbuvgidXZ6rmEJmn
I6ovikBGtRvbBPnaN23bwocWDMDnbnSbzThZTiVCQFeTewokkfqe5OQ7j86QSCBl
ScVo1Sw4sWyJfY589ubs1UbofjZx9wN87mdJVCmhI7L8hkx3nppAzkz+snZ84/XW
DTG5v7QOKso1Dx7HuzF8pQC2c7F4YMQti7t9jPKwYEysa2Tj40CRj8iy43b8aN/l
n+2f6t20USLwdzLD2lFSHQ+LbPVoREyv8B3HpNqGHyIQOjhI7aYPSAP3SUKY/bX5
GlRn9Ro+2q7zu+NrI4CNhAgKQZJ04nQqxUcDjYzoUJjFKVwVub/xSa8Ka0gB9czk
KItilfSimEmil4RSfu0ruiZhiK1YcIbSQ6z0pKPcQ48gEEvoIFjZ0kF9Qily56LU
bA1CuyRg6vro3naWyBwzyIJXr/1fSXImkp01yDWT5KV/XqYKAhzMQUNccQyt8rxm
E/dNkxuFNcU8vu15rg53EzzM8u520E40jOhadTyb2mXAj4e9rzjmj4ckX2watNx0
4y8uTT56gM8LEIxlNDVNstTXapqFY49rYSlXr6SbE0lfl1RDMSXYQ43BkPE3xGCW
7Jwmm/Vg2cELaaMvYH2iA12cDxu/V+vF4xmx4153jGPZfv+R9PdZrAnuRY+uj7PV
Wx8fTqKfPdK24nSDuzNfGLkicss33Mvhgghim3LFQBu/tgc9SpInBN+to1noIy3r
+mn7dCEBOCQltKKVN01jKiwUM0xqVkbkyjrf/e4t+ndCZ2e8jxWs18sP5t1ySIDJ
r0/hEVp84rOOmHo09nmZpXXoSD+PyFz9VYBl/p9BOl90tFcFNksDUORDBpPZOZ+X
Ish3vnDi9JebbLlCww6a0Onxdf8ugRcPY+GyMXme3NXNppnKmO19Ylykait8G5y5
W/mPzJ/6SIu7jhX1Mp8+gEwnQMu1Bx0xDtfFr4G975jh5Pj2gMBYEAYv6melt6Qg
6eYkeNypo0ooXaRhrHseufIGKzsMGoYfnt9D0mmNDaimfZ6jWJFhgGfzbpnmaCsd
2JvKkaF+6dXtvJp4d+UcTN6FqSkKI1m3pZEz75ZtCTUc/5cbiX9UceHRSvsxp0Al
YKIR3f0rWu/qEZhR8p8wDwfTg5lWbZhraGHM/9B7IoYnhrIGmg51WsmrhJ3gXHbR
fx65rEyg7c3cnWiqktMNGQ3bby/dzTCzmkvoul/aGGDgTf1MTlB5BHhPZGyinOFH
z3eKC5h8MKNwIO+Pg0awE8blKq+1IJBnxMKwa7hnIkn91I9rhOe7pdA1qGCyzjjU
X4THCa3UMSouCLcBQAJXs3Td8Kz5MtkUdWkZuAIX6VdIzkOsT0hQszWS+8AbZo9t
pjWCD4xKOSevEp8TeeXHUwAP6sv/3y29rx9DhemARuERp6m8rEkwITC4bdmCOKjt
ydxH4ODY3gNgKjIdtVoLW73HUd1LrR+wwZdgDPtK+C6Ar0skszrgoyYyAyCx5cpf
bEbjVuJuKB26Rn2fW6NTxkrGQZRhXK11Gj8F+sOBKoEQpjVA44ntmd8vQtBkQV7D
+O6JdD4cNUSiUnPKV7inQOmP1F6PKLggQN1OHmHTFuqS0zXqeBGjDSakJsUoz+TN
Cd7aXv+bmY4u90RRUeiMepNwnHvjUX4wl8k5TKYPnDLF8eAwKDEw46hYO/Z+mjcr
PoAC2wfi+1SNckw3+IS+T5Zczh3u0JGwItxXNGM9Eo0CU2ftnoomlsirWtGnLyR1
sFvfh0ccpj/WUN48OBL6totx8u25RtJPlM7K3SXRAwluBBAcCbzoiI0qstn/L+48
OXH/xNNSYyznpcdMUI/YQM8/SnrOPlMaqaJWzLpRC0T4z15IWVH40sjugoCwG+DZ
sVdzaELzowm8R7nkFFceX6/2i2cHIbQEUAP3Hv3OewiojAj4IzC+pLMgVvxe2nKW
aG61bZwstKTOas1CHhXGaAplIb/KYx6IuICv35kZIpdwuQUVPUbNnl/2n7DLOcR7
dDt5u/zJ5U0lY0D98Na+Ik5Ruk0pCdhdF8fb79rxTgSUaj0hy4iUzKrImgjxcRuj
rFR57M7+YNKQiGf4LabI+nIJdJfIsFFMw5TZk3QO40MkmgLynQweXXVmiQ6Bnlrr
SBey87u3ZmsD92FAvip20yR+Y/7+07hXpzdKsUsZLnkyy/z5eo+hpRFxhVF9Nu32
g5HBXes9aNCOwfTqNfky1X0nx5t/cU1IO8rbRdHb2sAAvEip7Rw4EHufQOaicuWd
pa/+g11xSbIOlCbBNb908ho6vrhVVtVRgARDDhQjvya/ol+QFfaEnMitp5lDxkFR
uJ6Y5720iXyns6f28hS5CbA5oEAViNikK/p75pIiblbeZI4BDy83kpTMZKh2IRxH
9QrbRKIOJgANnH0iBeT97xEiI4mmweLxtkk33tB9IfTntRNsvfwiYf6BlvJOJD+b
VQRweAnc1YF042tsWP+hrTlRFtVGjsaLe/4a74MP7qu6u+E4QwwtdlQ1NO9oSFyt
py/Ck8PjV3cP/zoCv+V6U5ycVSlVX0uuTh0htRc/sVSqFHdsBep9N/ZaMbCNQKKm
Ak+coQYe5iN6bzmbydYopqlgRQi0tcZuaK8OFHJWWUNEG/vVVm01G31xoxEg9guw
63F+CRjenDgQj8h8jQJBpyq7Qt0EsDYEpAymtq4YQ+iXIBMrBFy3FBzoy3pjdQ2p
Zu/oUnl1ZSWdN7h2f/YQEf30k57IuIbfAqEPT/zl1i5k1FVC4QNboeiw3HPMfXT6
EIilfbvuvb4mXnse8VtdZ63AKsbaWFJaHSm6Hz3eWpcdxKsSh/PNsZLnXq94fxOt
CQcCDWNN1c5YByE8VSfrOP9ScQmJN/orX+htPI6ckhVnxJ5jiarmcRxFP00MhCUJ
Imo35Tug9LZmm43TUbvbB7Ae6ZmDRukmL6LZQTAapcnv8ucAKAbZCvqQ0UtupIN6
gn3CBtFf8ORyoK9jbLu04eBW49ve9DJBQJ7YX8HSMv+YLvqDL/YpdQXuQ3O4Y7WL
eOlS/Ip0LlAUYq2cP+18B5wzLCOWuCibrkPR88Mw62GhbYn8TfuWI6+2str6agXK
147YiZl4RJ5XwQwRhEjhhtm87IW6TR604fZPzGvCRiiNlhVfWSbzyNr6lHYtj8Qv
J1Iv/cEjzedBF1RmaEFalODO4GOsKZvxb4KlslHCxtXEZVwNlUorf6eBQxTRNAZP
8BnuNzKfJmaImkNEjl+YR9CCmryfK/oJUQY9JKyU9le+G6o/civQuBG2SHQIKSlb
ATdeK4ol/ZOhvb/po2uwPDdS3/Kb+230zCLrlVfIuNLJdYkCPIJKiWLV+mnf9pDN
t0MNKrMdUY12474mTY4oFIlk73DNuEg+4zZmC8ie49mHSfGhlEWxJZ1qmRyikQcl
JS+YTIPCSmGLvlgm21lZYUY11UnXQmvqfO79Gs7fFrhdN8Tl289ayIabHHMEjWDc
MKKFeBBNClykpHA9P9LBu8c6H4vYvynkK30AJJJKnfEFzm0Ok/r51IfFeTMeknGe
sIx/nZwlXTqvHARnjw621PXbGiypd7s+kvgdT9xP5+CN7zytcKLPPBoZt9s32XSx
AQXB2Moh1f6IUFnbImbeV88fXSRISgS+9VElUfb5QodhMt8h2Gncd2r4B8FGYoeC
EsT2ULkIf99on/4TXPNF2Ankwa54Qnnk19ge4sh37JSUMQq3tlRAR/v7fkJfLcmQ
4FSW4oP/Q8B1n63O9d44y5k+yDxa2VIF4yOWN2hWRc8Ae23HwPd6Xe8Qq81UyiOP
kxeGn7URZkURhSSQJqmKrHPqoTjhSqC/a/Nsq8EXpC7cLGDMms9Cib8NbVHz7I4p
v8ZY6BwJOaR78KjyunGqwKVdYPi3T0Nj/O449BV4WjVuTRydZkfg02H00cSlCX3B
lUOHi/pvi0KVZXDmtiHSM/aM5AFOQ0Q8ZmJE0/6SNYGKs01zhb81wUaZNyfe6vZ9
uNfvpLEDR/ucf3fGQQ3S8v+P2CFeNpdu4vSpo0P/UlLyFZWShEfvkJh83VmXFXPm
ZsPWaTidcFaYA7NJ0gcs7aKIT8pMyYrkjywOVpZkGzLMi8HmLkBrDYyxLG2VY0zT
lPJxbc59jfPDXGdMg6Tc+zjbvrR17vQsKNhjXNxzE4WpTfw2tUqcP0xHN2sIO8bh
Zh4pbUP6E+CpDxxCB4yDH3sMoc01zby7l5RYZ8IV9vL+K/qdN1hJOraRMPXss+5x
N35pf0GzY+yS/+CQ7rdW7qSIgp/ry3m2Mq+wZ2mYHXwC4ByO1e5GIOfDuYr//ThR
JL+MeF6VUiWcSvONKwxXkrDEY8JxoDXE4HWRpMxKEDxLZ3Hlfr8WaAA+/LP4CIUl
6OmrM1KEnwT24o/iq7eN+BsrODjOB1ay/L2Hq3qgNQQ9dudLE5N5iONKabvH2jlH
a1A6npc7LD/8nW7DivBJjWC6GqubgPdpcjPxvdwa4i5LQa3m/NB3EziYZ8wiadP8
6127FBJM7GlNW+EtQSjLGORfUAXOzTdg932nwVpMgyf8NMbGYg0RMCfPRZHAMOLc
fIb+9JM9hka89+8uc+11knoa6p4fDR21M66Oew3mR12Lri6T3awJ8K82eQuGAWyU
C7E5CeULRNKUhkNYaZ1H3QEvsmg3YofdrA3wjcq1yw6royqJGnaDgCCD4K5nY/C9
+qxi1Fh8BtD4d5i9Bls+zxsCj6YF8X1qSHbYJDhjFQZ+wcTA/TV9g+ffbLKXa9Nr
rIElbCWPbIfVw4P3JDaOmOYf8W2ZDq2Xwgkd37o36CPaJdi/Tup6FCgtrg2J9cpT
e6HU6Bl0BSMMkWpP131tk/Of1MC1M0lZVTteJrKKRjSNgr95cAEMPSmJqwUpzgoZ
0+5wBKB1yPEVgSJjaKNwHp2ZxLFvwmaAxIHmuGwJnP8Aq5ceVksseM2HPMbEhNIg
snhdRfCyr70vY4wJvGYMQFt2/wnvS8ePJwc6JVmTnUrRfZwoSUb9BLuzFSYrTWRW
us/5aTwPDKF5Ni/lnAzqs2QT3rQUGpERkSiH0diVOAFsrs0kPNZmuLmenhHVmBYc
5fLgHWEmmNGz/K2cZV1rngs9WGX2cbzn7EFCT6wIyRbvO781PTk7Ug4Bt+lpqKeg
eXxTJ17dnMbG4IjoFw0hqW6Z4FOsvBDu0oIvBKq+B7sdsAyYzUcTuXWMzBuns1TJ
TnRUOFux0lRuja1PdeJQ5IuZoVAPGEXvLHG8VuooA5Q/nV2WlXTwyCBWgb2WPTr4
AQ0iMmWbowoAkfHb27wYtXwm3Jwh7wlXDOvU5WoPpiQ6EXV+YqDFLjJFRA32ODTv
RN8J4DXC3Eglo8EaG7M0mnyxSqzUAayTc8hhGZ2ChzIiN84f6oTeKKFON+DEh0NM
onZ2SD0mSbf4cJZ72GSARMeIYxlJgIKqATWchG5D4A83pVXjXUTvTrUB/nlkgUwM
K01EGJDyDncFxLC/AGs+yrIDR29AL01/qBP+PbiXVoziiJ/cPCQF91Ov6NSW99eQ
4QHF7HC9k/qCfeyDMBT8NkYQshjLFxNWEP40fv7gVeE5M67j3S0b/TMPPLFi8X1N
1z7qhDZXaRcP+YP2fDFalXSdWPGp9BZ1aP4OhHD9fM2xe3nij+knGCIzlVeh5XHn
6Sbd4AFMlXXNrV7rkzXX7Q4ZUCw+0hTi8LL/ky834yG2oOAmjzWhrAedOc0ZBWPA
KTLrulope/3/zn3yV58IVo5FVC1UHHwHPr6nRwAX3ZFRCbDwPIHmwXR3Y05zI2jY
RCtcU2n7p7ruAHn1w7VUWhVvZJQiy5ZbehodgJZSEqg77YdWJSpKpc1DPMDxJoBK
GAOixB38qdIDSV/f/uvXj4MWkAKSkTNXMa0JuW/DjVZJXSmLIeIOG83FR1ErGLgX
ZQ+Azt6cxdA+SKnnder3zh1uYiThGq8dItbkrhMZxgun+/MQzH7apSuA9PF7Ujij
P44ouIgX7hPW1KAeHGGfZvuzuiI3eAUFoNTJ/zZFMIlzuibdzBxVaEFN3jB/gedI
uwvvCAHDHAYdXh3iNX/3MgfZg8nKSjmfxQq8oyBrvWoPwqkgz8h5cE+1CXX4y8Uo
zpgi+CNx+0nKEisrFQCPK+qcDPYWlkAlm7oJkFunRENuKqsWc6d7VHDbUjqVfb1m
2F0ymmeQO98QFUrDcnDzk3PXSGT+NoWVYuG0LL0ldVEJyO+RA3o5fSrhOSKJETgy
GJkMwx1dLdmmz19ijeqt3I7+e26T4v5fuNXPZYxA0N9hqBU0NjSjkTUo9CoMINqV
LeYrqX52QfpLzB2rRB+uiwgEwp/iVgbazeEWCS7djQPG9cNXNbO1zzMU/Z0zWGE5
GjJKGOOxOG5gSAdFmZo0e5G01LRr5zIuPpUjQZVPLBNfOsbDJRuuDFsMNDdHaQA8
tK1yNL9phiBz6nXimPTBMPmlhGNbM3RCwhTPoQbLdDkik7lLqxJWsQK2jOG6jals
PfcGz1az85WkiRzXYBdXayJhBbQMFmVuM89FDgcHezTu6+eos3Nt46GIf7G3Ole8
/ddvC1d6hq4D4RYtkfQjQwQgwLa9vwujnAWDlu4N3c3EzqrPmxJHhNdFL3np3/kY
gD2G2fcwey2n9b0yrYrtv9QRxI+vqlVgUKaFK8rMmDrrHlRf4SmfbL2LFEn8miFD
QnH/Ux9YRlzri1k6G9xWgDF5pn6hdBiyCURmin106zuSVmavkuA9/eDADrHqd4eT
TmByra9DjoySRtgHHVpx7t7Ccj6mmWoZIPhwwqPFbvU6608da9hmHBoovxpB6JGq
RXjkjV8znaJDamU4wtgb0yneO0hnL9zQPc9KFjqxwqfEA+ShD8YIXKahSkcTbZXW
trv7ICqHc0OAZTY8oeElwtnITyGWrwWmdyicr/wGw1Pra23C+PQjdu5kKLcSY+nx
DZPWVNhON2b27jKA8ZD8YarFZeKdOWNcGON1y5hV/mLKM6Ci8gRXlCwlzxlkmY1h
XMB2NhZbDYNBA6aaAaPPVKgrOGnPIVh1LfzO5W3iWdkIljQzg2qBNJXIiSkR0UMx
1VgMReLQvBYyP53Q98VmxfwvIkCvFlMPvMRCEH13VG2Q1/J/YgieLWO7WzMBa3yW
muA887H43mF5BiIsTFe2sM0Ry1xaI8RRRlA7LRwu6LSbiJXzQmLt/R0+5TJ4wGcT
vV42R0xZG93yiR1oXvZpif6VHgrNZaAg4WytGgzCF9RfXHJbYpfI1E8ZvAiLYvpR
m/PFKhSPyHCm40cmOjTMsRYTee26VYfIDWYTqUY7HN+501UjGiUgwj8bhEMcFAh3
1E5sjQsXoRy5zlutvsOrmLzmXoOeqjEE0JEwIMM1Gt6VTnK3MHBp/pq/n8/RBIpg
QiM74yrPRl/JnxDnnbYLACQnciz223UnBYIrcvj9ylVn8Ju/mXVpUKZKjBj+I6Sh
CPLzUVfcXV/3/EgDFu36QfB3+EjZd9a4OieGGsCRSNfd1RQ0eAgdAqfVlUG1YTmv
I3L0DVnBDvjNOrOyuhBb8h/4crEsVpQyif9TWyqbLCqsEoZK2auKi/DTVnKFMnda
4WhdJ2U6/TfTIRknBBDkQqQ0XMBERgAzc9ap+U4YSErAhRRZKkZ2vB0ACEyw7yO2
rRdwdmDMccuIJexFu9ZnNLicibmnA3fWIA8vq7sR4QiTR8W17EH03XuyuDtew8WA
2FUaz3kZmdHVk/uJXbYbOrrbgvQKz1Kri9bK6Tc2gCsI/f9gVJAVSp7jcnXT9QPF
qL7HHSB53zA2bJUl0eDsqpqNyZT4iiIF9msxMvlgSYR0LQR6oxynHpktHVzbDpbi
S2pmDRwZuXM5GPIY0cVxTlcAfQgHiDclbb1tfRyl4JHyNq+BoYojNLvCX67ClqFQ
qeNjoegXvqxMuD6+7izYnjpSM/qOPE6xkGFOLXnsjgppqeOiHS/zyrBYf/WVy1mL
5dlPTQE6ftlr7Jj+NBToYAHFjIrikUOYqWnnsjKhfvVxkjISLh3vIKnujrkizbeU
5w5SolVGPjfyc/vScsUoggDf2y46gVbl2ww7nGJdwmwBKtCHVXolE+0y+y+Z63PF
GnZoB0NrRwr5fDgDnaaFjt+dw+e/+7b2GJC9rNLTKzab+7YjL2DoNgfB52uHPL5f
fgzAAFg4q51tdTGnjhASwRurBYadiGH+0xWoC95GEYE/slUZi4dEw1UyaKcGP+lM
9p0MYtxBRJV6p5nY996skbj37M4MLUGvXlQ6pCnWOkrQs6/z+eCQ7bFP6Xr84zkX
5y43JQX0i1AIIq1NjcEhPlZXn0HWUkCdgmm0l7I3TSH/oXUSiRBIyTnFjzgCT32d
+u+vg3IG6KhGUDjDQdccY14O1yGPDLysx2+SBZbhG7UvNHMTCN9W2m08YLqfFphR
scyDP87fCTZZN5uC3tvpmB80Pz15hLeoyipvsTb/wK/KTp5Z4h0flTFWmOoveJUJ
49S5pEDqaNb2+a926QfNZYM5ZyXpH1U4bRAZaQ1teIqU/NDELqT3fTTsSQ2SXhwE
q1QxkEmToQxYUovunhkgPdvHZ/itx8QhzX/JqTOlulIxnYB3S5dSrmGCswWxf1Ae
rRk6hpnKSFNdL90yKtnL0jt6b0/Zn4wHntQ8G0/4vHLcIba+mzszQ/JC6Lx4/Xd2
rxIEFbaYtsOIOysaeXxGbVEJBnyVVR7zk/6JhZQepyGL07JiKHWswfE07HRPObsl
qKaTG7K8+Y5pCllRUqQNBfkgzBxUYdGOlvIDq8CpFKCD708lsdBkVm/ebiqiDtrF
1t6YbSi/3ggClOP1kLfyBo+WWRiM+qA+9nv76jbKeV/DgGFcKIsOomQYKe3B3EJU
00tVyqAo2g9GPtvUDD9TRYh86tSmBt/E4LTi33ZvVCVoFBGG8f7lcfcRD/bih/b9
LYryo5mjbarzyjvucpbRZdslT8ixSAnoMbIUo1SiMEP0lJOQ9aKoYON0E08Ifg2w
Ye6FZMrd79C/PT3yBV2kxkFteeRZUFg3gn2O94JyezXpW7p1Kgdn8F3GLvNCUtKQ
LeQd8qQIGrJ4Wy4mh/9LyUwWGySRWlhlcArQr42cVoFy7f8VaDDM7GP+0TaO2ZYh
sTZYVu9HRiIYPzTQbQ7mGGit9WOtPLDapajav1D6MRH5LuvvWGp1MZ+KtmIulpUW
+FmxYVK6Ps5iTd2hcvbaVPH8Om+RWLetXHYyy/77up0Zoiab1JtYm7ec7WBNn/+r
OojxO4xkn/PuCjdjOVglGaiCMqN02hsEg1synUNTz/LDddVWSs68uw9djmH6tdMU
Z//TED3/LHL8OddZSjqaSsk16GtnHBH0gxLO/9q8FFwE7LJ9gBqiJAH0BV88vmeJ
hLv4Zce1WHkdbnffaAEXURBsSgD1I7kczu2NYRSbI3L24zJ/QcghnmiozYZXoOlL
teOBAYKTQ77wU1nIhZl/ij/bV95KNP9crV3jwwbWZ7KAVYa27Usbr12CQDn1PdR1
szzKpBo2thjyOmCWWtRoFFHDTCtPwiaRFFqXG4/xYUuZJWFT7BC79jLOxcctD1mW
h81QXHd6p7txDglOXze9/6+tbD6CTWJeSbPk/5NViIdjJmDLJ9K3keyFg7ObswLN
vt5Fxz0o9Gmjxol9KNPgY0m6tcao4mY1nGC42jL295d7sGH0mqzA2S1L+qYa3MKl
zegj6ZwWmzTQpY5IJxV2q1nc970aeS/vGqASSI+pu3coZPVg5byipkASTixPAv+1
32Njk9XTN5G6EaqqIeZXmITRK69gdT43M0Y14mKfLyn4G3PFElRUKxJQ+h+VeQmK
2gDvnEgwYQ67J/xHiuxN41cWGf0JSRiqly0FrIl4YN2YivnFfX2B1wkA8ur4Y7wC
LuDEOpRvmuL/d6/xkKBR1JM6f2yRLV5DYdWtiaqvbs5fa2azDSAbO8zZCTNc45+t
2ZZl5VEF5q/x4GSnUVYk1cPnmdMUA4yGtb9sO6GwJlqy9CrVAD08D13HHKDGzDoJ
wrQe2K9lwAan6bAkG9PVmGh2OmRlTtYNCWh3bUAfwL0X97qVQftShaUJYUavPeeE
7Yfq5PoM8G9kxzqv7SEE5SOVRgnBF0K2X0lxR/NIQ6Mt3wtVqDdABZ2EqdBMRVXt
rh3USHYGVSy58L1wQRPzifQCvY64IT53klOrntTeXXmnCi8X/WKkAHoysR2PbT5E
+E48bjmGJwQrxDLlaJYJVdqT9/ebg/WF00ciD10f9HIVajr426wNxZf67Thuu1kB
JX290rrYCbPcvr/CsBSRH0F0mPIhnELqfRjcyo9cPxQS3g2f55SnnvTh1bXgu6Qq
EP01GluQFNhflKZLMqtWWd6sZalJBCwrZKTEqv/LdV5oWbqIebNlUtVXsNGQgkKx
BomPEKFY7X75sv5gHdIIyn7seIuX747z4ivC4TqvLLUPGZa9lYKmdAKGfC8Y/GDM
tLKcKGm2Gxrde/mPLTpnUsL5N1Lbs/qUDjLYuSoMtJgH3RKPrp/Qr9iL6p36wT5n
Cv0zc+yb69lJb0Vs2QyGHHpwPwDv2WgO/MhihnEICzisDUWL7jgEKkbdoD287YCO
4+44wyJHsEnnPrllwJb6cquOFgLcdbd/TXw/zxN3P9oJVa39RbDD1Mc3rE/5M6ed
px9hMTN7EYZGe/g9EJ+hcbFDdG5a/oEqqVyy8iCrzWMpekCKJPySvr7y69s3/iIo
ZNH+/nNksqHtB4kX9h4s2SV6K8mMGqbuPhQyn/2XWfwQx1vI/X1DQMyy0gezFSMw
MZkfBX24O44U2BqkB/YmcMdDPwofYxs3vzPddw6DPzLo5Wh/Waz6hg0O5eBbuYqe
fjqlPx8jnTZW93/d2zK3PYfv8VqZZsJKR33hr6ESWhM0ItwYbEJ9yLkX9Ka6uTYL
kSO81oxppCgLuwuVpcjROgM8CTsNyAlf7SWyY1T5ZCMiIutokRaj3FNztL4EsAiv
nSQ0UM1qwzwp5KNlqa6lK1ab3XRvHS+Jw9cefbxj6Ic1j4c9400lcdDuHA1O9XpT
2phlwXNRSouuqnSeuZEEaEvKhsgo1I+lr83K3IrrMnlQNmZrJeSSrOw7PsMPLNAg
r/erlIuk/PR8Jm4TuNaS7n/qTLBGZtargL3NljaD3NJ9jyt8/6ZMXPM02+DTaNC6
7WWoON1pOmgASQxmpiMj2VNAiu9PSUzFWLuGcbhbWlpECjnydi06gmdLrZHMrT1C
zKUAuD0zlXsaIH9acAKPl8cciRDc2xhffIVjQzkmsrgcJZBZykkdgrI3itzlKyV1
odxlwa8FOHyBlSOMypOdyQu5ML+ZjZwS/7URsiV2dm/pFAezQhq7koX94PnMoKe6
5pQzM2397CxsDaLlzQ9A/c2Gtu2BnmrAE69xVPKLJCoE7Og72av8lhnxI+T8A+/Y
lLlX6POVZu89rWrwpV/uDdjv8l1wjoGePy0KiXNNdCZF2hg7FP5n3uQUIhjR6eGH
6/XTPc0RwDcDLUe5u5MAzR+BKGOoM+Qqs+fzUexaK/LmSd+RqJarv6UUBD0iABdH
UrCdVKPeb7oR2OEaumNOIowj/I9hir3QRmB8sMTcZjnhs1sqwPhyed3C1gitSiv5
pq0Z0edzcxqUcv85BF236n/8MwlJgdf1j6gjQdBGlbmqR2SAKa7BeCXW1Y+qnKhW
hctQcPnTvB5gp1ZI8AdeLwNtsFQ15dHpjU77lZtBzjtfSNf4gd3F6kLAQVG8NnYc
XYC2eLggX1rJkWqQQxTKUzSjaFvZ729Z6w3Zi7FVHBVrNx+vyaisMSSq5gJG3kUe
aUUXsn5S2fhuP9UYM2QfyLM00C1lozqUyuzZTTg+EYkUvO5l6sg3eaBxfK1zS7DB
ZWdGtqOU+PuaNjrpssfiPtO1qOdsYyyQ1/rnJpw8802xnDKqmVUPWHDdmkF6MUwW
N940GBN0CBrz9jgLlLlpRMNDql3hq+DlTxTu17FZYyYwiNeVCEijdFWcqMENcZhj
ZEyyApPeL3Pd8uSB/Oy1IIjTCTaCqs2s+NPRJiUXaPgCLyrw43deT/2kOndzBSAx
CX3vv7GpwoeZS+jAw3W4S4q+cse3qbwQJltr6Y+PZ3qZgAou0S8FFymrGX+DL8LM
jLuQkWAcu2HSf+ZPkri0Bugjbowpzu6foFJmMcsWDy2FftN8w62twnNYPBgYjB6O
QJNOe+JKvZY3lCU3BfNTRrPLqbzhpy/ncLZBhd89c5/faqSGAypM0OzqKgeKheFs
jmDo9lvs+RbKFHnqk5ieu0wP0Z9L05I5r1lhKnzgzkVxxYFiqA5sP2Kb9WHSf5H+
o8zf0YLy1HE/EgHvELTVqhq6elvpsnuCYRQB2q2xxOKN0nQlIloBKqdJJiI85iB4
RetE4IqAehw1ThavfKRTVuFDR5UaH7+QYUsrHyAQRu41CSBGvnilwiWNfrFmMAUR
YlraVH33aabMRlOJCQXTiVJVimdu6yWJe1FAMDJw1Eoz7WE5v+nRPYyJ/r1PuYFb
vuAaOiiAtF8DfGUH9huM5hRKXXsGE2jdaGfhuHHeIzeVmWDdZWhuIXXd167Zk8oQ
S/CJT/bNWz5DXYXLgx80tI5oZhbxji2+aGIRwkZyk6aC/ORXT5I5iSBiOgNhMtXG
2wqt4KXIZEVoyqckSy8Doh8qHc9+3rOy8FG+CfMD5XP74Rh4CUwUKl1o6/9CR5/q
m7J2cHFKnpehZ+aZ9ujirAOm14sH64pcrPbTGSr9IWWJt+X+ySmjFyxDC98occCd
EPUghb3udHG/8/q778fZLJlGZp+od4fvK6hNh+cSIApD4QiyX055F14dQ8UWALaa
yshA/oIjcr+oK9HtHwS84iHC73lSkGUpPMh4dvZyfUq+Brhb2ohcRGUEvSmqqfFv
imIV1wJllUgouyr17rJ4WD0KMMVaDCapOtyCW3tyzxl2oIaS+w8eFllhS47LeKjp
Xk8TAWpCnq8AhxDFV9PB8buJNwXVRMbPqFr4Zs6GUuvH6901KlzCkjBPqCxNSBvS
DMjVThEdc/RB3iDpccaLvYIn12AxRX1tmwN6ZW0+yxid05klMjCztE1cyMJ8+r0o
nplsyIOTWyCLtxDZClW5DQxmrvJyhGiV/Zo5uphgsZN4GoPp/ItatwZ9UG1s9pJk
GI/KIXDDKeDK1ZnHA8cCWIVGBNZuCbDT4TYoB5q4dp/vepP+aONuM8BxrW+7juYN
eAiV1NytqcWQCFqj3P+2FNqBeGWcQwEAp7jsQ/k15KTCD2C3i6+8mDyhua5TmJ5W
eJ+vMtSV0gfoSORhtZwDfJTV1JBrX1HXMpwrguQLTkskANrbaiL1LljL/lMmVpCC
G5DKbKUkQZtZn/KIFS1zLf4JqtV3GdvoXlFvJ2lfLLB4ZLUjkjunFV39KcMwz5vV
hCDeclbLK7NptMmO2qEMLj0T7DDBooDCR7pifhU0xgPRpu/65raGQpfpsuy4JI/q
KMYpm6j4bVVofeD39bIlVUYV2LKIW2cv5ZzE0viwkgtgHjg4mROOFesq8WVrXlFB
sfKmh4rFOkg9+DT2/s4yL4z6RnLUVOdTdBnmlnuXQcWZDj1DivrakCOXLSAYCtZO
z96x5amrHr61BUltT079+I9vls2hpP4ctMGg42/DlU6XCWwvAVKBIpPpTgRi9Wwc
RQbkN0FlctGcIVkXOfQbtt13Olh7LVg11YCiecW/0AU17rglB9hU54CW2w6d8jhu
jXQcup+6tp5n2pqNnadyuABAkFkP3M8sq4QxaKz2Qqe6ym1S0kHA94WT6OJ5kQJP
95JfbyZn+5dZPTi6HdYBDrJ31mG7LpINg0s12dfljt6z8TrZ3ZeiOe9+ZtlSp2gl
E8TdwJooX22PAiFr2K7b4Mi6PRZzNTkudZEKRyJUFMSObsqZWUcUselM2wx5C3t9
B8GVra2o1ztFioyabjY30wBlsjYUUSjJpvQj4xD43uf5p3m9/631W2LE7gDL9y2T
BbwUnhjp9NhzXMR1fvtN1il89yk14Vlv4mtupBsnNiZ1l4S4Kmw7wcNH9JCwAL76
7o+5U2OXDkyHBHIFQ0TveduaJKf6DgUQFwdNnMKWtg5YoJ2dDZfVA24qJu74Fdjn
QBL5pG4OFxnfsaXJHFm1PcJMTlAsad+NMNRKbbeAFY1Y9Xy57q4YHFgAGNHmifCq
ufQomQOg+MdMIzu4i9Ewq3S+IKYDd6uv+3gRqWG3jICGbjuye6V3HqWqRe7kbtY4
db0xUOfeIoCTBug3lTmiVeZEH2Fm8kkPMPX+jkGQzT48umg9XgSHlV6PyPF/OIf0
O3CazJjv+EFglUE/byXFs3dpKeQCHHnRyNCHcg4YJotCqokTMqsyUqzbYVApBl3Q
/Pgz/K4q4FFFbw91tKrR/2s3SMWO9AYyeqW/RyrvP6quvXEZo/X8osdsgoH4vdys
dH5xNtkcLCgHEZu8460U9lBOKnNGWAupzNx4LLO1Z6tSs/z+2YBZ3xjrNGozMxtQ
hrmgoUBGvaHZ6LXMDNcT8L56v7SYq+Ovr2VD5BioEDzAhICTOB8oLKNUL1UVETyY
IQ1Lxhobe+rh0dPvYKdU+t5Dz1aowVb+ZRNy59NezCE3RjGjyXvSCWAQXW/ChCw/
FGud4gzaw181NeWxoB1p4OzF3lCak6LaIqMXtH0HIP+GRKNDVgphvWTuLBb9Osfd
0GgoqBzceSoqu38x4eFDcM0yxFbGmvwg17a19t4x+jVsN7vxwKrS/vJHAzdq4Ix9
Ot3NZsDKqtY1CxrSVqVmArmCzZy+7/mEmo0VPY9r/Txgi5O3RS3eeCik5kIQntDU
Qe3IGShxXTcf/l6/NAEyj5UulG6ziT1w89M3FQW40ge+NlJxA13hiH4E+EUI8sFR
nR5psr8I4kTut/0LL/X4OZBnY42nzZ9SByWWaF4zOEsV60jBYeZ9Mg1ImbqsgMxq
PuwIOgdVRiYRtGt9WuokdDxmUFjFHEgI9GE4Gx9wFOlSXmbYAB7zMT1ETW/SBVZB
CVWFDA1tHBREQ5A+U0MxwdFU/LJ2Z3txAa0jqef8Jj/XQGtFMy6Kz+TZrIJmmHmb
NVdkJRAmVYarVz/211CnLjDIfyHKobxAucTr4swS+TbgQndD+T0owdZxDcptNA7K
D2M9LzIcbJKn0d9IjrsrUgKyoAXUX/eLvTzMzKQyy/gtJTNXICGr8bvRw9gv6pGD
tONssFqIvXFFvK/KVDV2LDZdUsPROUk7G9KW/u9CqsxVti7r4wvTTvQBzHLIpar1
RUwnfJ2QjnLPVH2rMzfUWnl7plQ3kjHrLka//fIcTD3us/EGnCD5sLVkZORdeQgS
i/BatUI+4JY9fQUdxelZRz/I6Dt4u/UtEbZi8M1wXz46ehLefBfvl+JrPTyiyGaX
NLzB4NADFnLrx5zWrZaccwjonA19e9hLq0NG2jwOIax4nGmTKv3z+OQz2Iv06Wxu
9mlr1ESt57bi4EE8pmUlptwtR0c3EsOh19DSBf9ojBSTKaIvmnnF7mgwOMgJNffM
bR9xKosWr94qWOTr1PrdkUDU3lQ+bQpLUViOYdCQP74N9cTQc/aV6B6b6do2j9Wy
nztTMZBXOdKbriLKYSnL+oogmZa9/VnIs9HdrQn0zkkC2zUT8rtdalzQzj7jJ0pR
SCPazQsQ0RIXP45wfaJG6qK6JvM2hmK3zJIgbyFBk6ydszEXJavaiWEq+2WeCJv9
Td7qR41W2QpHnGFGHvgTQzm0MN33TA1b4AUPk7nvRcedBKPp9HW1xWHNEplr/cpD
jJZl5vC/LpYayjGYB+7/K3HCZ9o67dtrX7ek2X2owbiG96kczaJXIx8MjdlaYNfm
2CDX+cFVTPNaP0vqfs6aobk5WTSG0gii/x16R9klwU8Zz4lPMf4rJiUVoLAH4esq
L5wd6X5RwksDNRQS7gH3mKUrQZLbtxk1xODxWFILZ0wgCQi2zJXW3XfDMsBLLX7w
UXX9naHvbYik0evj5C4nnuVbpm2j4lwmjj5NQBNyDt//Hkum5PLebVTJFeDYRlNN
svV8WVTUP6wcRyckMm8/pwvn1KqBplIGP9lq/hoxQRzowuWG9+WMjCkzhEuvMim5
C1kzXFUiqbnFGGOZaqdk6c6m8dBA+0NdHcxnYSfsoSKs1qA2NL+TdbKCtLaJRc8e
rTzALM8YrCj+AF9G4fpUpoUja4tKcoAv1AOGxOlSm09/z1p4+o3m6XjXzhtyEe06
j4ZggeuyqRK0rnVtwX1EDF+uOqndw+T0v5NJeXnkry2Y7VgHVF+TzXYmaocilwvG
rrnlDvDZw9IA0xSK2Om4hOEM7LoUuVmVqQA4JWztNbUSM2elO3xU8Vu5fAD5k+ma
WniA+CKw0AIVNQeFEdUHMoQux+C502PvrC7+byNoZeIYLYQpELKehING06oCjOjt
kEKqOvalutF2YPvXznA0fDe5thr5mBTHE6QTuBadQz6lO47lONHqrZIUwx0cDu+5
79s4BUs7ZmZDPzv1mwhJ+C2/EzUaoR51Kksk+nKxNVYt8RzVIrMGnqSUm4Aq+laM
XSfjshIB3CDX7jOBTduerW2WWltfBl3Yaj+SJCyqi0g8QwkGptY3eHNze2Mzja5+
YQ5OzyQIQrm3o2rLZabDSNHIW5WeVlrLFVF6cbQdXkACJp/wnUJkiEBQnoA0VQTs
5yfxwkFJK+g+rvxBnSHTU7UddP1F75KqNbWDZLG6sVqPZwo6qMCywttm7YJPk7KR
m8SF1sd8g9P7dd1d4sawGMGIRO2HYXAZO1AqH0gK8dEYRURQEWZAG2wFnyevllPT
W2t0mmMY2WyYfcpiQg5bW07J4tXrrAulghz7wimHrJl07ZajvBN2bdgtj3cnOgY+
w/dcunYdxbym3XEUi0OqCEpoTEfcoF06cAFvTCi4THwxiHfW9BQkNrmd7ZDGULJu
zs4/GNB7bmoQC4VdO31GjZYpvRQffpCtRkPPCP1wu2KmUbcSDbiGwFjZReEwP//c
P7+LviAzJLQmY3S/CrLS8g7AHfzEo4USTHK7pX9oXmTHN8gun2XgYefSaYVlic8C
7lgBRZGuWBN96uW7r7nX5o2xRD6bz/25CYoLBwjuMeZeGbC204cy5+czsrVFKpPP
W+9qn4qI5UH4n4IfOHdhfKO4q15hbo3UDd5U1BHKT9Oeih/bXCFC0NuhWMvejmQY
zfOYDmSPKrVCKbrMQkk3SFd0bSnkL+JEsnDy2VNiFfTsFJoTQpWtTHFT7gXBplpf
gfZL2yNf0vWsH0XMZ1rNwgTnKCkEDjkY8+vRTMC1j5qDTeCtxiu95e9A3UOgWhHa
gjD0qshDLXImW6PX5OTMkctc9gZP0Z/yzMS9s/oCuKnFiSub8jWY702xEdEMulI7
l9LeTVo9IqFtQIa2dp1Dtm0a41ggSskL4/ue1NS56BFOcjzICIFsRj2wZZpRop8T
dApmBEeyM+lMrJnCUFtlyTn8WC/IHL3yizbik2n23V+Glc8amUVOPwvqMD8WkjVl
RcPy55AY2c16QbytioLw7ctk6mZzXvNr0HzWdnp5o6aPP4obd+8A3CgvD4JXq/4n
z6xAkYbpqUdZzkjZdHSWp7qaYMroPQOZmk8UJPQiu/U/BEo+Z+cI1dAji7jOwokE
epB+pFXVIenpz+2sw11FrGx18gg8naEe42vvItsn1pqiSnoyr35wbObfSSJi5O7m
FLM1QPmsjPp/I+NWtmcAM1JFW/INx9/8pXagSxy+gwVcSmZ5gyhbwljeVY8Ej2tV
Rp9Vj3Z2TXh3cG9A3hhiDLFdcMEU2r8flWIDiqNUoUYwHuRpO1uWI0m4aISLYlRB
ZNTlv27m/U9vCtuayKWyFot6MuhHisoBALCsxA0PgzR1/FX1ugMTW6ifiC8kV4iD
Jv7zMAW/6yzGEIASUh/Q+RmATPLpVwT2Ag8IjvrAxStEClzPsQnOu1nQD2OPcRyO
vXJSLafOYzoi7c1iQ2aksThFonq2A9Z0BBsS6Csoxq8dAIMwRmbd7M5UaYYn5Ass
tbfN57QkrMkGitm9EmUDUBqEylUyHZqFzfmHCxxkJ7K8cZPKhJ97dIh9q8msqEln
f6/Z0fzDL0xbUDO8N0HSGByhPVVSrBSf6RWc2gPYwg8pedFUOIHOuynrJus23Xlw
EwH0arttjHnR52L2OU8hQMMhimmfr4ATtDucphW8aQvU4HUYoRQDP1Wotld/LHnl
E+69im8EaLV6SEeRRYqMFpg+RQIzj2gR6qlCbVcrL9NZxKBv5Q+34BrAUGCG+yiv
m3e3vi3a0aFxX8w1zIu6tCF5tJ/lRsrcrDgHdO+l56hm/JLfvIKYFW47QZC3/27z
K57tn0hJ95V8Rn+G3fI2gQqJrCXWgbZEEC9aPzr2qWvGT6Ble8J+Evsan0aNqRaE
ZlDLpjj9UGDhFV2eW+wsZGi8Gkj1g887pi90MuqIPhE7bKF6BKGi7CS1B37cLZ8e
FrfU+ORUrvxOk1+V80uoDhhLROrrCmzOHezjfMIOdhu4qxMOQlR7flg4FDX+1Pjd
9ikySJB4bmVmuQwrsnf9C9vQ0+8cuVkNWJOu7Ru1uUl6Ow31ggWEXURCc/VGTFxi
HsrtBq+Xisd8bZhEKXC3D536yt1Rh45oytmAGqYWBAu/WBMH+y7M0t8CUs3qDhMH
eqmBuhz0a1u6yCgVT1/JgfWbYqnXdyAK05c5hPKyFpCyZkmH1XTLTfigOl/NPB6b
R0Kyj1fBE6LufceVikErxO6+DoCr+DYZjSRklCrQOpsh2a1CxsIC0HVDkzxuGj+N
Eg/HHZr+tcFKz59bCic5llSGg7ySnYK7OMSByAkmVttynZ6qEwe2cyGA55cD6FEb
PR+beAicZeDaB1cMhBp5OP2hsZlLMA+jIsOGL97/ZjxfPyqo/cq6eoLeh8TDQkmG
UJOSZuFrCEaD0nEhmFXqVLhfQFx2gbj85MNkvWtENUv/4QiKI/hHxCOwsg1Klcyc
I+3Db1/gEiG/bIdQN1y+KVbYMYOy7/XI7Q5JArBV1aGPcBeoxUF3E7rX3U0cf6vR
0kHoI2ZEKfQAk9KihEfMtvk7pRhOu9EJ0LLAmAGsRTjIKfqUR+BP93f7R2Wj6+Bu
Qm4gQCYWEDlkZxfblGmuF3AHKCdAjxIDKs8dnEtPJrMG9gfQP2QQgUa4cQVkt3YL
hOWrhKRVcNdJ/7uphLNrxnBbrFYCKbh6zrbHeKENDVPbAXQsVYy7oGqBlbWnIYrW
ua9m2Gc24eUf5Khrp1p1wxf4Ze9PXfslCfKBL5gfilFptpPD9E4yMmXGFaWadpLY
BHdl2gM8LXh/q0iukN/hJKwC1UTYFw4sv0zXZY4JzRft4aov/IYV7+8beUcKVqVT
Rl/asji+xt+rgT6yyiWh9Miy1WNWjxFNPe+hCeHY8ndHnDdkhG+2eotuBeF0gF8S
LgSZiMQRuSDekjxTy7U1l5ZIL4LARZ8H4GXcD1UAzhJu1HwlMqLSwdN9EVmtFQsq
GXKcF5A4iuW6F4ITDm7GIezZl0/Bo1O2l09xeljAew3Uk+3sCO9qqTpB85CapDAX
ivICtYSkdm9hvEl3YjqTlhCArY7BMC+sRVyOlhARUtVUZ81KFWY/rM6XgOjqxmwh
yyRFkhrDn08ViFVtsA+g+x6AzdqoFaGn3jXiKXN9W91MEU0RJo4I54PMMAdig8aY
p7tE8FD9sYDpJOoAWroBS2jgDTZxGR+MvqazJThcjcqxc64QChl7C8EHqyewJVk/
30AF3pkADD6DS/uqFWx9kQLzKbGtPCMppgVTHGTwGhTzs2S+6DYHo5iHuiF7/+J7
cmm6QbNzNHjCpZ7djsvSoIf5j0QItXIDbv+1H7uCrCrJPwNOUS5TkPMNlPmadFLw
/TxDYzM9GueTEuYhSHFX87DasDDdbqOI1ICc21QHev9mUtw54h57wsUDbPtlBNJI
GANlFzJFXUPdjmQ1dQidR4FKUgx5cYGmHTvVxPelJm5Ea+53l5Jbec5B41bPx1Ty
TDVujva6JCmQFJYLV47X8Xk4XMjGvD/Z0hjuQ1WsWiAOLWgmyLoqWA3W2R5Ebnna
+KlH+oxxtUayB13D8p45FG90fv85Fvp2LvGi4X+qndtf9XLSom2PnouoBYq9f5wd
QL1XsQicFMoz2eabL7jkEto/XZGZf94RzcLVFREgyjBOzWiaPEQ29m1Jn/xuUnqV
iko93rPsKNHIW14BV5GoU5saVYJLwAmmn9l872SQyYC0YxABKJG3RAxhlJmXkW9d
vMM0wGHksBWhgH7rgnmzh9UIhMLDulpFzrret5/zJTHrF3GchFCokdIlV03FXjeg
wDlb7z/n4HdPEm1oJPLqnHYY3NspCI/onn5Wb4LBbxFBL7YFf+B5lf6m6vyV2Bmg
pyIkFz0nCFMDPfvni9582bUFXT/V5oYjWz/qrZEXkGI8LbO8o1pvV6uGTiJhgFtw
qjM9E/5s9Q3+9xK3TgPRz3FaWu28Lz1+75kSfXlp8zgtEC4pdhD6XMir9b7IXECN
U7DR99l30ykPWisb8gJ00IvmcNC2KM+k1hIaMaQIHSIPUCjhYJo+ES1qeytMFTK3
fIIdQl7pi7oZUJ850tPEJ+g6fvBPBretY4f6AZXNNFE1LFlOrhlAq918O6FJlSUW
eFk0gF8YtkwuLPdNlqlh3k5Zyd7kGa3sDAB9YYydA7Yhh57bNDus+xZP4nczelt5
YUHZ02KV8/pCt8S7IOsZlLhpmtKnKJJDVn27yse6naRSSUYxPy7TbJwtxzznlq96
6AxF2fbB/PjwsxuD3ixL7jxKXRumINK/aGAH0gX7q0giQVzAyfrE+l7NHgf0ubz7
0aXwGCixJujSvkXzheRhlNosjKlRrkOESub6LwQsQ1CZysd9odPvOAX4tpvPR92m
OxIDhW4JuBU66GVyOVYqm9Wiqq+TUfyvbTVI1ebBICg47gd83EKpXmeirhnM2U1A
NXu30pBGckChQk1GPCntFX8ZxAY27uaDoHorbUwz4Y4pXByvSnDF/GFEuxCZTuHs
ATmW/W/6ubdqJieqkrzFDPZkELVhmpseDrmtbUDhwKEDIxuK+CDYj969RfZPB1ya
1kc8FKFmcUNAV11Nl3ZrksYgUufOlXsama5YKD7meMkmTmw7yuCXMO1/UzVaE8fi
GDUzQHqf+Pw9D+nAYjTDo1Ek25QniTLR2I/+MZtbcYiCMsNvLR1HSIJ/a43PxAar
3/5endm4Q4EtiRGQd90UL4ZZ/9Ugi+hzHIAFJ838xq5gVDs1CRb9lX9a5HOoFTe7
mu4yT49R0gWvTsLxJEdVTM7GxYlVK+LuTYuq7MALYqPoQ/qECX6CbH/tzANBf9EI
WSj23o7SUnLdhpHqG/z7L7OA56GR0s98v4HL2a9CR1CZopTL/QUYSxRpEAE9YjZV
VPVVusW6/ttU2ak3puAsMD2iS7wX3OUCgrarZcnRi/i1GZKfbI39g1fFWq+ATFca
sz9Uzd9jTns1MSCJy5hF5fNS8L2sfLT/Xxfek3/WxFFU6yn/X8eHYZPpwoBcZpSO
L77d309Iv3XIXRDyIoQUd27YaUHUkBWXyGtKd+BmDwkflXeI6Hrrr/OvhqNQlcnT
htChENcwyh2Fs1PhcGMXLxlsbO4REzSkMPX8LSWP6y9WnjXvqBMIkuVcZiGewT4G
n2BQUA+rhp+1bpU1TpTwX5QjoFrUgY53y4VK4wuN2eWLH+nk4RqMdpgIt3Tbs52w
8z9W+O0zXtPn1XsSjW+VFt0wZgjc35fdJrWP+lBvY9ArgmKLEPVA+kti+G5tPjSU
J5e01PmDYERAWUE9S5w+FyqyZin/zXgJBllq5L52aDyN0zEgoCDN6FT0AXEZ0MIZ
TYK1y2Va4aUEArF8GwX+lQnpJIiU0GS46RQbx29JkfsU3rAaqj5JQMyylAEqi5/m
9/OMkDD//rR9Yj+ZzvJAI+RpO05GV2Lsy54zHUH1+qO8bWJJFizypLN7Cuy4o2D5
UeK/ICGklks9MkdTm98cHsg54HxSZfJSGTG8bcpLrWz++kj9sFAolFlKxilUuCfq
yS6aJhf2jcRlLtxkSBB2NW0aCFnzHhwHQjsAYnLG9v8CrbUnrYvG5+osSA0U6nsm
olojCBPOqTWtE0AyeoiQlOcyGxbW1t2zJ0KETiCfbf62p5sOd/EN88F+HvE72rz0
vVir6XoDO0x19KmL310NyGG9uwYuS1323+DzcJ7Rihn+/PK/vilEGh4vScZzwYnC
eZwKlSoJfq1yKhaEObaJ3p+ilVKS2uAkU1PKsV/xh3eXqpkFdcVk02zcWqlkC7Af
U01DnA7Hm1jrIZVBj3vmt2HSHWL6efTcL6Q9KEg84lHjHXoFUdpoKsbjmHFAuRdz
oNXC5BAlLidtHTXs8BBgPewLqqOC1gev3dcNpnqC9Rj0kIAvsNTFJEwC0bIXJ0XW
ztD/9dYhzWi9dnRSgeTQR9/l4Fd0mnckUAXvFkrJs0TYQ0FF1nL2baEUa7r8mMpn
HFE4ALeQcFzSZO/yVcuSRM2U6rz9JsaE7NbCv4bhZcL3BYTStFWdEIPaeiLNOEBY
uOBDBqMdbaxnZNefam14WRLYHxuoJhEh1o3mIRak+8E9NOZWhWwGQxvO2qHAxK5l
/tZ4zIppQa6Dsz139/MqY2of3WMS8RHZ2aiKlqNrtxcDz1CytJXCG9YVtFoaavW0
UCoGEN+k7qKMCYbJ6IIg6ImwtlND1LofxiQH2zBAAgY5t9V7WJMVonp9RZ9MIHMa
ZRgt4Kg1/1rIiW+Y4tHvMjeBkiKYTHsCJHy3Ba+YGfsve+Z2KOdLjY9MidV8JAkH
emvXbiqxGuSkH/m6Eaasf6kld5C7+Z8TCYqOZuE0Tj91jYawTkq85Ngc0tVmkBxz
0gnd9XOQJHU06Ak+4xdaLz+JYs8cTRipPhyPMih5JJEM0x7ml7tqTK2N2jb2g76v
NYtT3G49WqBzaqDnBdQAkku/8QYwZr43XEDLsKwgXT2xaAhQE1X6wxjzrxz0T30Q
X8MxzX9wtNOvrWD5lHyqQlETo4LU3yYeHYLJB9GsRtkC34oaGxQA/+rJXqtMx8Zg
rYl3H6eRjmw8OXGliusKjRvr3brZaXnuEHzoy8nzrEFWdU9m0091xLkqYLJbUhsZ
jgkyixDjoBcMj1bTIFXNREm7re26XwLq3Ztg7Tu7wVV0U3dTM843ZtDcRyI/xDAs
ZdW8Ck0vHuAwRwESq7TW9paohZppnyWOHjJwYgF21BqkLNu1+yey7mceguzbEnpt
lA+8nrcnK0pe1AMQo4IJSvhhl+j4ZBIf3uyl/k5Gk+lXJT27bzpXLXko7GGX88bo
tTXuGSIN/1IsOpgHFtPY0Xldaz61TMnGWjiv0RuVuY5YgtvI725/OwvvTltddaFJ
QfVXWUOS+AQkYnSOrP0YR3HBkgcPYuK5tbVG+Vl2OC4d/RFkiqGoAghM9po3PZYU
Cow3TMRcAoWjmCyyr38PpOMs8GAW2Piq3eDi0n6kS9hXfki4TFqJfcU3xdhiZ1kn
vpE+Um3ajXIpfdoDterQSDuIMm8l3q5xtRz4lQ3Do1NUBUFDcsNHk/tRFdPjz0Fr
ZXelRpxqHOutpWx5+K4xsGcQzRN9BSaTp5k3XYAmReV9GbewNplYqCMNz8LCQROa
xMRMuKrzb81GrMg26UH2lMG5Y8HPNDacN0RdO3Q19Pq7yQjIkmkApiLaeqb6hoKN
PVc5LNZVz99HJWAx2c8g1fegTXtZEyhn+P7iiFqAi7qeZkefeKfNKOavzceiC8Mj
8IbFtL3/S/msHGoESggVEal2Y8ZgguWApRyCYa1lwptYJhhIQ3fIbxaLcRemP0vu
IO/pcv4iPrt/mqoaLvyEpjJ+IugdSwd3KXaYz1fYYKnz/IdGYOXgiMh4PG/S451E
lPCoaOWl/WxwPDTSzUBv1xi9Xg6UmHCigoamqR8t6BV3nAbo38/66dCnRaVaoioY
pG+XEjzIUQvixoo8i+MqSqdB0xyuJAtY5ip7yZ4G0s0R7pdGz21LJOf8yqi/Kob8
knJ675ROVX/ykRQoNGvD4QXTcVdyUrK1g2Xya52yQxl7Ky07k8yCtT5krbJ1EIfq
omy0pKHfiIrY++8NuiHDsgYbFXs3gqgqGdBRkGNLMyVIWhXHDLAd59joDqLrM9nJ
NZOWTDddS4cODgqVfpV/t3wGWtTX8jPiyn9zzwQIz+EtyHrt/Np4YDtBn9HSbOoM
6VafwYFqGzZ8MoVHHg/URySQgxE1atuTNzsMTQ4JC9fdKQp1uAohVdKdbwS4NYPu
kRZM59pW8Vfeo3H8t8/itli4EOBmJQEpq9qiV7kQ1umJvb0/uC82bSeN6i2OtAV4
LpA4QjIiOqv6K8n2MfKt1/nZ/MjMvFLZejWF00cW91q1HmW4Y4VxGJvwiE49J7V8
MSvC83nPND4BU9LGNVDwi28cI3bDDBoZRQlT0Lr4PczTphHyCdMxMevUaY9bqUMK
1jkX6tngUc69UblrcCWDi5iULRvhIBoE8TqoXyn7LBu43t09qNXHodpS51+/fMXl
flJVh/JlOoUGhOR9Iv4frSEZqJ77u7NGJtt+OqjZKskNSZY7zYrPp60doO7ghSqi
lD6leM89qzWFc5JZVtreizrFf6DjjJ+5HFHdAs4HHxQ2C9aXtzvcIwrjH70dy/KV
IBQ+IGVuxwp02cqnKKb60khz7cgTBWY8EpKQ9kPWuxowLX36plN1YmsGFvN6NXsD
ovhLOej9zO4I0B5mzFD4EauHfhwxcPTrr2fACybTmDIm0MOQNVhne5GwYgCtoWMZ
nRAJjd2dp1IdjMLwbfluKwJDWp/5vBIPhPXXhd2eNvyptngmED63Ilqp50y7DYLM
vhQ9nQcDzc86eW4yuUByNPaRe4Shxln1BLvnR1lIDKjlZJdStjcFXhF0D2tJLNv6
dosETnd7wDkXon4qcfASsLfP19LI8BKU3cubAZGX21RB9CGFc7yq/iYE54YsGm2u
dtDynKYLRg9xxl2GyX4uM3yW5eOjODUbDk1W8g1B4HRk1htv59221MMrMZxG633C
f8DDsevJouiEnfGx41jKvyzACsRCAgLbYQgnwa7dU1GxLWMybtGWcP29S6u3d7v7
OK0ys3gXPN81YAZbiQ3nHTyKaU0BZTvpFLOK8vNsvCBPsrRWvX8OD+fOLGVQW6++
6gMmOeKUlTcLDQiIPDjqOA9zV5mUy0e/cKRVLd+Yt7pZ/snCcAe+fepFC/O+7VTz
SFntD4cJY8hjXRWlUlIAuSHffVnBV6Zx2xqd3w5rW2NpZC3p/KHWwcCSYH52sqps
WSbXBTPogky/Tb+lgMfLE51qDUT4LrqP9KvvLHnA3bCR5rpauyXNoME5fkOVs/40
I0dgPMXrmPKxcszv8FbCZmUdyCWiWvnsWAuqkOe7MZjDW1PtXWq12G1KUqNgLkcn
GIVa5SgLnMBXfTCJhJe59ZLY/QmjrY+z04A2vN+K/Vec7LgnUqx1nXtJeTIGo0Qs
yfU8cNU/2gc8zPV97VkgnG+odOACie34/2JADl0OiaPZgT7YHAecYXPTz64qtjyK
01HeiUM+ay1VXu7GuQhimjzeP0Wk1w123B143Qr78xc+ZRGIA4LY56mnwlk+BqoQ
VynABnI8OZ5CUI3r/mOvILCZtyS0yCsiRMdZJZ1benNCc2nqW7TvFVg20uU7395a
bl01hh2Kux7NNfY0wfYbPuopPtOclW6GWUtsoGewiI6nle+E8PwJYV+2LWx16LAR
I3NoXPUM2Q0ACjgZIhKB8i/awLL704o+CpCxiUK5Mxm3NTwWunI4XrWlc6hAzyP8
sp0T8Eg3SPUNu6xu5aQnouchtpBboEEhd4hlSRTlELEyQ6sUB9kgPcRAMy23a4Yz
BYEE9CHjjWQAJiJ6XyIAFSdnQpxBYS++bZboQGktcIIq0kEV1zKUodBFf3uWxXyi
6tMehO+UvoJHnz9xJcaUl8NI6CbaZ7apGSnz42BUtYzfnLvxONeHqHGNweTQbqJF
+VYk5gasQyMabfVvvJYJhWWWcFFnAP4eslZcIuuE+GdBiJhew4rVLA+jkWOf6lX/
ET5ql+yxbSyyY+mo1IdOWiHnLt+mfjWmBj6xCeS4bXFO6o/Ug66CFGARyo9TPUs/
3waZzvEDSKTVDA28B+4PCgOWxyNdnTbQho+yqIb7mis0v6Qlngg5BB60jGTmMgvx
bq6A4fFPJSJlUNJ8cFbQzfG6wEU7q7D73z5ksSG57hJbRSmIXuav5oo+nhTqlbn/
crPEcf0gj3PNkc9I1DHzE78k+LDPftQJwwQTUUdPq2IcZBF87OFh/Z4H577JS8sx
i23/hEa67MKvM3oXstBH0Prg8bsQqYBeyHlbbjBfWulgTFjew8QEnJZtcM0s0RLG
Fbk147OBtBD9PkNxNS/MaITDk7IKxqRSqgj6lgVw0ILcEZNSIjV06MUbvqUlPZV7
0z9+1mqliUDUahGnWG5z20iwA3MNG/ZN+23NIE3WZoI+iTvwgcd1tCe8QixHP34S
NsddPi/SjjEq3JO+FmADx6ewiXKfaz008iig21KZSkFwRFHXwfr5i8Dd/CanYnQp
mqRr8gEAqybujZwPzIAGVYo43ZOwCv1fMEHCv7hG+PGe8Uk6bkQfse8/TE18Rl7N
O3Oou1NDQS58c9TAYDHCjB2Zc99KDlG0A8hv6IyUd2rq9dKc3Pnm0gqXukonqUBd
4tU3Gj8kuNtdBbH0VSkoP+gxg+8vOQZQHgtL8HKqMkxvATLeEhSCVfhK5APzQWaV
2Z2RmiBmpNPGW43zed+vp4L+MoSF4KpJB5me8tZAA8s2M+gd7PUUtF4v0FdfvToP
aSlXeOYyNUElYyrPm7/1xxWnIvXPJ5ATAPpFrJjzhbifnACHeHRoTF4cZQxrUdlT
rTKH09jaO5yg17XQ/kwEr669OdSuGHjVVNGDSHTNml9mNoFD1xmVrZEhwzlNqGTH
OHZ0Y6g5a1JYOK7RUCLJ1W8xr1dPNdGy994OhYrHVKVEIdyl4o+UKLbs5oAgX2yM
MX/uoTighGAgju3JTjQhUQqLZkRZa4AVDJQh36lSUKAOHlYnFzZadHp/apRFklDq
HUOQAiAV+HLV+4lo8R9C1x2kVZ3XAna7O3ssy769RIVJjyVvK45LdeXVKYSB/BgE
ngYwFlJ+gXl2yJySf7UhgfhJNxDLGOPaFkiFgOFaXUMylZyE+4HLa+V1wgQNrs3c
iHIVz7CDDrtgHxu5Qsv4vajfaD6NJTxAAv5kxgvpngdpFUZv58p/pYBToQo/mD1d
BilPZD9PYOrTzaCgg+2SZgHxTYNsMIPt0RV5SunCfTMTVgEPL3vC70XIrKsy5cqu
1fkspbWatw6G5THHQ1nqKNe41+EYr43dd4hXPv7Aql5u8g8mZCT2IVPa8Q2gVsPG
RSyjaJL7wR8gGmJjKoGy5mh1Iuz8t7rzXK8rOFCoej8R+TE4x0jbZrZDuxpS56mF
FVDeUtRYimfVAyOCvtcwMWk4YRH6n75g4Cu861iEbfy7JHT8LOJyqIz6ydK6jiOg
R2jlhe3qLZlo/4Y9ReuA2a7hXazyI6rPDhn/PctUw0FAkafuSvkIPjGhaTl1DdP0
pEf0r+4/J2t30g1ZMFLnTmEOcXI5mKPXE6cUNJAMN2h6fuZq/WbFMuDBCvX7pAlZ
Y9yELVyj1N96Lfp2zm4sTB2ZPQzf074f8Y4mXPG2IPgGPrjltu+U1USwoQVDA+0h
ROlZkiQqSZ/H8ukOBud+bnKfvsOMxbB/4FcGvDzwE4StHixMT2Kkq4ZttAo2IC2W
5LZM8XUObsCnvaZUds7BOmxxjFKN7h/lIvcDnyRJ/J5RlXIlN15wurpcNQpmra0a
krKhRZg5KEoRRzz2fUxP9qAkf8PLjB0RLW2v4MBN0UhrJMn3xaBwi0rxNFmL0cBy
VhGxUdcrXrbpBRo/sydAHZ79JOIrp08TryUVyCMo3HE+JXZckx5NxtM9R381Jhr1
p/JtHq8QBvG6rTGULaPogttkYYzPRFggm2rtjecKxa2YnrirYqVg+8Sr0lmqZUV0
zYbiEs0q68H/vPmjyYfALg+W6F88Quf5BX6ItuvwWtbWBb51Dw8Gqm1czEQB/rsX
hTsxQfoSVW0J+v/nTS/uZjUUKbm7bJSE7hDFZX0BMeKFNpk/uXuMv5aipzaKwgLN
XYEpRBeZRgsSyi06twQ6+D3WRJzMB9ZZ0ntTHN2ri9Yj3k/iQVGDSKmM7tc9FLE9
mLJ7dBvIrEa5WgguH2CnGWH5WckFO4ey1/ODwZLkE6/gVK2fmdOF3RFoZKIWo9PX
RgqgY0tBW0MJW6UhQzCMTrtix8t3Ymv9ngmtKCYa8x5jnPeLJ7ogDRMWpebQmSi+
fC6f38MxLveHocEtccyCllQddibCZFG34WnZHlq7KLaZVza//mG9wWs1IJcH80uJ
+XwPDP+4LOT2GKAu5rMKDym3RCUOyA0VOh+aExTkJC+1SE4VdfxrvOtkdWhuYm7m
F4w9spwD1JrMCdevnVZuqcvSgGEWHB+3dib5zAPJvvXGNa7V20Tmnbo6movLUImv
I2audPooMROZmjXoj/T8oA6x6M4KBoBqAABimOhh1Sp0Lm70OLwR3zf9xH04RrWH
klc7wfIS35ZhJckGDH2BsTQvfGUforvyd4jUsP24mfFZGvm4tI6A+PQZLyHD8bwz
ecq6W9myAjX9rQehvjhPNQEFHOg3NMpO6yBq6tUfuGSdkpqhezTxfmoyXe7qj84E
H3EQeTN57FB3z79ogD0ovNsJGLEXTOItJabRuPfjC40wKLJ8auA3C8JgfK8/ueuk
eLX9h09Zevm/hXADy2lbMbBhDWGBVg1yZUZxlvWt+zkmOBd1L1An3gAIKfY5Gwoc
J7/04+cxpfmfJPDiuzcP1tCdap6lsIErvNfmbeNHUdthCeae5O59drVQE0L17CCM
DTMC/umiWZCLDNRBls6IKeIF43ojukHBDbDKwe7RHjNlH/ExRHm7dNiFmga6XeaI
KyFSuLNfINsaksq9vu+Y1Q/2Bs4aB50BHj2ji2wEnMz8ElthSYwjBED7UhCU7xKs
ASpmeMiA2X7FDUGKTBeVXuBfhrjAVxTbWCgWFVldgjakWhS+l+gZYaMUtGD/b0jp
mKr1gCwKRY1h0eqQwWnQzY+6TI92Hzx4ODy+yPczo5l44CFig7Bc3l0Pyj3Kk0ZC
TUCaxEvb23Dj5oRNS8jiY85x8VM1JNTXIcQkh5mkJuNJ3bXpeTc31vZLkESpsOCO
02XjhLdpL3S9Nv0MfzLuNeec3LPCVkzfcqkkB4pCBSgUAqo0HWAtefb+yzqD+3PG
fnU4/sPASGNHmkWk8CGayxXOJRt7CQd1zmSMmyIoDfgSB32vOogNQLMTL0lKdX/8
HUwqREeOAleIdXdwjLwuXPo+lOQbYzjM6DWxm4BtKHKAGxqJ42NqIBJi0iPk6c1L
oFZR40jYC2K3NXovScDmpZQO65FKNytscTgaTi5fCzDXAhQZRX5Juiyz47+G5gMG
baZxwiIUophYVMvBeyP9NSE+lnxSsO6u89l6MekbV1p6iSAsnTqFa7365kZh/iTQ
DBjoqzuqTWnWEAuCUwc2OdtFgYo5DUk7OeunHZbI5xuYRn+ahOxUk+nmOZnAf4lh
U34a4fAz1auZV9lHCGSXyZ9oUxN2FmllpuERyqoif/cjczhD08Jnbj2/1cEMpgdW
X6RYpNWV0HCucL8HPmutqqwv8JEbvsVPqz9MS3xwBLqL3R0FucQAkMs9LJNeuFKi
K4goJc4/0LBt7gX1fxDSGzThDfRmwzF6OKZdHYxxeO/pAQ8NkdmzmT9WxXZbnHBi
9rgLXRqdLLyiDa+tIMfXDmosU0rqmmbMz+Qyzorpfkl9lISUaOMrLGIg/nKmgAMW
5uvgKdq89pvDj5h3vgRbvcE/fcynQvACeq9sjGwlw1Mop5/Y1VIow6N1JhougM32
7BHh0o4sf7Irc3X06SDDA8LuKpsyl4wYInIb8+UToJ2QESYQeIzv3UI3r++8S8Ur
WNI8la3po+LWu7+eL5nk59q4ajq2nvRPV91r4ONVOyV9NXvE4saJ8ygI5UPc1wVJ
qP95qStG91ftMwvFaEW6D7LUGyirHZdnBWYkY7f2j93NwbAD/xb1hjVklX5MQ/l1
P8MCl+XIfyG/PXc8fT9DPU4PL0UlIQ2W+NLz17dTUAfGDmiLbgzXZJksWhRAS8gh
pOMMSmqBRe+zy514F4vg5WW33tLPrbc+CD2cfJXvVyvPjyH+W3unC4oB5yOz0XBS
gKzPdwJxb4dMITXxq6Mnf6MLKVxOD9WYZQxk69hC+tEu+vr8uTgs7IgJTDeeGpId
zB6a60jISPwb/4J7ysgkqdd5abRDBF/jup04u78SYg2AMbWxoWL5x9rJUyXQ6RPO
DbKeJoaxybFGW9zRXuSstWCnXheDn2grfS+8bc7mqi5L40Sc7cuz9ACBKp+cGacX
F80k5Ml257yFk20UPEz4rfe2bvUxeie1AAziX7UB6JT+N5Q26IY+bnIevxeXumnl
1S+u+lyEjjEA5c2tbzQXQeYsuO1qdbVibPGPrgTjEMeXrlGrXaXyXAKxFPYI3bJ0
W8M7ubSIuPEpkfvAhdq5le6iZGUGF2wWuuS1j3uEfFnlYItYbl50ZRD8YR9HUNkl
uTu+IBLTeP7dvBfLUnaLjeQd3CV9uqpQD+q0w2GfyWt+w/EV3XcZVm3g3A5NnfuQ
Bj+wzTKvOVM9E/5v0EaGnkSTq6qOCjzteBKUlV72eBsmsT/flwu50Nen7s2cYC5X
LkHMSnkWBFQ6ziptW5yEK9XSbOCndtxhyYF9XPj7v4qqBwe+Jv+2noeoc0tGAhEG
Gajn8Ex/z/04TiVlX1c6D7ofhaR/DjSDMcxutJzwzQY0O4S5PAjFngXbhwM8fLOp
nRwPF+RhwnVe6s5CIaS7keeYu5V+TWEFbJLXrI57nfT2qlsUevMAudzysG1dA/qJ
d2w86k0tPJ0PbaO4m7TltbmXqM0MbzYvHiLW29a1zGbDERGFOmoZOXaJ3SP05GDR
z7f+4ZbU02XH/up5VMlogpaNVfHKUJknP9oYoJizNld0bVuAo71604Tyez7D7HYC
7j3dQBgqbOPX7cH5JyfhPivjecy/DDa9/XrDP2uXTOlBQJEYrNvUI9uJoNay2aUb
5NU5XTIGbRUoxoyaB+O14ikOBk+bW9i+FkC4jihHmwzA9ShqyM5SHtQB0BFJMln0
4GNCwwqIAJ/N+iNwAP8//jQj9n/s8OWF+BHeEozs9LN/qtCR3K7QQCjsGr4aRZcb
Zq8PcuzLpJzSo9QX8PO0JS5jRzdMTjh4shdJWkVrMJamXAY08MjiJiAzlFgY6fRY
7v1HaCK4/Sd78CHjVFeqIOKbjuWN1F41OQte/IkQ21EJsMGF/HBq7pBqaWoMo+DD
sOmkrZcHvdLCMcI4M70J5h8eOjAoD6NxoYt7CQlYm+orsWCSb1ce4ypOEGq2mnnN
oaaDqnkM+gsGMV6MnWwqADBA+1xsGknjfU38mnxmQWHn2GCtc50/E/4e58V+QTdv
fK6tk4CuX5t2aUWbceBwSP6eEeK+DoyCbFs3Bgm2IxnTbUkAIGJPVnnUqODqtELE
/7cDiWRJCnzz7TUfXfR6WZk5/KDk++tTppcWxqvx0noi4ciVgNkT25GgG4sJhm7R
RcATThG/j1eu9cH1NgHQIG0pCBxJEO3h3hO4SmnVvTnVzr/OImrapLi+36uNI5rG
AjMdMXBYNTwiReN3+pRhn1PAMJeFLlH/kbnbIcXrTtCbpIkReCx31CBrF3VS3GO4
6wi9V5vW6hXIT26j/zfBS3P5pftdGZogLn8/T1cA71OFjDCQAxgxVfcwJ4vC78kv
GJeSvswg8GvMskV7Vf67pHvE4MT2ZOHr4ryGmaayHxX5E9DxkIOz+JtoQa1k28xE
d1POlbKV9sEiovazkCHBOnGHON9ihrlFRtFAXHor2+Yps6+950S28EYWGA2RlpX4
nOm30BOaC7tWRLhzRwYCGdrvcxzdvcizvzqnAcNjuvrZSLokq4VkTnvrfbaeC7zf
2Orfx+/DCX31hAKLwdhhRQ/ozGQNSLe2IG+nm/12ZE4F9zUQ1F8MXTZ/HIMMdwOt
lAMTcOVQ5zDrs0MK4ajaaaoWvzVB3OS2jc9BpPdjek1Fzc/nSoVQ2+VJAJdfsLDA
DeqIxW8PEX2xXinbJvhO0lWjkNnwOiQMDKMKqRP1EosYJtDxfQG5d2mzwg6Ie0Z8
kVub5f0b+SaFM0hWRnerxKQV/c/CUVGRQdiPBXXV+8SpyPyQQD/fLrSr+NJGObzD
rljUkhQJYgjY8UwLdRn39PI9YOesqY2YeZjsGSqjJq4O5UlFt5umLiSTSI0OVeeG
lXfcnY/m903op7K5Mtu/01qcdzjD8/Cp78WGsyhni96aw8b5Gy7jKyz3VKNEETro
kwFAvhF0Ki6UIGSrR/3f2Hww+nvbS9EsMZSSF/6cOsO7D4nR+1xzz2b52bjG4oLp
XvRyFhSGFpiWDO43cPnkdzeWOyOVe9+BCb3rE40k7UTD5Ax4QCHvWymlKsASeqSK
gBV1qwSLtIZ4MLwWd2YGCmk2v/occKoO3Kdju67v+Waw6g6gD6l2b/Q06x1FnLYE
uXtRrClzyrslt+NZzdwhovlSu7C5QxgylglxOgmse9XJE1Foc7U+ny4x4VxNQIm5
G/yEzHnYOTqpjjS54E63yA9Nx9jj/lbrM3nmePxn2LXHAdMM2xctpJECcKh7kOw9
OnHc/WlEp5KIt3tgFjoVOxyUH+NXDD9z74EtUlqlYg1ptv/66FPE1ONQBoT12L3/
xqV/nvhX76PHtQOQ/mX8hiOby8Z1at6rVeTKgsuwAUkVErSUEV0MC6+2vUky8oM8
3Rhi4VWiBoqQKO1w3ODRr/fTPxtXAmqy5EMVj9gvphjMPusWNBFDClQ69j1rqKJy
CVNdWkTLgZjIcDbb1KRnSkLo6Siw51H6s88YMUCkUh/yfjWSgzG4i75jVkmYH9sW
37p5xlW1hACM04BTNuDzSxUi6vVq7sm1yVb9LY7jTNuDIjuAPeO3IH5Q//UQmx5/
QNC6HCrSPyfI1gE+/a/YFTZA0eRt4r5IpGMeqFzxaPJmjyo6D2dE3T1p/jnt+cH4
G/7wsS9ZoK/9AILuP6C5++zuGh8uR3YRyjxTXTuStKSY/GpnAwEvBxM2NVgxbcCD
ejUaWneUoW8zT4YmU5P6YAQZdkFpt1/Djc9yOTUy50bLr96gANj8E2F883Aog5QK
GFX47GIhqejeHbd6J4Y8T/+IdhpJJ0+SzCvXC2dAtENNl2d7VUAqUmLgqW9XYCVr
/qi9MeKpM10hvT4NzDWkMxAGv9Gqwsh3PwNjv3MJRfi3HdGTSUBkXmmRNCOHzoec
ebV1f+whUHgO5Nn/w4WKIyQsTXtzPyXpJREQF9f5NII4n2+6GzXqM6ua8CTTtbjh
ArsLv1xKcWXAfjEpMUFgG6I8IjhSt3Bqi0GZLYR1mszU3VqhmNNytF8PEpr6sNNq
YjcyCkeBe5IbzD1xGgCTyjO7bgpLHO7weDbm7krVBhCZftb8+fITTp/rnc0VuqSQ
yBXm0XbKHANFzZNPJ+IwgHG2PlfiYwB0umXpYkqDeeNKENGkf5fe4DE46BY0dOqd
jNfaqRwqGyx0bLvk0duao+tssRh3oP8dBmR70DA0QWqGyr0Mn1VYwS9WzVM6+gru
k48HO968YfTVlSHgjgc60cwWjnrmVrFo8MiJ57GCgq4s1PmJiejsT2IZI00Y4Gtg
ga0UreKiH1t5I19zwfVDWsRQc32T26setiGf4O2CNF/oAd+g4CRdwukDRkxaYzLy
+BihD/QcXBptoWsZv8ji86MWV1DHHZ7yzKWh19/Y54A/15pf0yGuBc4jZYaAhlfW
8VdVs3TrqTrutwir5TjQRUGpiebAE5ubiT+rLRJqp0cTLBiFjCYzJ/+wqTQnToJs
A+/5tHTiW7VgQ+XIMtrZgLb34+0aXx908E8TTRwwGZVpYv4rvQvpWVZq/AjZgJE/
ZfJCNt08nfK8qqntpMfeoaz/gGeqe5//jIfCxjWyzNHS4/X30xRPfRiUroUD7Ki4
qBIbRM6ywpWjVb1iaE3isyxBCxyMDCtLmFcDYRRaQIsUtc7gYKzJalztWLTMfKbj
ILLZURMnxcRK+HPO5n67qad1G8hf7yPyRlKNGGxi6IyigzOW0ikVyFWsZfXxXsDE
18y+UIUrlV85eYe3BnAdiHq66qCK/Jl1yd+rIVceuDmu9X+jnQIhTyh3wz7UZuHp
pnYIHGjnRwggOc1JqdDjWvGBYIBDnFi8TOA3XH3ajOv6gt0S3xAA7t97ahH5udZ9
ij3dLDUYmLnUGBml3C9Mzhci1hAHIxxIvxH+L0eyMBSJ8yImY+C6C2kjy4n1oonq
iC23BREkd9tWWSF72qDtjdpesJ7oL8RHM6g/TRoijF3S9HJg6fAH+WkLZfz1L9Fo
21SHtnDtNvyfJzh0QlZUrF9D95F4ak6INot74y6g50RuaUYhs0AmXHnf3TvaIq6v
0VobFPPkNHZDAmL+XdF0aanO24fYyjQzXO+sBG0LuhLsVTY2ZsEhK9DksyyNj5l7
enFHdtrz+Q46Gy/4PkUzOM8fJRiwOCEGLi6nD6dINL9bHNneVYc7xPsjsennBVfI
FMMK/LFrOdI1S0Y85e+NQF1t8aBX1Zd8ZCb3L4IQOC018nME4iZzRe+EsmbuIaY9
LPZCNeE6GTL0P34f8ucr1sK3TnLsj1tlPqTAMNyoxeEJY4iGQjJ4WT6zNuXNebBh
Ihmx44v6byXNEtEgn1jsJTaJD7zpeK2VAUzl+iJeRhFYNZ9DeSfOstdrIf8AT5LQ
F2c7waLYyczrnBF0TVxF7CQp/h1Cf2p4zFYQQcd25f9T8Etc9Id1U/w3TlIvuzbG
PSKjJdUdGbnIT8N4poXT4jcyiGKQ5qX7AKr01cs1X6oc7/b58Fto7pZk7JfSf9Hw
psTOo9/kju0RYiOnuCYpuMIMyJjuA6HSLpYDiYMtu0Db0pbcTIxhjQZ3kS5RnmUA
aJxqkIyPXD3/NtJQqOkpX3cBk9+LKLNnhlylUaXMnHYIfIM/mH8HY8FvavIcgIhp
IgyUcvOIjh1VvqHuJEKhzQLPVIsBrs+H2bVsb/ZU6WNS7fODHivGUkcjJS6tuMhw
3SxDHfsQnfsDsxo2T3R+vR+Ls4EOKvan2x2HO08+1SEW2QreiDijcNZKWR5u6AhL
suIQMo2ZNVY9pa4Doiurlt+a0GHZ3OQwErnBAp9igQw3xW9PUc5Gm85apLY3gXUt
kHIlVNOjbN62TJYF9kmvDCJJ32dmoozsvbxN3L+ErGA9bVZTzmrt8sAU9gQt7vs+
xCZCloSV46j4yUgRpLlagK1ts+JmbAzMSe5DG5lQCQgoORVwIwUobGlJyFgpK5C6
1ob3jITpZI7rKRvyZqKjOyyLN5GqxlCD9hpkzmAqkal49rv/PZaVdqj07YxmLH97
ukYILBXPCwMDnVruyWRabsF6UIXWv+Q7DljPAfpFdnAp4O+ela2+0kQpUUHiy/X8
blUQKQyq/vRvSMJToxRFANuXlRsRlW7Du+YcgOFbVSIHP1jtkCe6To9gJ71j71XF
ODCzGf/JJCZ5LOU5lm0gcGUInHOCDQ4zUB5lExxePgAfeJa5o+DwYqf/qF3ok3SO
iTLccTriAsX5VLt+sTEKaClyfADlzBvlgSBtP7EH9/M+gJzbJvglyKVFhVgy2QqK
euFfK8H2FITr5NDa/6/Av1ZC0KbVMMWugAWQrsqJIolUeaWXpjZdG/Q2GT3Uxryt
R05D6i5sjvGJxxZvNIu9DZhOxl9FjCcJIZHbZ7C0FVrv70Myzwz7fnU6yf64mity
e97wTbj938EFU1rnUaU6vuPip4Dueh+adgjfj4aZ55VFIONhLXURn8Y+4oAWWmcM
YNKB1wckCUcUBXEEni3FW1w1YmRK2oEPgp8Ay025Th6fUFxPFw/om/mceJ3Kqffk
T5pa5L95DjkphF25/NxbW6O3/5+SgFVKubbJDEyrr0fiNKpRupBi1T3ztR56scCX
oB746YwJxEWhfQBSff7VH5Hw+fRej+oULgjWscC0j/NpQsnD5StlH4kuIdJ0M+gv
RsCrrge06JIjkpFwoOt+mPqTvBdvynZ2P1FdGap9bLmOqntEWh9KLp0m3W0JCYYV
6dP8YaE796+rER/m/A219O+NjF+EkwaYGm63rnt5z0K/t1hQjdHgNEENec+bA4rJ
SLPwiz/HFjqQapZtYsZZYZEX3DOVpMgdhBjxjUsc5EyPY/6lgrIEHVt+BE0u8qp/
+w+o+roWYyt3j6tNFZSGxf+26rIBBNGfy4T7QPYCnZ0I3mkgshRD2KVIv9KukEXV
smN+tyi91ZJdzSPW8EDUKjkOyqE8xZYeDNTqdY3/DyFuopHdVHD9M3cIEzOPEMNP
Wrc02N7UHKkxJgAhLkIAv6bmm6CwZxk2+mVvLz/9I8jkB61C2RW2CragfL9mqP+t
cjvZ63Q5bcL8V7s9vquMogOhcdXy9xWN0G+su0z/G9/jO1X2Xm9xLGR00XTQqzKF
2iAEyMN+FyiGfqHbIwiN3OLSqeRbxrsKKzcol0qIENa2fnF62pdxaq9wGq2Gbh6+
JhK//l4irEeqO+E85gK9ZD9BSaYe5cnP356a8MaJOPuc9uMY1LbkAl7vxbIJteQV
zJhmhKDpkJAvjg4V5jW9uPMsv5Hd2kvzhpqMas3x5/LKQfIGxIYDTrnT6DIk/3Tl
01wuKcR/mnaP16xeZLgpNwr40esly3RsUCFPQKlPHBFibyJ+N4rAddAAV+thiiSb
QQsifmEW1NqtH6wtM3NDUAmG82Yi1PQEj+z00CdnY+9FUKHaNnWcWNf3yLM6ynq/
e6JwBs0/igANjngnHGhYFppVWwIrQZvgCAUGe7KdHJtej18ZUE0OdeXU+Z4s8gTd
VPMrmd4RdKoP5TkNHFhXvFl4h7OdiAtLq6eN2+k589FQ+fG6Z/XnHiY1GOiscD+L
1hYr5pCAEM/wrEZ7+VMZyl1gtWYHNPv+Fn8JbjBywyvyDSGe3zwxAXl7RXBnA5Hn
abs9Q0SwLzYfKNvcTdIsiOuSwsk/90uATA7niLunOicbW4i5YSBWxOuGE4UHXciY
+qYisoyewIrwtkXu4zAIkO6crTXoPhKt10qGu08CYoL5/SzO1YFglXPnf1c6Nhca
GZMB40JVzTu/FIzYJKfhqyDEGlCsHbJUMcCql9UcvwiQbI+T5aB17kMQ9loUfS1l
JP7K4DJaNKi7c6k5k3vhr1bgzsbt3XSSmeziQ4yWPwGp3IEx2kR2IzcCJIQLCjm+
iex51PlzbH/IGB0cxzWc+hVQyz4XMBUbqJRCVoXR6rzd2R3JqXMsB4D6Qk6+S7D+
V4+Lkea80DU7Oug4nmNVpg6Vrd4ShRRcM6Mxok63IJMNNO3e76TbbsNbG6sqR8J9
eP/pTaA6Dz1Q3noz2K34ZZIh6w4oPZNpzm4NKMyHEadQ6ODQsfNXfNAywMcQCZON
yUzkRxiE0vskoZa0lBrvgSgx0odkqKH81GVnFKiAE+BJtmmXH5zxf0xNL5tjdr8n
2djz01glR5WX6qko0NFZXNAoRnKMPOHc/TNn2CuyJmvfv3FdbA6o76tnnJ7k4xVl
SgVVNqXNOWsXQ8JwGfJH127HIccriXMvTGADoGbqJBGPBbDgUaSfbVJMTbzc/Wur
R/j4YIZm7ChnfUrXh7EKOXCKQEekwvmfa+ipELtLoT8wnjAkLiosmoSQ7Lm52yvB
+npQJg98HMgam5ece5P0zz75x0OzEFyk1ZOeAJ/Ouk3XbpuBQn3ZHIlxJt9x14Rp
S0GP4re9VCqO8ZQhesqKm7hwcAWvZWBgSiGyvf51FTEMwyWGP2X4JND446r6KOiu
G967jbaV1NHwz8Y2TDnvNQMmNfu1y8iEZ/FPPzgR2PcO4JzsRQvBQUC1AK9SsJvc
+CxR2bQSeXxBxyJL5Vmc4+08TxtwYzllYPziwrlH79igkp2hdekmiqo82da/rNck
lEy2W+aB7RmU2w9QZfk30HbR50CHBL7l4e0HF/qnDCiniLT9OqYiawOFPjiDiMJ+
ORnoYjD8TKDEMAkwIWmFnVt9xrplvdaJ4+SaUm4rI1BFsxTN76qk+pTjIdg6F0Je
Fb3DSF6B0yb51mxpx3MPNpMNpxo/qW+EGEBRBKBZ4EciFIVRUmLz/LoAke8yNeHQ
Pe/B4bN5Qm3gF+XNO68hlD6SSYvTgpAXIHUrKSEdounnExTeDQyV/ciimrUQQB/S
Pw935zViWxbuahpNLpLDuw5HP2b1NwYO6QKj6NtzF3DxB79MqGlQqzERK46YNKB+
BWCnOB01wGTwVsifCu2K6goanMtp5/s4zRkoP3Nyga6AkcY4JdoRzW4s0cmjZkz5
R6V6DxiwDrEVJePSiyfJCwUutcXV8QYFF62NzaPk0SAMGJwOJwEjDBydmBXAURcb
x2uc3DQx8ewZcvgiZJ3yzrfnSeKA+os4YzpCGua1Sv0EyTNgI3Q3Yr2eGmI5ZHZV
Tdq5VbYU6wbNMKmlD+2CLyUQXoobvJzeuv92GMpLm3+BdLgsUCfiHbwkiS88B0vF
JqSLYHP/lf4zdtI8a2qvDB7BW/hw+SiCXFWxG2+GYzRwHK7BMgHAZAkfo3hxaqIN
FLo4CLa3HnE+jP3vxrEWqAcKy55tK5kNDmZCP/XyZbcaMLovgctQiNLTckWUWzwv
C2HI97sZWsA6r0lbES2ZrdmZ2NbrZy9w4apa5cczZiaHeaeItdgD1quU4cFeaBXu
BxJ8Td32TYHgmZF8Gn2jk2fZzDkF98A0Kp3BxecO1idurTWJw8f2vQ18d2GREGHX
O0XDKStcCf1L6hyUjIASd7dh1CMxjWdtBOIRamQ361lhOdHpeZnZ95icEuVAbMAP
1AA0W892+5aylhy6DENkiT2IG/BCmxjrRkLN8gqKZf9tJtMK4RAQoO2ldxR3Gp+i
77TKvWq8GoEV2qySPtNi4V1yfZtJ3zya0IsyeriMFSLCM0wHWSMS2+FsPton5Q59
lQA8tmnV53e7xwb4T9P4Tf5hTipLLHCrVw4xHHjemoC37PC6Yue8ZXrJik4pzkJy
/vx8jFFpMpNU0OUJAIPRV039KpXSLWDGJZky69R2IqkBtMnsYTl3qFijvc81WA+Z
zz/SUUsOQjsyJsHk3EZzV37VQBhYPPrM35rQoxPhVF7CxzlyzFZb3/htStckmSki
tToEUWSdGr5CfHYRI7NbYFuBXiZ/B0vZlEHu73cruWPbXA8bazIKwzwpUJns+Tum
jQInLLsicfYsbS+eV5sIasUkSNVu4Xt4YbjF435SKRuGo56QactxAIBU4MP4uWmc
Qiwg9q8n22TuA4y4MmG/u8qlXqLIixwxYgGJiI/KidccVQKb/sxGMJEWRMIcl/Ah
RXjijcAxWfP5KY2n+XA/S55uuazfbB5N0ojyT/BnebcEVwm6KzmW100GkRWdaSGC
7vBXTGoZGWsbq7V4bvysDP3wwYe5CZw2+7tMhKeglbrBELu6bd0u110QzchLFYaN
pUksDOf07UxJZ1VmSBAdNS/7VDpI9RLgaAP9+sbICjIUjGcYkIicqis06zJDzS4B
jXNTd7VtLTy2QgyFXqkTPtaId+PzuuZofxzZQ5EkX+dbPGO0fAep214uawtXcHT2
OpWuMGd/h+IaX2Z3ohzqPeO027uCR34evtRt94Ic9VpXCF57nE5+IkB54T4Xpbm8
PxGPUbClzWYkR6YSVNY9DXu/jLQyUAnZgzAuLBY0O0LuWVULnolx2jgbDTfx1Pvn
e19c6pqKIFeVxBDK7TUrI7gGZFrvtRonVFh3EwQ2kvK4wrRB6vYW3GxrEr0ubeT9
9O7fZznE7OGtxQVd66MyVs+MIMOZ2e5pAPjrEkbuuxLJklUaMW1uvErUyTQkZjmx
+YNna34Cd0x8vDkV02JuEMP3ra4kh+DorNudIYydZ95cRA6PCTNaFQQrPOMILtMv
kdu1Z0f5UzZRVViBty4p7GqWtaOD5goH6ybXybgw6Yskf33gRlOEXzJgPHH5eVZa
v8en2+v2LSPYFSw92Y6qf1voVAsIyjjnDA5QPUd83zNau4VBbEwbWacxAQE/3lf/
DC4SSY7m6vux8kIPqU86AncccMCYbbwX0YuRsEkWFdEH4nzljMeo/GAH0m4bhjAJ
AqIFWz9zWwc60xAJhgp51cRo/WJ/MNbzrx9hIEke3QJQFwyBTYo3PumTLmIKOaET
Xs3kjhPRqboWfTJ0wS9gchKBKEHmMaxA4ms2jVKKXAM7Q4zGBQS2eBXjr2B0G25Y
tC5t97y9h0iARbpIYj9Xvf5gC/9T2hZu+qhW+dR6UUMPPDX9/yIi70l8I1NiatpL
5rorbXmKnDiYGm5X9Mhv+MBSbv/xht0JRb3BS4WgP81uSSz9Ge2DKc74DDzSSuYC
HFULGExhJ7Do7HQ+PDRd0D9XLRejlIoz2Qrhd+LRbyAvopj2L2gRPtd9cskw8xQu
SW+OaLNJcId1XU2yvEQJU0MCn3zV72jXYMF6ST0KQB/hVm0JfWMm7vs9u8EB18JP
qCfy5lZQrO94Q1nmVK16ER7QMr+xyJqvYYgkQ0feesv43UlUgPmCi4UwwhvRtAIR
XLkEBP0ACSb1i7gFj0OTJCvLtvLzvoPMWZCWh4J3d/JAgKP+7HjwR+pK1Oz+TjrH
4f9Dqqk7EWna+mj6r4U6xoWfxHpkVCRHkRAUkFWD/eoVn5m2gwNN5rAyLsniUg5n
c3ogsrZFapeIFoDwMPiIQyKesOYAvHj0ou8uWrJphfkC3ZFN0lp6nzWOWu2KYqv2
kmpea1wHohRDWWUONmxuIh7NX2Iz0vOT92VyeeULt4G75OzpWVmUuALTj14zwHiV
NuI3xpu58XCXsLFWsr/reRz9hH+JdHEo+U82gS3uiqhpA4lfP7r04YXYBztqlxYM
QcvtIvLJ4ae0E36I56VbCYb+G6ee97l6hRZS3R02UVL+rBP32wMcHDeF4W6FrVrn
vhB+LCMjFUVyGmr54rMXp2/bs+tehcDq+k/9xhdat1fMftW9jooJhwgJQJl43YKE
4wBRoFVd3fM0D5qmPUJT/aibQHQuKDVx6+Y7FCeoY0y1S2GhvsPxeugUs7vrwCto
I9PxdoYvnCkK/0GQB8iYDIsFuIiAqHc0kKyEOm+dfzMW6rZdRfMM6aZ4nlJbppex
SuepzrhX1zahlqjeuhw2Qtq2euOaiMidWFHRlLR/UWWgIhskN1aFQRlef5DnnhaX
Xo18b3s4OZgxwpz0T8AUeLP7p4kUkeR/SOFGxVHvTUFaQZW+mSq0TaGlfPxaRtHN
5drwNNhKR1EEoz1Gz2PVLZ9Lz5ESO9c6ylNEzKlxnBPx+cNt6u+7OtLOdjZ1gwVC
5YGoFxy0IK33ltPC+rH9mnLLxZIixRab++pOo5JTsvFxg8ED5zqxRd434R8GJfa+
oC6Pq2M78XDV0jVIrS+jKdUX/OI9jF2D/mnByNbLDAdMW0+uCzmANRCO2xj+wUAN
UpIaz3O3TSRbsL0mgmxgPLmjy5dwoumVodcQ4zQXmuzBPY8usjcdwI6mE5yuhUiH
b+II/wuweeWTuGbEOepajRbKsCnBMYR516c1mk4MS1QEWIYPT5Tyf8nTStjTAnHA
P+MZDAOklT75obTBO7WmrNPcvVrvlAcQM6nP9L0TAw72+CX9IsdWyDZ27YUA2qJ7
IkudsOL6ojeUshgHjYnT/PUVMK4i6kZv6IZ01BxK3aJQBsHFXGFeFBTUAmMzg7aF
1mmgXxjIA0hJ+tFUQlSUNrYRtJ7kbIYTNwgwkA2EvBWf4C14n8KorA9+1yUSPlty
+kBKvLHuYchl3g0yFRretVvDLckUiiMkXZjA+oO11P51AtdOnmIfMRlDAm9yO6Kv
Amq0IwMcMn5WxV5YKOKdda1TlGDSRFgD/DS3ZZYRVpviO9T0eJ3FbB0/07uNcn/W
aoveaLUe8QtZ6V+9OsiD6P78MyZUTP0wmEVAzlA6MLVP3vBOV36vrkgU3ZQoUFcb
B0xIXMJR8p74KBT+d+xWUx/OmxMxaQiruXUUR3LEKFPT8BZrBHZnXoXF814zNuSc
dIYdJ6cgTm+nd7mkNeYMidMP6fmsxm6J4sbkJBLaCc7yfQr9HySsNBP0AX4dWBoD
3DghTZnYlI+8aa013WvZG9p50z5Bw9DDLGLkfX9TUu2u6E4ikSkdHrWCdy45fD62
Ufir8tys8jPK5+uQkdOvUbVVox/wzSeqZjA2FUXosSEZojj3KWG/5ros0o3hxZKu
P3uZD8lSMeNA4/aY6W1QbMIv8V4ZrwEChrJ46BiOGADSRwRMi/B38VUvNSrVEoPO
6GhYVInmKFOu36KKeguybz4B37MfxsySxFrZNAm0cearpoGs+sn3bl4uvwixV/ua
WWJUA50s2Z4NrkBwoY7SVsZQpeQK6mjEBM2T+gFjkAnO7D4nnV7DrmvTf+P9sXEt
RKkrvqECYHki1/+pNEIKMbu9bqC1d+tKTKEfiZrakysY94erk5XdoYZ5UelXdRVC
PNpZNLuRetjolEwOiyG8+unbmVC31GwsmCgEx5xC9V01kJvQSPAeMpngLc36pJj5
aFRY7SP6WsnsFanAV/fe5GU9rRBhrHOa0YsdmBpCQ5S3bQyuBxOQU+PdM/RvF6eS
SVuQe3zzXGFIgrHdjw8erQ93VUT7NX7jbQ9ev+rsJIyUTiBD3O5WIZ3zC4r42hqF
IfKnweAo3GmqffPLNIsQzwdRm46DRTznf3c7MGnJYSqU9W0ka0OfhCKTZhl3kpw7
9Z53vH7Ajdz02IJpF2fPDisQQWrJ2bQewtj+SRBCXGKfT/sNNTyhGaaCm+abqznu
qy2EkCXfQrmwPUuCaXw21bIVqHkaX4ANIUezSZt3jw7Owd3SoG/UpZ1NYg5qe722
f4cSsvpztl4KHQ7s/MzW80rMfsCVC7OyalxMHpgPhhhAjI/UmWbKUnAzgI1XFFfr
7SohnpbXPnMm49p4YkArCilq49fwj2LRIbzv8mutufyC172UDr1K25SP1gKSKdXj
CILlFgukMICoBQRTqEWPqapspOAAQFq+cU7dc7ROqrxTLjgtEF4aORAKWzkgox3F
y6NNNQ4QtvpsFKvm6lYwPn7cfCzkGngdn7agxlRy7N89192VGUTlMVTowNrb/b4z
UVnXQtuRjNSg6KIzKP5pTxZHyMd9K3JSYo1aXlH+Xds5RFMIYZYkprF4iWw5EVQ/
lhSR3U6DV5oz43RwgvnPv+WwGOe0FCUy9rxYrP8DMIASOgdoBBiIHsN+GDYvqwg4
RGIJ4r8L0pYby5YTGtBNFl3pxKlrMosAAL2kw6b0ZOmW3y3NIcpbyOVc+c421m6I
pckplDXhGZsA6g0J1xABHQyHAqQNRVcBKD2Mp6qXZZ6WdJn91mX4PPuc+GRH2hiG
2qb9tBdlWPg/9nVr6AbjKa99gf+HlGMWdwdwl373chNrt0lsxR64lkJx9cZ438g+
U4fMJcdSEqwphrm6Zclt0Qnhe37977FHtOnXlMOwLfO7BvtMuvAWNbWkP7FkZDYE
pVgmEeETlUpYMz0gflK5HxQNFzf+nPKI9exb508cDAOx5uBk+8KtVp3ffOI/0VmK
edE9pl37u9Uq0hXfWTUXXU2RSZjT1/bPfVq/2E0Ox9U5OajovKJQIox2rLHD3bvI
AGbQiZjJ/Sv9wUhrQLlTYMAsynp1EzjjRO4grfOLQEwWJEXopYzUb5KbF9YTMqnt
SbNtfFLk5Q8N2O4AlcIwLVMtAqj8fQZF49TrQtnokhis9D2CCfz9uftbvi+8Gs/L
GiaRRddXR+ZY7dmzpIObDJESnpKBr/Lbkyr98vUnBfSenxPusNYiSU023oZ9Yi9g
KU7RGENUMJ/e4kH5ScENDgBQ9y722SdHoHQ8nUWZmt8rrQxc9ugtkqFKgZKDbWiz
XGNgm2iQ490rM8G1OY7wUdGTKlTieuzpU0iycJw53KEq/1QjjsAjVcW/r6TCYCLI
ap9W8GzoX1fZvHDbpvq0TQo3q72fI/pjBgCIssXmkAaUgrtXQNNcruqAbIyJ+Tc8
Y63wUYztYBg0h7E3KLYBnuRW9jJARxbKErxrdrlJhF5VUxIrylNIU3ycIdGmiMLp
Dw6gyIG8jmiDdFbHIpDDtK+XmdGBKemuww94ZQwrQkFiHbtTiw08946XM8Sp42nv
NR8i4X1lbQXowMrij6WMfq2B8sgNbir/DZXl+r1oPpAhQqglDwrFbuoR6M5DfCjv
za8MxLNU8O653RaM9/KzVb9Ck6SBsAF7koAtXqdI6y7MHTlzb1f4zM2XGQ/mvUK/
iovcTr3efBR9AjSkmDbJNQOlSq7sqUro0CaLHI6w6pLhsMLnASY5unG+7Y0t42Sy
exr+feRy+dS4LJ6KQr2Sq9wNYkdMu9QhScqIJHEDkPnT66PKcg5VpRPMWis3J3Ei
Xjdvhe46nDN77Fdt+S/xMWG/R9WLRogtVzUF1qp0zyd8jzc4Xbv1/huGAyAjFpem
SBQNuUP6gKE5GWxOTVYJdq/CslXjW2+M7u5NjUzVKhO9tNZKrwrrK2gAsNW1z2hE
WkCRB9BKgDRciiiNORSUE6JyDyXR7FmRQK9a19yaf5hH1SRk3XE3uBE6acGR5Iii
T9AgMjzmPWDOkNa0Uc33fyEiRhH9qWUIIYQAWdBiXJYbmYHe1sdRWqnE8j5zCo42
3mF6e6om7NqZ+7T0lGcgFmdwQrFUqqSsLJ5+56gTEIZ9TgX6QY/XQGCaby5dwBqt
HFMgrcMOC310Ff1wj8q+lpsP+GtHTgg4yFClnwpeCNlufhvO7/yPzhakpbAtMgKy
W7ao532+5twtp7+n4swkqGXH1wl2vUlKvevdM9pkfhNzpp5SaYenCMDJWyIzT9iJ
ak8lr1HH7CtDadea0DR8sfX6Uh5rr+Znd5byyY5uB20UASmkcOwUWFAMCA4flbO/
qWK+HS92T/GCa0wvMQ9olFfxRukay4MATWB95dyJaKCM1m+Vn6wzaWXfnEsVRKa5
eewiAxAfEbRxdL1vIP15pE2BvjZfmOC3sFNITp03ZUrKEYY/ZxOg0mg62O/0NCOL
yrcBSKEDVwf03vFvyskuOWiA12qath0QdWoggm9vQq0HJ/5EHvdfPBkwFv9O1bmD
VhWxuTM0RsUlhoBHq3lBB8H69sARrK7edeXrGNTrfZkS27xetPhR/NBSf34iqA0R
YRYqsZagJEGdiSSy7iCm2Pz/7rTOnnTe3Ip/fASb4udF0iO4fwQNtVzPEKsjo4qS
Pjuh78RvULSoQXN6z9h0uaceZEt07jTUBVGE1r4MlKFzD+ffIrEh6nA+t42AauNg
v8Re4a7Pif5bQrHZJunpCGICbPf+Avk+OsSEcKr7qV2Cg08/xAIpr+F6n3O8ltYT
BdUtOBrImejHUaFtJjqTP0zVBPFZE43/dolB4crguUi7hugxMtEk/Qxp/Dm748yU
fRVUmpX0nfAEh6FWwM5pEzHgjjlJEiiZZ2Oo9mbp3RkeWJJ6tSypu5GG+k68XdQ2
mWUTo3sXwdsblcosMaf6fiQBVIJUI2icDJrrikdFHtus61afRt5d5cFOrwzA0afm
V6vByeTehMZnld4Ut00hIfNnN3yXw5pjmkoAmslHyMxTU5bL3LN927cxvukiAT9H
qhDGSXNMmdDGhlXSrGTmP63WRw61pmlGSVhJfs+zz7heojQXBHll+yJk2UnnjZ3f
MGNcHRnzlJvQ/ap+DLbRi+hkg3v/65PLr7ZA519C34iMZ77UcK0ZgCoaGSY+c7fO
WdL/MkOxZExZHiAGH4HrD36jxp0csPxDYKWB2At+Iwz6wlMORyeoT/PRH5HSibY0
FoS6Uit2OyJxcUXNL7qh2BZExvbRajcK/MhzuC39KNumWyI7lenrXsOCH4NfidMR
tbrebxh+DAcHSBiyHpLUXDwA9U49xuOwj+z7wnZxp/97ebEjELAmLrAIGqSUhboC
9zYPETwZNJ2kw7jw+X+K+agKdAbED55c1TXWP/l0+bh0La5coUqxHStpZGM2JluD
r7aJvU10/q4CY5RURYALF3ziwe1Q3aXCpLY2hFi+1KqlefgQYEINla+8JY/uZZYz
2b2qPZJ4Q3JhgbT4bjV5ZhWuXE+gog6gyYAJ7OVUL0B3A/o7+QrV7XWAjR8q/2q1
/UaU6AYfuPxr7bQDAY4OrdNXmhrrpKCq4Tn6jnShphVGIxi83k1JubB6jcwarlN/
IobUy/eWtStdaevOp3wSjuV8ZNFVO1xq0cit8D24OBKrkYfdBZLzZJ9LaFbOCV9o
WFYORRZEBf+H/AcZXk0pIzurvTJZjyLSU82x0Z3Ln4LOaqw7AGwuiwE0pebH2EOV
iqJwkK81vLYauV/8VOc0YfcAv0k87Y6C6YWGmCwoiH9yhR2CZEAFxNrIZMcVgW9d
C9PVZSAo8qhu1B4T8ar+1caA2+/qme970vlMJKd8A/EcJRgnlxlV18IV1J/hX57j
4hdpJcaPLLVJhq+NYpXfxW70+uYTvgZdqdmh9WXP/mioaULAfj+jPEQL+7X+9Is9
utT9qSpv7O5NrxZsTtBVdDDDuX3nrxCsOTUHCp+CUAE8EdVR8Q4T7cWkUtuEINV6
7AOVnogXJBkrozdGL8+zfZ8ZrgOxvr5BBtQcP38TDl0Z0oNe5n0aoxGlli6x6+i2
N+c3499dhHLMFuv5XVjpVxEUgN6YuPHhaQa+UrkP9r28hgNFE78WHxEvSQQ0UKZ2
xyt8e9DNnH+p1CbqAsTdYeLqDF6odFn4ctkDxXo9DAHlh/7ZeD8CQKVsKBwq7H7n
iXaiEH7i35Rj1uQisGgA6TOc3PnryPyTOw1HZpP0PNnJx21mSC9I2iVTJ1mL8nWo
R2I2L8BIDj0TR88yJuUxebzKqfz3bS7ODIOSpKmYk53f15xyO6SJrHLAwBtfqxSh
WFmLWbGBD9w7l1FoN82zEhwsZct5RqeXBgqWr5hebKehZcsgfXKwe2GJuRjiJbG3
azqAJG1C1Mi/w/QRoByz3GJU7qE4DSiKlaev+Sc7i1doydmn3B87jBVUmzxptqMQ
ycOneK8fgV6F2Ufa0fM+ZGxZm1k7JNi5KDrYFLzPNcD74LhhU1d8looVR9qlkWzv
KwcoAs1iXXe5ckX4WWoqfT2qAHr7nQsDgmWz7CPn6fS45gsSmR9cxq+ZaB1CPZis
8sqbvjQcooDCbhRGIG0GHhiXU2x3xfHNF53uIjwfX5+wnpj5xW68fl254CdWOlw/
QNxPByFUYUhuYoF8a5m+GaJqlB6MJXS80/jFgR6UZNv77qWtzRD2meN6p7MgPAsa
8g5S0XWNISgjxOVUPPjSzszA4Lk1KCUWe2+uGndB1ucsPSY2QPHQHI6dh9sghhS0
rZWVgd5Og9vp4xKB76lClJDnHF8lJpJ9OmwhiuPdszlq5Ls848r5Zir3kTlZNHat
P+AavriFaC6AwSQ4GaIy5DR0GzCIp7EiGdB0dWk2j2iKjiLOAeNmJ2EwaeQyEpZG
U7eU8IB7zuxjcV7Q2jGG3kgiC6zbnQEpPk/uKwtEOU+d4FOzx+P7aCUm7uPxF3mz
G8YDF9KTG4r5eR5kQgJ/nvC8Xx3iSP+3suxkvEkT83X9V3lmLbj+P52UH/VwnFjW
snqKIFXMZzXmy7zA2s0zBUjIBR3V3RwDCHTkGLu9Hr21oiVngpveFAjfhNiq7V/f
HcyZif3GKl4rLnQo9ktqY4ReFEM3SroD49MgBW61EQzXqgfb+FRQAsGAfizWSeHK
MfSIHE/3hYXaFVwqkBwLHXY/uOm3ITRe6eJQ2WFB7IAxqNO/ecB/mCjJa48HJi+K
xmc113i0j250idCf2fbF9qI7D4hdIMmbI1dllvDjPnO7AZKVqOHszrXJ5YZT5f08
Od7EG18G2hOi1evoJWTC737HPXlmOcyR4nKgGMYlomStsU0jI8pjaXPW8J61MUzC
WNLoVxMq2bb+stODdSJynLegrUq9di1nJw90ZrAhztUgz1aOIoONtg0rHZgVdGmK
i7Ns8p+JoMY2nrArIw008KGxCr7UlMND+p4rqOgvolv66rKWqBlMmvQ3MvQZLIDP
gI54CPwXchj1PPPIn1wvOgmq0jqESgd6edRSfFKclgKlQm86u7o/OOmC1nJGh5qA
oNBh4m8Cc6pG+zVN+Fm2vRGPqWjrVrZTkkDgtzBxDKyrBDYtb4ULBNgdQ6RY2+YQ
wl4TrN5ELNsmjwUILUS9M3tWmyOXxPPLqYldPASmmEne1oTYPFwaDGpE/BjXglYv
2fGywR3T4DYoc8XV8co9oa6EihC6ZLGn96Xt0N16KCuy4kQqZG5kEC1njeH/OSgP
W5EEy7m+YfQFM7Fm102STU8XQ4diNeB/V4LyOGtZJAinGukPPTMxXshy30jdb2FQ
MaP6s29jbdK8rx24yoHqeqQg3aA7JX1/wv7Wx9iT3rrNLlpUBny1IXKeUlZAXKKX
a54PsZ4tEMsYXfZ1Slr0GIeJqKuisDFbiwv3PTOPN5EBGn1AlrPqfcsFs8RLcnuM
T5bzoq9jyZL0viO0CTnDNFaEbN4cZ6ek5RPlHvgB2uU0QfruA6/TKAbLQaFezK+q
f/lDLBfnoN0D08IOedz1pHukHFx0WrIVi9TDecBBnof7hDHNNocRn4QkrOEJjoDJ
UR9yF1nH++lWuG9BLSlArclJL04OCr+oyH/vQ0rlBjFcEsgjcoHL0MSrmoq4LjjJ
i5i1lhym2r3VABlO+CM2KZr4xBGbRJiFwEucPbG1rsSCiB3UB8BQCPtUiJhwcM21
RA7IFUSRm/n0Jsn+0wRh9mGld9sZSXY1qOD7sIcB4OsSyq9CThbwoA5BDUdXhGGR
rj6S6eJ3ia1jor2unQY88xUKp+U2dF9ePzD9AN7NdkUKEJWHi88xzVghZNvHvyeA
/uxLT+KT0wquHkqqWKCzGYei45f6oseziO9qsT8TOSefb/lAb5q+OTTZcQCJDZiJ
brkWSP1NMbIeIW3W5PdY5vslNwlEUUepZYrLDsCd8LYX9ThuQ3TTs9fE8dfIY3CO
rst8dFTHD1F6D6mZ5AgXzQiWLqO0cMvcaRuZt9sHfelB6XT783kh+DmhHrih/UqE
2NGnIkifFTcLVsTfXChaZIjfDdtOxsNyebw/GOOS2m2Xkqm6yNxyQ+5uwmUPZ/TL
KKGt4WtSilUOkmrSZEc5gfFzarz9K5bNNRGcezY23Bhoaaxq8y+cZpGdabPXCXAZ
0Q+1hAYkWMcABRtwdSifRbUwzdafZpBqEB5teLcKofj/PfwwOnUQgDthD8hEXaut
3C57h9Vea+5KaDagvGTtXFmXh+axHhy/ONWvyE9LaeX0jwMtLSbLUXmE7nsZSutC
cKeCPIu3MYC9LokPmPVidmYyrh0nU5KYJr7FEXvSU5nac+2A4hvOJ63N7Jj1lqGP
BvrGSTTt1ACOd0DnJ0sgmofk657JYhq/OHiZUbeCKYH/H7VLuLXH5kYONY+zpJM6
/Ywawbyvcju5sYbLAjnWEBPwmwX/QhiFCxx9LgCTGcnt15D6UHPH22Zw1y3aVtXW
X1vL40gr9RlPyNdNqBCt1mCeHiQocUTW3WGv49bWu4HhDYF2JFnJJfW3kAn75eTs
fBzIhcnWcgLJmuLV0CVBqvj2ZlqBN4tfpQCY5NMaD4NPJltblKiU5mm1WgeIr8Uq
NqNiwHbuZ/TztgwGRNm7A5yFtWPH5W/uctvt1+4r86AQUYUmb12djIn2IzCL+4V9
k8ucx5pPwJgLSw7eAuqyfdkzErlpXtn5TQ/eomwag0h5nm/r6VeR8N81m8Ow19bK
rq5AKTvoKPk9X6ooD7t57/8DO//LBHhz82Pp7mm2f9qRP3IJC12Be+RgzCx1Pg3j
S6JfmIriVzxDA8w4FdSVc9Kdo7Zr9Gh3lOY5dQUiFzdY2OZNFccjMlJAvIDQ2ogu
ovJtgTS32gLNO3261M/4HrENPSuohil8ub+61oj442565LyuR/k9sCM+D0HlYDmZ
fW5HhN/o72nXPTVzzTcYyOn0N4pBNzC3Zo7FMgCWmel0HyeHBr1AXy8g6lnKavXu
gSAT8afiEfm4Vw9w8blJDQfkRI0rcG7fLpT4rawBof6mQ9IsPpVWfBZTqqxDBSPh
6O4LuXKIdQjBkv8aDP64j6kn4nKqe52EwMVXwzyNfM5VrViLTx2BE4bVuGs/Xbh5
/hLIq3qNkpXK5yIkPdtERfCQjIbcPezYkqIp4tW8ELrRh6HMH2a5KLCkNqBnLlj8
zIrRwsMtggppuNHmvcZuiOsPWom+M/TnCUjz4CdlXRPn9klMUue7hLkQovtm2nUu
SvrCVCdw3fHDlIpKF0c1lKOP+vJpGtSXMoaN1r+qeI75WEBPjlBxx9UVowjNRgIp
ubapX96YbAKhFpPBASmUfcAEOi3/nn/YJffH2AH3Lt3aROoeiuAQtn/2iY/4Lr+N
AYOgdoi8catrv/uNyF1gq5GDfxYwmsBFeRT7cMjx1myDUGhoqKIZZj49Qmk5co0C
watrnDKef/4FN0zEGSn+xUhgq9IQvXCpJVD6f1jeJRc8+PyZ6nN7iwNK/7jCo80g
ILO+Fy0RnBufb/viJiRmKTuU5wAISOvllIQ236QlL49dQGzgUVC+tvJDgFn99f3Y
57Nv0hq9q+M7kfRZgnSqgMgC4FyRjgUWUoQGK3Z4pdRZ/pqrGvpOoUawroq7lcVl
CmFFFV1l6iqANVE0zfsM9AtGIMucI2isQgsWk6E7PseAwaJz4tVZ976/PcKlDpdW
EZq8qYuWmz+oGJnVZLumUkCovICxdQH1YYRy5SLH96A3Onjx1GidJZz2MFStZOBJ
pOnCfurJ6AJ5jFqx9avK9kjyAhLlOToluDN3AVkkZ9YBZlX+hRpPCAsP+HmVMpta
EdfT0BbNq8aISx2ID40lajKpn4ISEq29eJcE+VQ1Rw2PJn+E18HnbMA9xQD6/oFa
xSGXBnSlDTMQvrs6YYkFg7qgWvzumJGrykAW9D3S1DeahV3uvNSGlN91fsimM6QX
kndXhabXIT0myQpdCEOYDlOkEaLNeY9I47NmeMU/m/TdzWBwZZsqGDiQ1/OuxAB3
ukneAGKs1yxfQc38tHgNa81D7YbzgTlCVZ4j5U40HipFg3fjdmyheTcsQCZ7smL6
bsPXeKkE06PzD26CRc05Tnwhkrwe/4jnpG0cdyPcCCtrX2RPALk4xl11zSUmYvuZ
lOQAr5oC4wx6nvH7g1hh/WKOhP4pv3L3c7a4GVpKvXaNtnkXyf4Y8tOWf4z9Cd1n
qV4HOAXAzBHp6X5IkXAv3j5rZUbBA2YmYHHtkT4GhHZFueZ8FmYZc7K0EvV/TUJt
KGG6zPWWxTMWPurBDWNTrOa2k8Y0q3gkbHuxM8kX/FEa7O8FD6hqdavCSPNH524D
CsXoaP00xPjFMP+xzW5OPN9C9k4kAqY4SY87fCYidQZAJMMpU29tbqQPdKq36Qyp
Z5j2uigXl04Imf0T5wGs3vB1Hx1occERImJwlMS5e/+T6tCLvnjPZAeHbVxOZAFC
S8Jtv8Bp/pFmm1dnoLuaPQ5t4wg/WwuB225+X2em7owP83qDgCzEFLoZ2n2dWVVC
8rwhhk+NNeXdFr4rNu43v4XjkgNVd0JpGIVRtLSyRA28J3P0fWHQjoiitxxbTOy9
nFBDYYh/tUkhPmZWosVc9pQguruk9WA6INWMpHdfuKCv70isuqJVy3Awdg4dXnXf
dW4gv7t+/4hngk9vK/9ZxMVjjSP/48+cRdbwIWL7Ij1Q/kLNCpQbCCPcKLnFz0rg
nWLFenFcN7IKRaAA3mHtMGt0qSsmAUF10dyNxJRVoUy+avSoyeZsc7UuerUSr2WN
0BGjPPD9Ve+9KAObNM1vc9j8TlcfZuXJxvFDDChriCnyMCd1O7H9Lp77TuR+HBBz
eABz93Zo3fKG2OrDh+4FYGOPQ4NE2FkPGY6IYp0AIIo=
`pragma protect end_protected

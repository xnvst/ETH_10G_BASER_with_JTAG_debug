// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K94XVGcO0gM25br1M1fY9FFXGeRb7EhxTOug1J6x6O1+QB++Saaeio81/1+0o79S
BK0z6Wxpg3oXnojAswew9dWhIJ3zymtuA+rVZnnskCX7F8xOBOds5W4xyKasNRHr
vYTqZ+k5ScCUkYcRdWzim6AWuum1kBkVxPYItM0E6MA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26288)
9WqWE1t2R5bG6hEj5UqtAg/iuWDmtODbYbnMMxGs+ZY+xV1nMQVbPeV7cniUV1+8
SbrBexy56mN8o8+ZvTPdXvrHw3nzZ7C1KIT+/BxjEkD/jzFdwNUBRy1HlOEi5cUv
CZceIcVNLg/aGn8CsBsEJIdymhgWljJjK+QO9w/W69kEEH86dkSflsaL3j5pHNhx
YHFNrlfHmtMPszo70cZdAkIi0qEOk8VAKpREZDYUzaga/D0Lap1mrW5hwWndDJ2Q
GsN2O6tXCoyPa6zZCDrdoxuChoWAVaeb3h5Dcfrmh7f6dmlRb+3PVcCUKWhfaSar
gzcEn49NZk4Pg4O4tYVxAoIhrz3Txye0GnSy1Fy2sNCQV1rUyh5Zz/uhUq1Mf8+2
1k9VxOmZ2ozSzGK1EWhtTQTstF/WoCQXA1vh8GXkTKVsVj/XBODVmih37rnQbgw+
U4cfUPWWZ3kV7SLWpTx0zm3v/OZHxQRTwBcY85NwyARK3aaC3iuf9NBeuJcrgeEi
Q/N6MGsjNbYZItS2woIXnMwLvWsG2/fNlqViCnzAare6PNMIUFMd8VXSjicypJII
mbmn6FKU2BWP3ixUV01Pe7Puq1sppynFORtofdXEKPPw/nmR6TiAdrHh8SqHWQfj
AGpLPEMNlL/OQDZ5UoEZr0wowE3mFttmLnzMsU96VL1SICGiaIe6WInN2hVoDIR+
OiS6wxIkr/iSICOy6nTGPGdBGohlaIBvrtVNSYVkyX4/n698q6/3D45EeqeZcRi/
kyh2VG4VtJOf3vZhT6+haby/OHuq4T31rUcThuE2Ab9I1Q8h2PL1TH+HuISDl8R5
idhqFjyO/FA/Jbyxs9L/VyyV66r01AvoKwkqsgkhe5vrKj/r0VtA6OJErkkJVcI7
e47Nh/ddargnjEuVzY3PWqExPHb4LUdt1qBqAhVykUKP6+cba6dYhM6aA4VqEiXB
uGuMXtyY30pLQC9UZE51zPJNrBgRpiVkOa0h+Fv0SaEUHXJa2QMgok+T48J1/pD7
dUW1l7EiH3Mv7gdMSYS4guVAv18AEEXI4gJTTx0HoFqguJyDYNitsCxn/s5zp2Ev
mVS69BR+6BH2q0E4adsfwYhwnO/SJIPexzGglwjSkBv9ApJ0BR5WYK2pyhWP21Ad
U5mcA1B+AIDL8aII7JTU/gMU/3ZCbbZG2UJ1BLLmvQZ94ZesCdrYo5BYcO8pEH3t
ubva7IGERAcOMBeJjbZC4IJxjDvm5o4avcxWwJ7csMID8UudRxqBY0q/2he160cw
Lc7qlEJcSBcUJBzYQlW1VOYocKLT5CaH3IkDeA0w37mhh6x2UqUKt2Gz4HeFiTpr
Yvh2gycQt1dOnWqA/ZIJluquHjusgU81Pj/FRE8dNGKaiOn4NLPCoKh1yfcAvHgC
qx1hdj52dbIEY1w9OJEVAsd+c3o93BZbWEwcrOwJQNQjqiRjLKK4hSqDYiG1GVLR
Fjc6T3vmt/TDfnE3uwSvi/skmzW0ptK6sAOolQg/MQUHGVVKUJUEm7oqo1weaszp
YkLnIqn7GjfmiuB1WC6Blo65fqRmXsGZGO5aSt4NAycsiPSmhM6Wl26uG4i6IKad
0W7oLXPPV0AEBeLiSjZj0698ya1HpEKSp2aROjuJMumwx7wVcCSwLbEtXeYNtD8X
uZl/cX7xV80EVhyZwu9tLkfFC6SahbNFMkWsd5yC7BJOe1w0BgAmf32MG1YUT8Y0
c1xSt8hceWmgtuMmVkTEPNV5dwHPGAULjbBLChCfsWih/MoLnfHpAwLeii4KbOqm
ziRMSE2gf4ndeHk8ZxYue3V1uy5PzzAIxyD5umRNkY6fK8045R0jCqrn/BY5+dkG
9ZQKT53chQw/ZXt+XHwHpd+Dfb4CpwJpFLZT529x0o9WfLpNNVtK6jaZMZgOmIor
bEmCW8tISABkRcUuUbC80DkTt4yT0N5/XOm//sKbqiJIZooDoKHNg3MjZSMy6eUl
Mu07U0NvrnHx/GAyjronCF1B/rh4Jq5C3DvoPm7BL4C32gXiI28Wau7OuNRvX1tp
d8UJ5jE2iuhrdkZ3ndYHyXMG3YjOPgMImy9Y7P2/a8a7m7GZIw1+0A944vwmCrm0
6PC7p5M5zNdx71+jyfh/vkQL9E3xsrVxTmFhjBntn0Zb2QP3InJHKNCeCRMmQKiQ
wRwoy3ODWEjWHuWnLUn1LQAFRSlRdEVSWW41+eI82quBbVM/GjNsLUuUARUIvTfr
WOLiUjWiwGyjRI52wPxzRQgC2sdjJReiN576H8sXmjhjdvNowxxEEZA5koRafT/0
boQFWjot1KhYGa1qUItBohs4IUoVOR1X5bhau5DNF+liBMdj5B5DeIkoCvvIi2Ti
SHIyYsBRJBUwPi2Ggk+0Y43E2F3SkXEV8tOtqOUs+o9mDZ1w5RvxcCkHlJzpDFQb
E9sf+nAeA8eIxNYW2qMloaJJQH3x1tVJe3cuwvtsk9dk11PFxdpbnXrwZ4FdwSRe
MTKjUSW4n1aryOSJSalmd8yvVHrJadTYKKg5wuG8S2+0bJeUoGIjDNmTHPifaO6n
4X/e+31A4U0g5fWI6yJ9zrybSpjYQAj1jivuGjRJdxI7tsNaImRzz+bmuOvT1D6H
mSUHQaKg2WXDT0C9bkpBsttmIGezJPrN25qUVjsNVNVfPPki2bowctF9eUZyPv+i
7cHO2u8OnusTWBOWTK3j+zPuqbqlA4TQa5DQEN4uwZtiIVWkA6pYHOAjZExcQ6+o
YIBwOd9G4fIG+Gu50fiF5pW+gO3WSnhbiRJ1tYNHWKSTK+i9mEGzGlUBgQXmnz5R
rxpFMotKJYQxmA2cv62brjaU4Lg7P3AB5aaGzUU8nRiHKHucZqaog5N2+m9fQ2CY
MRYTs6rBTRiXBCkXekTgIYLWnBZlaPy+VmyRI+1U44l2UlalzLjL98UGlNSbJIny
kUEwqfb4G8/I8FvOFZA0KyvfEpbFyCb3fJyAuxkxfskJLy0RuxL6Q3cf6uCGTxaa
nng8lORhZYzyFgPYppjccTg8nYA0KhC+ImjwWSxCUZ+Nz+1Xi1r4P0Dv3HqYlMaf
EnCxswyN777Efh+DMt1OVQNrTEC1y5r49NAeLx7GyJp5Kf3W2La8uBsADp8G29bS
LZEXeUSes5bz778ZnPk6ReAXMTfpQ0jVp8oZTrrl1dLqkDOZLzvYoHlJJ/xa1yGb
Zlm518R/frGXNrBfQ8Y4ChsJvn7nUDYX7Yh7DkxTjGrbols5biLhamapbPe+9Gcw
8Fddh2N/ejCDObETThKRuHdo9XSGKR3bZK5bqAEoFbGLhuj6XkqhuArwP5jI8n7b
bJGU9oQlLXlwnsUg4lBKgvlT6vV56jveC6eh9j9qOrmfuwenSFKZxbn9UqNML1KY
gpM0a93E4aBB0shgPaImbM+1mWSu2nUyCWI4ut0UX+X3kq0pasC3zfGjXngp5YWO
cKCO2KaZawaflf5F9cGY8r6mgN/OFYAC04KF07Mf4cpaw54Qb7tpih7Mpwwc6C3j
Vz2n8hY+4ShCIEUCsDO15ANIpLupu0hlwb4PC1sfmjhhFsLQt9FzEegHpN/k/dLI
15iKfUGYXq+ozE1I/s5JhbvytJuAJMwOAt0IO9ZpziH1KwKlt3MotvIggXMaGnS1
pgHv9GOGzyo1E/aT+jDFEJVLNZSqjUUERRqyJ2MSoo8PwVmb3fBNZSqtEtmKg41v
RYql2Lq5zQf84MDojsgiMdKL4h/Su0LarCdrcw7AfwsWDDnhNlBxS6ayQdda8hRw
f8KfUNeh/H41Xbe4SeFIs8B+iTKe4uJggNvvZvmurNOSIER/VJ49lN/lOHuvHR+X
6YVm9m8ACXckmzyBtv2usWdf5XMRyQm+2CcjfXej4OgfCiCM09sg2VHeUM11ROvH
EHZtkNhoNlA7OclsgR0qDP4JMdKuaH0Ybtb9vBj9QLFiVMv4Rt2y37KFAtEeWC67
OJN3spYii4TvlTocdUqhp0bMJWlSplF6iVSzl2KIS8La55kfFEnZUm1YJDQDa6WN
gjDEjGqkG8FE8xumQivK/Jww2sxXKVzNUsrSoTRNZP2LUsjiqwSxvdZhlJ6KYDpo
eBgektMXTDDpwbPrnsSQm2g5p0mpmrLwLIimqxxADvndnC9jDIlhlqzXBID73PYZ
kHLY1PW4OQEOLb0y2WY4Y9sr9Cdsly8GFCXHxww0dUmeH4IwUJyhB+svOiXEx9rO
5s0qSSV7NMJa//VZFn13XhTD+01MTvvtT19dcI6Cex3c+bzOQF5l8oducZLOqCGA
Br7q6WK5aR/CjhwBBgUzIZ25xzpAE+kCWIbVzmv6Fz4j2O90VScjde16MY4BjZhZ
nqesGknxZZ3F+LMMYAt+MbWlOceRz/AFIkxuWR7+R7glPQ5PdMLPQX7kKvXrIzS1
3WZ8Hu5tY/yzl/MZsy8slDRnrwtFR+iOSyd0jT2WijgZYjDQBqBTHJXbzrnbByHy
dIVKT0fHB3ihLjzMZgpInJnKw7F251b/1r0UUrdGxy1niRrHecs0xKMILOtQLo0d
GOlv0cWCcrLFC5OHFMoarhAD2Zu7CXG1PO/wDk/y/96CpnQM0074qaATlwWHUox1
rDRvjWCkhouxq9eKnEiSAKjpMjR1+QME0oqbwDJeDF2dvIN7PnIhSzrgw/IBD/rL
qJ5YqrPDmzpPA69s6cHzkVJs2d2CONRuLalgsHp88IfrhHgs/q35W3gihxdKBIrq
TOnPOb7upJcrIxJ2g6wIs9bEQ1s/XTNztXZ0PtV1CAOSVAtsVTzFfLz3Q13C25Uz
5E1ODw9/i96J5IkAAPgm5GVAarzCmih5YQ1f+mg8p6lnHq5NKw8MHLgCqSQ9AgRQ
7dtsGLLmq0BC6UCKaieO+A2PsZKmFUlLRpT2ailpV4qY2ew0QLQWQD2FoK7Elk23
6OLNjcqtx8f3iaJ1U5DCHIsPu5jkp2Z2id61EF/1IeKSw+5UJ1/N5YUFOc/6d2Y3
8Qd3ZpFT/KHTINTtapcrdPrE8YNWhq5kBaA3x57zlWbedAGCGsdXBW1v4JEWsuHr
d0kOkLUjVhw3hWDZXZh2drDZprSbRKwV0kx+Ed8nV9NzKWcf4QG8i70syVTDruDQ
W35ZONkq4XCJw5mX1iMVZRp4xb7B5P/TzinPJv2t6seYjMwFMzgQinborqTeFGSB
WA8y2I8ENyeG54Rz76KvGvRQs+hrmllwjVeJS/9wC8ZdcxQrYqqL9+GfrFnHWrhd
rSZa0DJ7RdOU1uo/qJhvxynK4GjQx4UU8k3tPGK4xwfY0IqgnXWeAZxZO9UKrGMo
js/EsD4MnxrNUtliiP1vGhD/4ZZ1ZD/TXBfnO1t6G1VmDS8Ae2s2IPR+tYvDzAfu
DS2NLBzSUb5Iby7VYMu2ztV5tDOWNFUKLAELho/sa/pJEmTzoQptr9MCzjH/9OqQ
J68b/n550gp6XvdyECdKW16Ls4q5ZYZL6rYbBJruBkNz/x4ZOco2RI8mmNKr1nVP
KeeQkwayWRRltm/9SI8LCAzpRM6OkbNeTLI/6Mmwy0jsAOQp9spRgHZMz6fWY3kd
wsZ48cqZZgZhT9gYlsdwkDe3+Uf4BwpUDAveG9cpHFOS4NHHhVf9RhH8FBhCn4Vo
DAYyjdTzCo+z65iqvj+f5MHuy/6pyzn6v32l3SaqCji9bGaBVVqrK4X9/Ys1dtdE
sIOAcL25WXkifnao8CfEgttTbSc5UzyHDvFOb6y41NIGgPX8TcnznKcQPum+jMQE
F9p7sBT/0HsHnhqzzN+Q8JLCciFHh4R6l13OyA10xI4D304308RYoXhsSkT3y4Bk
v9RvQ0GM9JLZjA9ORpkxol6sik4nz3PBxhgRK/LeoZOcC0JgjIa/Bh5bGa1nXeAY
Bg681gimnGr73y+xTu7Ts8oLAYFgrlF1W062LEgAyKgputeekHG5ZgEaymA4sf0A
vAKHjbrNSpmAoYIZEXlbdezg34ZrMMPqc1/Fv3o5UwA3SROREsnKa6tzQpNRf+7K
0SHXGCAZl9nMwpHP2fpBsXuoHetDZ1QC87dSOn3jGeBQykQJJN0R1ZqoeUNdC0q3
8QEG/RGQ0OUO8XJuUnqZj54QeZxI5DsApNHk8lLaUS/0jgSnkeTzZSk+yaYY5EA+
S9410OtexxS8cEFdG8OF6iQZW5qhOb+JmbOExQXNSJfUYkAGfG0pb/UxCA+9x10w
lyC0qeyU0eUI7EcLheGlx/dLOtkc7UIAE7rBA4g1vE6B5JdHLf+h1V4si6BHVR52
evcp/PWaSx76QzHqMNW5LlZ1FN4Up/OQWcg9Cjy1xPpbU0ry2lhwsptpA43Wi5De
Nvm0JB2KrqrERfnwiGNGp8oHY6QC5bP8dT8O46Mb7NkC1Dgbu0HYUFh+ndgpR1Dd
vkUTA2Z5BUvMmZyb7TIHn68JQ6XsXEEtHwG+xgKIz9LkHpbIWNbfSZaWMxTcV15r
uH9X/j/bZpBnORa2kYD9cAI8jhseaFP0CWRbMVuvf/tcbard4qcnAqlrVQ2lwC8i
qqyH3YR6vF0/0AdreE3LUmx+DwIur6pHJdjBDURvNgaW6lGQW8rtEM8eBiDVz/XX
NBRFqGFp6bRnDE+33868EmRvYWktMB3rBaFCW6KZtcZuk9qjFbYGPYhniruCA2cG
atBYsM5BUzKTSD5lxZOE4Tr4L5/g4JMKEmB1labztf9Uh1M6KUPzjnwgyu+n2s8E
0U66LAm9biXyxZpFU/b7vKKjYMoHm1l5CbV26XVpPXz2igI7CymCNwVXFngNfvPx
AmSNR4gC0DtHGfUUl7yxOQ+mmxgthTxUGUsnoYDKXp12kpisgbm/2hxx2NYNNIvi
raph9UhOdCbX3q6gLLmb2Ze+0/LtFMIBkWBms68OayeNs6kSoNQuPAz11Gw9/FQt
IIfftg9yzvJaiCoQia85X4yr70N3eOM1L8HnCo05TK/XT5DHwJ5tcTIl4mWd2fmE
4QpWXBPkoBR4XX+anvPXxwYbZ2W5Oyb1zWqRtzkL4XuNtjUlTJjibuSxmilnQeXz
eQqIUq/mziaXAAK0NaV9Uy+xwdXfzFeIBn+Eaj9hXWe/t9yP0mprk0aqZDjwrbp/
RE9j+1/0yciLDRuUYj/79m0DtR1cZSHid4A3aCLmixBqlRnWvCiYqa3SQj3JKkmN
1tfEibN11hLK6IQe47xLXd8c7i9gis2Q+PLh6LuqYSUDyJI1VfkYsnpet4EIR9dK
cnCJcWi28ljLN8sqUdwwgYLNGpqBgL8A5gkNqatFuv0XfShnFK9rGDnh3I5J7RAM
dc3uXZZaCiAO+TzQsc/hYJLdevr99C6VpEIORQnY1vp98VHfX98I6hpMVSoHoP2J
faTWqWiaej6x/x8Si/TBIHSUfC2vXj1hy2dDIXWiJefgSN8cB27RoSSzJ6NDG/or
rxD1NY5nCQxlx6hjdI6Z65pagRXaG3IYhbfrJemL05XfUFxh/NqaDGm/QKr2YXT3
YZjWa57mIee0/XSY3LftgGWxiaEIRofPSpYC6l5GLFNUMJ9SX1nvFyWEG/DafUMP
85rxLTOlSYVmcWxCXhiKo9fDyeJlZ1y/uMsJ4AoA1l/XLG31kIjUQLuf3Tlh9R51
x3u/0h0EtzAbioTd+w4y1yZR2TD242sG6l7Jx6EonvSW8Ku4jtBiUbXf0P/TiBV6
mk2oalG8cw62Fv+edtI7vv4/PEo8VBqN2hg3A4wQp2pd80fKF5UnYSCeXra55YgO
HKDET79oFDw1BcLkNv+2kzNeTgmcIP0hRrvRrVaZcfVZeX2ouK6ibZdBQnc2PD3Z
bEBeiPUh3iWoEZYHzzls9SEhZ3kmETN2qc4iUHrR7o6zo8R0v3zlJdarMlb1fLVb
ma/LPwHyLv6y5NjWs9ZR+Xl3CmwlJGbOBHEyAMs+XndUAcbOsIeyRkmZ6GuYGdVq
y/0YO4LJiPLGgYODK+jAPJYU2NDE68NEcE3WnAitkux2RAyGYQT4UK+fZkML1n3j
Y9e/Ql8kjhktzD42MQy1RxFXdUJoK/GUUSCybcqQhpwFbZtOd+P0mBZRoSI/y64e
SP18hF7/IlM5/Bu6uZsIzuClhbjT3/1czAPuRR6dhowWhV3BrlkCmON15UZrmhUE
eRO5xMyTt8zm+/qHe7fdWLW8fZXGXVcHBF4a54+ZfCwf/R5rsiRgNbAwS98etCaL
r1dIa8yQUXWFlKCsUzkIfjMXw5rO1AQZuXMHl42ro9FlFEjJMwYudgrJTfjpINZa
T2YPUJp03+WPtTJ0OvEPsI55whfc6XR6jf30LceJyKIMQauqUq6z5C71J0GSEdmh
QwPbcc26EJo1m66kUTQ9bf7m6vYEL6jSaxzqOhyAe4KTqFwjkGDjNqNGh81QwKny
aXz70hwGcoLh/FE1W6i9S86KIQgYs/af1bPaqd6jB34kTwu2gcC5S9vqg+GV+yCz
tsczaI1dPd0v11NXhD2gbE9ncVflOk1zcrerfcRlTXF4yzYi0O+JVyLJZLqWiVPY
CTSiY+cPUP77zpZVfQnuyB/L45KKEHCrZcddZY/x8MWF17bCJbWBuVbVvu1NgxPF
O/zApWNcqdo+FOvTPAbjpPO4WIduTV4hrnIvolpAj+YqnNgbnVGwP5/l3CUyjAkd
6NnLxS0R7ZwKYRDDBfnx7eFgOHG9YU8qWC0GFHDwPo0NftGvn3Cnerk761CuDiqM
O4736qwVCHrfAo/1oU+8CPjyRpy6L72ltnKEywEb/RmuJroHFNjsbV8Z/WKJ6t62
w+VsVLT52yXDxjMwB8Z/y4EDokB6sJonT9lGTy89RjSrX77zvVUMo0C0/MrPXLlk
7XqwlGviDcrddUORASbMNksbLh4gLCnWjLG4OAJhrIQrQZ1WvCHnr7/gaBpanB0f
gYmbIQ9oKJ+rWzk8uXAs4n0XrS+qm5GkhKT3fUNXa/fcIpmoabCDrhwjweJvNDJp
DnwoHgRlxn89ZYDizOcIKFjWW++n37J56i1f/bybW7PhPcKR4e6dowFcwJGOPG7T
7rHCM6scsMgcp/jH1LnJZ8I57+EbVpla2eNrh37TFNCzfc5tKr5te5zgtJlzsLiV
Iiq54yvSeIWca7k+FZeQg8jIoEfusV/HV9d8PSbjpdmi8+XtrvnC0oIuMRMY/byh
n7UQyCZ5jO7fn77JoD1mZpNpHBQ/yR6Lqa4+BUl1KdVrhaMyPn/BmPyJ+jFsA7WN
iXLqqoNKRB5FKERzPXPjDfqoA8/zHfFW/aGWdcnzEZgOQFPMBqqdGS2RVSHtaYSX
tARtCagtRij+/yZ8uUjGfqaNyEpLKhzWNnLzeLuG8pwkRPf6w0a74Da3Anepfr/g
dZjeWycuZF8DZbn/OmvS3+UiqN7JaVtpQd7iB59TABTmLHQtNmQr4uz5dSo4eyra
Ssm763QvG73H18rq5BePIIrKvXIzcMJ+r1iMQUh8tEpBCaFDl/zzsB7idFMGUgf/
lPBUnc+kcnOnUbLRMlbrQxOIR4tjOd6TS67TqbUmC/N2thUS82nJivizE8ZyFKfO
bZVHuve0rLkyIHQJ1fJwnoMqiyUZyamT2CLi4MeEceOgTS4c7x8uXdw4EzDJESUz
7c/uondjgJi3yeWglPtBehw6tX4pp1F6iutehJ+mqhTbevkso9Ql0svLVwEe0loL
Hv7UYvt1uCFzSNL4zbJ7v4xvMk1yFGCoTCGw/yrr8C1iN+KFvBcGxoA5Fj+OA4CR
xcw3zMWe1hndUyoTxUA7lmp34qi25hFNhrKCpxwWJfbXUNmlR2WaBItFdU14bpE9
3R3c11xu5j4pRqx5mqROrF2YzmA+APl3HbyW5bK7RAeWEmg+jMunTeTPJLPd3jRa
fEjPrWrd840SyATtEZzsXNbm4hkzjjsw92QNEa7DS2VeCieC+MPhYPjrrC7WuP3v
BTrsc+bnQlDUm04WXs35kL6VW3e/SITiy0U0eKDWcbE6fvLApNsBC+vLVN9y1iH4
keYJF92Gr6cdW49+9CjlwH+S5FZuxOYgjhAinh5xbgy+MFJ/pBkihVf6M8bTwIHZ
Aau7ahXsLj8nFk0k2t8bI0nzClB0+xc4Zf/7rVGwWn0RK4sshP+vd2FY3r4wwoUq
bpRM2EnqXPY4ATTAJj8s5fXCdxfB8u/flr30xhyGwOVqXHGlWIsXUpQds9cphUUK
ZisHEWuRFIJam9IXce+bfAsLK2g4To4RomfWQlr7x5uX/M7f4CFhsZK4w/CRMOPO
cvn3er7bcgY+39lCZUkpB2tk2MEQtQurEC+p3CZT6f3XHdqLWkLpoBnzLs74IlDb
zc4XEH9qXMlxyGqRfxXTE+1a6INbFJSW8GzeN6BKG2B8Pej7Zhgt8nlzp8UiCFxw
Xz3n7wHxjQct/KWVrPw1L79HEbeVtIilIv6RjWsmcvLzZ665zzKRR9L02+zmD0Fc
4S/9Ak8W8GuBO+9Xo8Ic20n0qAWrswvKANOa3H1G49dfmOFwV2qfluy4QJl3BNvd
3MgXDbSgiw/N9UuSZvtlInORvB2fQ2+e+rLgUiv122vL2PK9J0yn8QpSjsVn3MK1
GizxGQHrFPQpF7hfEvwenLEv76pUmSUxq55ZnE4wCrN4f0cQ1maqbbmK/n6En1A4
FbJKfOgpilzVH9Kc5M2DOfYjtpIIol1bkG8aaqkzsgv28lWakPrVoFj4ger40FEt
5p7QwZ9Qw9EaG/7IwYxAGsGWXKzXdrR/QfX79TIVZK+ZpY7WsKoXBNVqP/BDZfRf
4wULSHG+6/cPtV0Fy2TlEfl2US4OVtpUwzo9GPbWTyS5yZPIF6xm3HfE7tA1RlGo
5Sq1/HpkDIaDLfpwazFHzGiTGB0V7HdNAVSfgwu9vbKPAhlw+/vWAwJskrbsgefO
wFzoJYY0yZJ9N7Z8wTdmdvQg+cBYFSRAC21nJgp+NRCEzX1wRngUljxX0AVde4fA
8zGBckGjWMXlOjOsHrqVgVrcEN1n9+dbPaSP4Ga4IjruJQAja8oP/TGih0xZdKrx
7uCFdKoB5E3eT0q+Emjclh3XUr4W/Tg/9hvRn/WstGB7wnIQKAB5f2qA2VanElVn
veD6e0bTHThE7khmJ0zO1G+FyEbLbtoPEsObyHW6NFsmSPua9IB9ZRnt9R1iKewt
ROKw2Hek1klkXiG67J2D1nc7HMDwn33PEyRkYDSRXXrdRoR3+0v3iHa9Sab33nSP
9Vrk79HsaGFFYyml3OBlOB+dEPxBzuve1pbzWPiUoTkZuGz6x7TTtTnQ8Xe3U4ka
VRFEm4jHC46GXzo4k740GnYQDEO9v0NX1bE+N7gDIvKYOq7CCEUBO9dhe2vKB+oA
l6y5UK6EbFEeINQYVBUuX9uOvlN96Kf+m2Wl5Qh2xwq55tWeeN0sfNzSd5ex6v0w
9pZCOg3nRTPLew39GC3whWj5Qbl2WcU2MMX8O3/660OtfzNeugG0n8gUcnFej9b2
NwujYxncWRi/WwWEyipz5L4Jxt2ny5RAqr84UgNsGI5GYAxbVHqdIl7dmjRJ+raF
xvTP9Wus1Y2FgWSoDJiYvM9V+wUHzK0aTtBUekcHqfrIj7iDdpdOBtgXEbrKvPjo
/TqkafldhT5zZxUW1Gi4DDyPRIJNDWeZK9tqgLcEBm+mG6YEjGkqdFKOrDXINWlV
INa/lhaNWfN6ppLwfL/zXhtQY6XqMjOhqOFyQmL+3IlXKjkTSf/OtrBMZgNh5kNm
FfxBtIGA4iO74NL+txvP5t4KiT9OAYqEQvyUKP51tkTICpHbyAGCzS3YDBOKwaVf
wzED+Xv/6OGynwmHF9xl337ehGFPMcfnYbEZiFetrmicBADpIxt78OhEfnWB7TbP
UubMpgzZX/2+S8s0UE7P3vAUPcJnCiJnSQK08L7OK4uXeBoArS5v6f8J61Ok5wxq
3tls6CQe4lWrXIcJHXhTnV2MOKxopdfAXsoYkBHS2aIX7hL3tS3sT8lBfowdO9G9
dKyLgze5AFMCR+NvMYQiCCw3MVsBFW0rI0w5t7M9g5HK3scVzSSJrJGE+I2WoRj0
cYXRQLPzHXmWrVqyrleWxEiIPFojWiCDGTtE/LA44jBrMdeKrYcYStVNFmFE8M2V
PqzqQ/6AYBV38zHH+uyHjVD71oD6hGp8kCJ+WyPRpH3G+ihLMVLaeew/2q8cUH//
xOfvtxZQya+9Dq2t4/Xt9Ct85HaiOB/8787v/oxJGBdOpVMFjetLWwk+azWxPE/m
e9amy+J1xndZv1l1I/Q8S3ZRff1c1GTQZGiezkgflGxXCg/uc30ZEfE+XMoJLSNb
8yG/cjJZ/oJ/cdlLzBym+vsOTMIWidv6UDUZP5H131+bCYW9qkEYEfbJ8IhGcBLL
5mUZQ5kS4crnwp/5tn65JmF2Oci9foSvvtHuFg9/Qzxl05XY89cfXJtru5xmiu0P
jyIQO4C5Xh4xT9FGGNUScfsc++Wx5nMBX5N6mrD7jdosFz6DFZrjJHp21AKVGIMJ
ZvdMbV+4zOUIiwJwi0RnENprcdLUgm8XJyqUK+vbhxx6Pdgf9MhBVk81ONtR/uD8
My/B2r/Xf6EvEAm7qb6+ECH7j/VmCeUTNYCBZSODqPOU/zKtzdH9eFarNiC8pIkK
XG4uwIpyPPSe0hiwHQeTl5U0Lk+9HqySp86Gze+IqxTO4JGWKtO2lq77vX+joBx/
OWd3N+WYhCCteQGN2uBTvDXgsHBFZALvuE/VNUQYaRdYd216VSZqsAMcmfKimUvy
u3iE/O5CQ5nK5MGurA77lbZU9Of+Z5+URXZ7olEEwWdoeOmKZOeYLg2Ce1QAHMTF
PDR8bXp2z2yJKUTnSHXV5+779QDdq7XI9fnmW2WTAYV/RYXarTvHGQ2og4QqXoiH
6mUVfjv/ETWnUm/+l+9lEeDVhrRUNP6Yllf4waTEMYYaY+fuQ889m7vHn75PVB7n
0JEWomHja9LIwd60y4ujUuNkrdy/D9Dnsdi1/fVDiHvhz2pndzTQ1YdIrUyfr4hE
mMZx9cPzFq79yQIKpD1WmaR+Bv5OlW91lzA3wOCi+jrHnOE0Ri52YjEEmwcfQ8W1
n/JAhQYU4r92gHeTyL56rSkC8pzhb3iETCPz5bS6TN2nq4pOgBEv8yAQnRltbxG0
BkT9raZQLdOpP94c29VAaWlRxVvSxlE/WDof3F1zasFbKqLb+qutr+MC5RzyueTp
+KsW0iUxB3lGXrad7G50ksYnXeo7P6r1suCY/F42O9F/o10XtOAD2mEuZJyLZnnB
IN80tucaG2o6h1g+OW11xqzdKZcybUonkps/D0+dn/aoDiBG8Nzq++n3RHA6kKDi
BWry9S7yyW43enKAF/EGOVIYJDvRip2R8osY0J10FBf3j+bU8a6pxcKTQeRCH8Gz
TLfbCwbv//uu7LTqRnnR4BLuLSzXjMbcScSM+gSESExSZaWtkDK1IwerO1q61RWt
NJRPKzBrZ+h8wis8onOuExtbctqRAndrjeR+4soVaP94ay7FxxSrx2q+gwmVUn6f
xy3dsYQatp4/+HsL33YCPaQeW1Dc2C64dhVi/bsGwUVzY5A/8OWgzVMFCjHhjpAd
ulO4Pa8/MrYwZyjLTxiBuw0P3TBXO6lmNz/MfIzHooXFkV61lbrbKkEYDz/gZmfx
WJvI8OW8xPR1t9+UJuEHm2OILmSCkoP9TviOKT+6NB+bTNfpaFoJ7DIvQJi7tUqm
C3NTXxA3zkUdQ2cf4NCtw5/K7oi4sJYb1PCwrhrSzQjBUmCBDQYdYQqYz21GJ9pL
0rircjY1JhD0CWzfx0ip2NLPWkMv9C8U54FznuZgsmv3FFv4MBb9nU6CPDH1errq
jPXjjlrP8Upl5FawQxRTWuAmg19zPHIaVtUQUgF6fOngA62s/Icv3j85o3KrwLim
cwwOEDzTZcHR0vDLppqQLBDmWoFN6L9HOBJKa7tUdqVB+cCsputpzkKaTNz/hIfW
RnOTux8gpZDuHxTb+1PTw5kcCZB18+bz0KDcz0Clh9qFADyEqMjXX/qEJNnNzTZ7
gNeC4KJptuLfD/TyPPJ0GJx724NJZ/xzIZtj1pMbWlS3TzEbPBJrvNNFWmfy1ahW
sOc76y6Ck+rF40RXZ8gE4CoyLfpleGrFDCiT3JCZ3QW7/mV9RJw+XVPbABn4coEF
E08obRdJFVyFoOJP+HEPtsPcBzyOaXW73CNztvakmyps1gqmds8xnecWCI5tsFEn
FFuauKm1LiVwrgmHJJmIvFjqlKaMUC/Gt4862TAenSFrcZYGYu48JawVktAoQSpZ
8P/1g+2J9vlnz5WdCxZtk6O4D/VM5eN2xN8fPQDsAdHjwEMZ9ebwK8RHSfp+XK3n
Bo5CYloPK8lKEq3D5tQ9t+3CMABh+aWWjBJbx5489FwY1RVKCPC8ZNeQe/nZfddm
Ll1eZI+zki/d33gsDEduGXPgUgvDVN4u0hD+wrqbKC4FXacq+ES+SuhglK1JWRav
tmfhxs1QNK5nB0wc51iMo/LgejhoxGq3LQF/ghtYVCC8ABAieJQRzhZef2LD4ouD
mMBo/0+tJx1cAuqKvz7jzxky7TqubqEdqVixdR8k+++6s2cwjdof5wOixNa+Y61s
a9hpY5SStT4rVoD5Mfj2Q+3JsMJ1V+f1sXqY3xxiOygKiqaV27EmY4a7bYyLnnJq
l2smOFPzrRQop2p7mu5ubVRvtRrHi7LJW+OQ3n/JqUYV1nSt7E75BiuNOvcIIhWZ
Iv2UFZYX/si1KwiLs8zx5DD9yoS6BQDn4ml99on2FzHxSq6ezG09Kv+GzkCqEPaW
7Ke9BUIT7a2cfQCvsokTmCNs8tT+7Qb2wec5Ifwif8B3Bg2ET/F6SSqssSrvfdQT
WZcPDpU1KNvi49h0WIQx/13SDWxqsgnkf/3jxRN1TLOQciTBcLcVeFmFO0gWI4eg
1W/BGB645rp+ACBThzGQG3RiFSJcI/f8+RxJVoYt56zG6lu1m1UNPfUTczg30xyx
4xfROxabjt6iUV6E5SYF8atLd1+5KATWePw4Z9BpabRN1UR1D0YVUyykqby1AJxx
Xr0tj0sFOuY2+3BCWH3sUcA+ssdzFjMRQjlGPqB3ht2fpadB0UrzR343VUFZPAwE
n4mnWIR3fAmV4V4ylzz1FFX4jJCYJySApyUtAQxpRwNaRpnPWa1mUT1/Wl/FCZxk
uEz3aszm176vdkGxnWoyODYWehh5ki36WY+I92Hpn32PZV7RcRtQMTSY88Yan78e
EUMEwlPPxyQ7sfwiFE1lC9zK7IPBBPPsFi083YtlCk7TQ9PuRpCFU/5823xN0ujt
olvjCVYDs1FIBmYCHLlktH+oIEJ3T41OoT1xj51rwioyNg+ZgOUQmrA2Zv03+2Ut
WxPj6ki+wMGpsaUyne4Lcrg52qG3PbFJApDNxW0PyNWj4zM2oafHIkzZGDu1u0IC
ilWb0IC4t7qlKknzPlgChwruO3i1OAOCep0Nm2My9p4Qf/+d6suNTnwCFsg3Jr7C
A4Y/NKSgJSmEuDd04rS37UJXtytlBAMi4vtKnAk6wNKOZpTYMfNHiD+NvoDSjIgC
eRqFB0a/rwro7tmH77SOgvFJUPropdx3ZgYZfEBg+VZ2bXZ/7IJ+5u8ux6KbOY/Z
WdqAalki+uqYdPzQ7QbNGHI4LNuPORv/rQWK4Sk/wYk7vGGiok3TVnOx8SdbotqX
8nLnwYyfq26frE5CRcCe0Ajs/Qa7KUM54DQkxYITosXSHckZlgc734WGGs14Zf3W
PH675Frc8ebmS+kTFCnLF9NsKkrApXACYR14FAe6eiVSBO5/8sGg26Fcqryg+vnV
2h+bxrxTKhW49AvJjfcKNof9a3ESWcfeWLZ2wjA9aOLEGvhtBKD6u9J8HVktoqPs
fmMi6sbLpsUotpTDrL7i1ICf3pDbzodbhFG5WEmmpL9atEYAgdUGKfkk2aT2SXhX
4lYRHBC6TUAItmxPThZJRmyclCfHPNUV9OG0BnzhAEdTgUKYbp7rimNvDCiZvdLn
RIG4k6lP7PjOyBqMEjhocoshh2myc/QCV5e5JqPdHuBBe3qIg/8qKdlkk4FXbLeh
9BdvULdPho3MgLUno2P0kf8MsQsNBx+ys30GkG5JZaqw+OF+kb/+JFEkwc5A8VcH
v2VKx3llV8A+jWQym4p8Mz3Dt9AbxPepZvmWocPIr0gA43RrRXy9CVps27yj3V3u
MIiCp84Wpehku7Tifr1TutPxBMdpTtBMUcx+jiWjV/0NmDLljzBcbC+f19D6s7Pu
QxBzAinVA05IivqaVjEp8FKty7aqte/IwTDHy1EJm+XkGitDVDq4Omn6EU/dKYO+
PAJodMvyDK6JlDUa/n5NjUmtafBEsNi7DyKEfFgFKEBA3sJLSxCX9DtV8gTeBLYL
g/NS/j2vqzU+oaR++w9vrPScytORI+B+Vy9TlevYOAHV8ZjlFaufcDNdWJVW4KLs
RTGP9f+3ZorzlY2PLz4OujjjTcdko3y0QKOkCjfDRXiKuuzxI7cz2NJaSHo+3kje
fgrdyf0cTRFwQ69I/iluC0mi+wttRBqNIjOEiPN50KJ2hKs75jXi+k1FPpOgw0EH
7ZjV+VnxH09YegmaIkbHArQTV0ZUYfhkW8pf4sf6wOj4OFQchSy3UNGqncB3ROLN
NvA4zYlUc7byOfbh1j9UCLVCgZe07HAfOhx14IkIAU9NkbJ7rzGUwP+vS/QMgnQT
eraHSj068qKUrImPRxydcW+F1B6a9CpSCpRdtpGF+N9Pdkg3FXui5HkMexMAeiFv
Dc+NCckOwkZWIGwdkHZiBEp7zE0L+OW5uPwIQSAApZy2cEtXsJ4gLdyoJQJgAqN3
yhq16fxVTKfJWbXtaYV48SOVXLMhzMLMEYPDPqpZqWYNGVb/WWcgc9kLZxLW2h/u
Gj6TLTwie1ILNzMOhFC588hEN0VygAMuuaL2QLap3lP9kMrilDL/Ndm3rqtCbK2c
WEs37WhWnT5f17J1iRb5/xzYBaGgqYvmhGt0FTlptkGSFnnyw2Y8D1XdEJ3cCmMI
I6OcpFnrD9EIBwp4Et9jDuPdntArZ1Rzo5iId2TY5SoBhIB8v0XU1ISluHvC5VR2
3Qg+3eNRdDj7o69R5s1q5kcc0/3XtTYbe6b5DpgXB9LUXZzUEKao5Q2go73QjHZ4
tuQmIBtTfcN5vth5dlu1g7Kuk94u5rY+bAgAXG8NZtJRFMvBJHesS5tuzEgmx9FS
TUf5TU/nwEEPg+6NAbQ39N5bW9jmMxhGSEWjjzY/1m4K4qe36x8VxKAaJe+xgs2/
nK1zdjINZ75zfnkHAgTAfkgIDF+Wwdy2QGCpBAx0wLDLBKXRLTWPh1UaYatHHIEI
CL2PSloAaUV8OwZz67t4bH6pkDpHGCriAKbCTfHOujECA71u14fKOc5FpIbe5oRM
flpZtzXalrdXmk0r//5vBqtS0asEmCrGwXM8moemUMjimMNvskfw8J5/JvRUoVP5
JAIqsThYvKuLZIkKRHp0RhD4oFnoKf0U7aa2ApN0uGNv81MXxcyDkxYaAnIpKYaY
P766GB3Wu75ip04jgmP5tZKVz4guTQNZLt0GrxU/5Fkyz+M2KZGqwanJRpZm8SAA
PAT6JG+qawXUy6tJwmg9EariE5fM4q2zd+IR3IXBTX9oUZXF6LTtT1hrosiSWzlA
5DP9pnTMeENqTV46yjDWyyAKJLK8k54wQVk86v+zmEhVx5pe1ZCQ584ezJ/0X4sM
ipkXbR0bsOzCG+56OTOmhG3QxSAq8WrKsyFe8TXbVSGgoYreTZK0NpUgxyB/QJ1n
C6b5QYY9nd3jgMGDBSMdMpE2fBbrcoLkEgmjQoWsScwdefevRm7AoKyZZwrjX7WO
Fo/6hu9qx8LL5mnPGRJto+3hAb1c0/SGSvv5j4Ys381A8HMfq819riMQvmjDilBi
w6C1Xp7HeFoMd9MmkgGfpaxnJSLz6pgKQCzmGSo761gNvZVeyvqhHm3fl9gj2TWB
GLN8DjprltCi2RnekPkWKWH1jLghcT/DxhZbfImKUiH1Sk7oRMowwy3h8Fi/fnyy
/8NkeFlXRKPrq572uAJCbyjKZN5fRPWMhd4UVG61QRTRoAzEB9znBIqvKsSVmVdE
IHdEtaYQJas6YbdxRGP/00BtqvVcj6M3HRQj2NfFIFhzUcmMjiq7d2hM8d0Imz1g
dPgQ993kva50SS3ytrVQSBROI+c/5RtBsTXgQTPMDadsMV+r/vNR7yCA4W7JtDOi
GtvHjb8KY5oLyKPMPoR6mAUCzaXSO0t0hXCiHNrEXvojU2I9jy8s8d7RWX4qo4zg
3v+kl88fYjPiZ9dwYlZwQJpymEI7u6Mn4XSzg8VSH+S8arlz4XcFPBNjzoq4hW7n
gTY7HyKWxY8qbM0XHoQ6EXQ1+4D4YH6BLY5nQbf+yTyDsSwaDizlHUN2JVnGZ2io
otC76QZXhdbo7GBx/IdJorPsQw46tUjOJ4lQe5SPyJ3HX+8NGqYArdJOGbnRmJJr
RupBZHooHdEiL9VO3SzjUEmccVSM4j5fZ5xyemLkj29TfvxiXigXU6vxMBFMfmUE
xkMzjd1ft+B1aQ4SoW5fU0LWNCxYjaYIbHmZO0Qe3v0l+jlEgPKXkywRRczzlHoa
g48tcIOCaUTN5yY8Kr76n/0WBN2jq6VkFbT2TABwad5s/QqNGbm+cnpgipZvbBKc
ndr9Az0RP4eCBTFwpdRiz2IavKNdtM7GNJ21lXhlJVcokCBbK8d8GdDxVkDfuR8I
bJO9YOReC26fS9Vc6E4oUMj1xpAOUzmcwTwHGBwKbr5AO1gveVncUi0P/XsULrbp
TD7Ki9Rd96bj6hFZz/rmc7w/yQLhskApXmYhGyDqsyr6pcRcsHaIJKFXkfpjY74+
mf3dQ1wrDIp8BVqIWm+wCZKi2Nnfx1GyTU39poJZnGRU0ECVdx7RgCaENu2jkjuC
GdYFjm1pajbxq1Zk4JhJ/16/osSZurE4/Heba9GTIcOHEJ9XLCJv1Ixb59irPj0h
A5SJ/TWPyOS8NPp8kzU36EGUCO/YmxfU/llf9uutK6PuMklF0zlZz3UEmx8DuY2V
gQ9LShKRpoRJWRHUxystWF7n8IEvpOfvwzaYAkipngUqCCsEtcs5KwqYM2H3nCX5
KPOvB3AIw/crra5ccQsrBvVTB2vDvl6vqvVLrFF6xK5P+w1ta2WSdIe4w6M6jI/U
TcAJCY439aB1+KWoqMAWrhZ+t1t068O2jUrb3O2PtZNYLksJt9gz7PT6/3Pd/JDs
TqIbx0LaP5Vcu4fJx+HumJgZ4zr9Dczxd5WKhofsYi7k/yOYFQ2Hb8V3c+zUxE0n
WyHJwE6UpXv1id5aVe9jbCb4ymTDB3tc1srRVM5Tlh7QgHdp2RIACu3s8nFM3zoX
S0qC92c/RD/nQcSvUBXUyMIa/uq3m1AoyyvpD3XK4/IiT9NQ7RQTTXKj6YNhMs8j
BoX/NB+79CtAo+3AlfDm6Gc8sduib2UqcBE2aMTgRcaUqE8+/JjfNKg/CzoxM443
lmcD9DU/rSPRj0Y3zu//awsSCP5GnVmdUSojAN/3PFOwXfuJsdhPFmygEylRwaEy
a+ctLwHf2dZOjVt2wPqXan3KjSJFtQbrW6B/ZVo8yj0ii8y9JbHF3wJqyzgBaUN/
kvO15QN9mXMgkk547XmGK0jfrIPHqhOk0qs0rN4t3g4RTq+sD7l7YjajAVl3CS3I
Rj0Q9D/Ok9VdKfEsjWaisuvVPDno7NSvl8mHIQUlIcfvHFU0X8Wsnm/b1+1P1NLP
w9OKIIMg240IaRC4sqCbkbgFw/LdL0TVfhdjAFUWEwNcpCExBr0Ip8Qunwyba9oE
b4++j9NmmshTQsN3SJMSOIc4q9sqQOTtUZ6bVaRI2sZEXhj9t9jXpT4gIjCqIQZD
DTHFwDaV4SD1FHtDJwuDC7ST5IaLOjaXENay0xFmxb8gN90jI3KheIBbgw0CALwu
Z2BFsFL4RvBnlKRfqUAUPel5oOE85S2XBoarezBhlnM7BZp22MKn6ExUMYpdy1uM
HJkPFqkz5cES9QE2X4a55G7FOyFrUmNbKiGZUjXXy/ajCrcdQ7ft88xhKcWUi7Yl
EU2jXmLMtOtvDTC1V+j4AT3Gp8gXr22Jo4gerQrE1wyqRwNhmWw8ccgQC0TNICAk
e+b+SOhILGfMv6uB5G86rASpdXFt+0yZSz7MR1AzJzXsLutwF4wbxn7HBZDFDQEm
rK2vMwk9yNqpIBGlFynoOdH4IGvSIgxIeoDt9wVaQvFLZYdXAf97ujazLmM2mEj/
7mwXTpSX+q0TewLAtxyuXbklEsR4DfTjLDffbtWvYh0MygMP6+QsacLrS56Vd568
ErsbedkIBLey/S/rSOUJ9QX0tnwXbZuQNSxUGOJR/4Vn3xY70AY0rPmUt5Ou7MbA
hjfE8LDX525phaM0R6Rc8Zb2AOd3tFZg0rjPRK01y/2PxykejXaZ3jr5K03Fqjrs
4AD52VbJJay4w1UxZpukqPFBnobA7ZUPXb3/AomHFxKKiaAUDYaYkNYSc0NTMtzr
njTfruPiK12DcG2JoMBkucO1dBiIhlPPqgnOezC0D2nXLS6FAmtOSNPvN7x4Vnpo
cdwAmPtW5OG+IJWlJoQkB8eT991vQFxkpk443AK/OsiENQbdiKsBiE6rmR5tbFAx
0YWbnERwYQaDa+S0jyUlRgckdV7PUKdBx3MuzvRQpvaGPvtpwK43Gx/FC3cYgTGa
s5hT8Q+mVnPBthNnS3RwSh9sSbQqXpfHDppTFNnHCJ577Lfqx23XahJxYb/+dOIf
OJdqqgstcmqcqJVKQurvHFieTEs1G7sljQf/DioPxSa/Bbkj2RIQlpleGCcpnMLH
PxJkRHntj983bcF1xkRfVIotO+XLEjy8YqNSygyY0hSkkJ1MkHkIFpl04MAuxAP4
vv4U5yUpO4y6PwYjz4/2pXoslDh0ZGyJ6eAkgnAt5agmyXvx6hgrmEzBIfBjEcEC
IG6Gw1lDMQBMZ/wRqvTlPRjevCdJoBk4SaUGucnsD7Ysoi39gUt2UxEX34z5W3K/
ZBLkaTVQXUM89grsWWNj4jxfwThIkf2CW+2IirHWTc/gQo1OQ0x2l9LUxTuRqxb5
XmLnigjQaLIMLp/H5pU9agO4E6zqnmIMsy0AuoGaytRUBqK7hroUB8XJDlIlq3Xv
g0ycvfEpvtPl6hnQ2meDLnPcGxL7ldq4AJwXjqRc2d0YVFIrRu0pKSdGDpbFLI/N
krTV+VjoRjZmrMho4NcoIhJXbQpstLq3zBkr/UxAdwceNkJEmtfvxNvPZ8x9i8yC
iF5xXylP9ASVG94P46kMOTMyz8+CrdE7f9dTiT7DbeNaZbAw3M02ddMR4KsGdino
ugEk43iC1WacEfs0mnI7/1m3Z4wOr3/Du+l0yiXfMd8U8htrhF5Z3AldZOFarJM+
dwKGNDP1wGwc9Sc3h/Yn/4fNZpKBq06mfs9wclvbeCNbFkYcdNbnTWdByhAc51bp
KJwiN6QJxqIrNLsOduH6QUCdpzy3+Npu8cl7ICA6G20TxAK0aJ3bD7WS+/un3Fyt
Ui5qbdxvNzKPPQu8SK03Zb4Accx0dWRRsemsxNkTBgzVgWuMBm/hzfhUaeMkkfyJ
XVm6Z9k/TplvK2wieYyD3Tp5eATRinjWYaPL9TcSgYId1lsUUSIpvK7b/YIwBq8W
/tMI2gI52colFfhm1rgJ1i/HhpDxTcmgEe/Vh+CLwNDoA8lfsUoPkNKdOIWHI2rw
LWacP/yeTRKpK2RM8uiZyMHc2o4bhh8Wu8e+cE3TgrujrbXVTw502MhZW23vva2j
wJkUJGCLMQ68LUzX7OCIJa40usB5BpWjaAR+EM85KuDrRrf0x7kdBJMhI8gEe6kN
xosbwQDeqAB0jB5sr2d2GfFOO94pc2dnK5rhZWHVM84jzb1EA7bmB4JdFYrSpCnP
EZBLlEyiuhsaqPDXBanKd6ES7lCQd2FNQBpzSmb7buyRzr4cUbhdBWUTobYO2W2/
tcmMmVHdhE15+Q1qTRo/DxC3pGmwu4wTjsnCFAXbmuZcQZaAFQkYHsuYX2TMvueo
5yulsVM+85bDGEXW3LRDxOHf3Rgygp3yL4pzhFA0OsS75cqEoPqWzTM1Y/wucSdm
DXnYQnEbL55qlps43OazMkpXpPGsDrySXlX1yf44W3iM2cS8DzXvTpTbWy3orPft
IcOvl6UtfkwjUk9uuLr6IPlzAKkDuPUu9FSgfVbBZIh0UyTBOaSYafi64h/mZOyc
kUSP5DN+0hKcur5GHJbIHU4RqQUm2QBxEp5c6iR75P6mp2DX593IquE6DtBm+1sw
e9UOSUBm5cA9SOGkVqHwmW2jMZ9p0ZqLrkOQHpbeF1nG8AsZ4T9o9l6t4dk7idpg
k7RfzjzKy0bPKnvyiVTVQnUc1b4EKYSkdrQhDlqKir+ARxQX5l/YHclDVzAFM50Z
FRriumprUDJ4Q/4w4H92TBIeNkZRmdtNLIV8Hd7YjuF+KGIgzFi0ewpgAyXBAhJ2
PF3+T83jWhMzE/tp328J4AsQ8CNEXYZBMVs/4ntaXbYFI2cfxi4Ca/ihe0/uHfN9
AQYFzLq8P+NwExq/nqTma2VyFBFcpmlUAbyYrqyvfy+yvT1bhHm1fHazfvCzodrf
k2fzcYvykCfbAb1KLocAjYtk9cJqUE6RU1SX0gf/pATiBkk/RDsEKQPyM6PWjYNL
kLSgavPOjmNqsLafSNOikl/o8EukrfqPPN3yaY9iWQnkQoxzAtzt9rv9MRdrCTHt
CZtYlukvSA7wTUkmIu7ULJ2fhhLwPpJhQtveiC0TX0az6WdEYGiso2syWzfARRlG
GnVU5rxioqMNJN/Ge8mI5NYDP84y0UEVPmzdH0N+EcGdVl3WdNV0sUa/YKxGiAwN
2ocfMQ3Ks9SiAZjWxQ8xUAKTDU/GXpTKUstFvVLBW+QSMeZ3M1OA6lZBKOKRXW8m
yj0+VsPVDEcjSgZPbscAdPEABbKg+drd0TsZxuh1UsBZM72M47BKZT5XDLMHNufz
TnvwFhZIOAjXgUaC5h0tjqH0Ha5ojIkwiv4fobFlyVIPHK3CYe9vMaI6jYDtP+8l
74TOklKsbq/5Z/XblvhC3Rd0DdVB4FzuOOb/UUHIyLpYPKpqZ2RcxSKPsXsj9vvn
aKsZs3X7M4tIUnxFtzZJ4DCTWLANnCLdIUliC8l2mNSf8g+fxj1h9f7mzKDLelaG
rg1Ee+Df6wbKevLwGbTjAsZv8S3GAdJlmzXI+rBv1qX0uYvanHZuPG2vcrpewgyR
ao8O33ca9X3XiP07eKs+9mJV2ZvuInRA5F9dXlZRcDl3yKyFIBbP4c1ex5SDyD8f
DXt9dF/szOZl8GiTcn552l4bULn1Hi2ZBeqLx4tcUnCJ1SoxZIQPfs/17EHfZwnD
bdjnJRCa2yFSQOsxi6TNPHFSoOXNiJgOVEYBgAonfxv0eVhVpn6/3Q4gJzh9kNxP
43usTkO65yxP8ALbgzvD894/GY+mNA0JFIUMnOHDRcJcpwaU5MKj6kR3K5V0/LCW
j453oDQJB9l2EcWnw+kK8PIPw7qXnR86P/xPEdukiBWUWfAShN0qM5bhKRmSDwrH
y0ehIUMvLxaN5dcSUTuAaP/pOsQHDb5ivqnpMP1RLUUnA3DXN+h2EzcWvw+DfKca
fXtF41CuIrZw2XLw2R+UBJ+CKDE2X7S3HXCSQl3ILwnqT6IflvzfbA6a2pnTLrRK
eREMC8UqmcR48jlyLbwGEenX10VUR5ohSxTlB4qQix9Qtcyi+VmO7+eGNoL1Nt1d
yn9DEye76Fx887V+/xbPcPv9nTBIoUQUZ1HV6THRaEcbdDiyYM0PvOsm9GD1UNKJ
405zT2C/ZkeozsSW2u4ystHcxY9wgvJhHqsCGrESZhiRjV9fEW9FBxjkzYggGblj
wwEGzJmwJ1dLCoBn7ooDfRRxLlFhPm2HTnuqs2ycpNh4MKdtrygSsqpqHtWo6hkt
9fCfDReRDBhVmkUU7jiZhw+y28AoL9TrtxnBPQi2tbFVtDLOxrJ9hg9cP3g/VmmI
+OrwDPj8s636QI4nh1LPJeAnvWm1qhltjhRk/uooahyabsTdoWYkIAKt9o7j3Yuf
PBLv9or6HVfDDxEAIyUK9lsHjXDbCFhne8oc2ywK2BPuX/vVHke+dbKOgu/5GPZE
VcdTm0mq7IdNnm1xWllLk143JoqwvVQVew//iV3zZbqIWsGM+SQS5ff1m3wcDcj7
2cLy4qRsoIMrJD0kM58eS0YO5hUi8LDZ1L/Bx1EsYEj9anQDAN3NJmStvWw0R6fG
pF0muDZTzeG2Umk2q51ysvXrMA76Jh4nEh5tWN9Nh+ute/OO8uXdATSXGi0g6R0b
J/fKVmZmFpmjFqB+8nuSWPLcnCuJdVd1vf9mu8ZlKIFYgcRsWw7H2MVOkPg0fDLq
k+aYD8SskEG3691AQnLo69kEg4yr5D/ffLjSzyxRhp+WRRvba4mz5DCuhCAuTFwk
VgtI8EBVB+Ysxe6KgaLAwfar/Ivr7bXbUSOOKhXTsReI1c32spfvO5I1mjkfGKcb
+c0PkBmuhXMKfYFuoECNcEHNoS5j2UF0iQF1Un7hxnrB1HDj15z0YmeATztoHQ3B
oXvRmI+McrQoyTljnaKN/TVNSM9ZABXPTId+JLhWI41ElnTzEJeLHBfhW0aFzlhF
FOkrGSiOot8h22V+W0xIwC5+YZ1Zu6Gbwbidt7cYroGjmHMJy6vFd6CqBtsh1hXa
mBe9XVyaizbrNeH39JFNCAJUn1sVkY9mQ+1KM1NGU0EIBlSx0GbsrfMxILIrL6Zw
t/aBTdKtdlnv0dD4kCC0bzzTa9oIPgWTZkFo28BfiiWCiSmi2JRSHmxxYUbVUFdE
oHHHE4Y4uS2J26wMr7b9FmbugHwifIE5ohfxbO6+0unRm+e0VrbNi5/t6D9XPhyV
aOt8BRU/nuNtuCLg8uOhJ4BMfN7H1wfPlnK4Nhh55WgiHVPcov0QYNQe2cU8OM6k
qs3pGK7+2vmUaDJzhAHQ1vOFsk8p27m4LNqw7oCWjawsQcEfJ7FuB/wQq+5XAWVt
1j/aW85btl9GAUVAiookQLf3jZzGPi/qMyd2yoTaGvIAKivSTdFOgcoJYSmVR99t
OzbF+9XgVQN+MD+79jXzCxUR1dlW/5foGhxKV2E+IfTNAiNq8FWG87vCzdN0Sv1U
sBxTxeJXDwo+99q0g4v9LOAwjG9nzPbvt/JxyDh9brrGtT7UR/6DvcJeySDazwJH
5oWBjkxbnDuA51BDv2K/6X0gQZDz22Uwhnl6mfSMF4ZiXnQzqe00F37ckj0/ZLRf
/e6/iYolNJ4CfuxiH6n28BPAnm1hTOKSDxjhLkK26wH8+1yc+rh6gYhPPj87faGz
7oozVGSfqo5c09coa5ydc9byg/snifIPmmGXzq1r6thPiM0EQECmLyvYFPCVxRfs
S5b3o5bXiPSF4VqYNhT04FIoWDIbfQNBp1tAGL1Ujj2fPI0ybFwiYeBhORkP2any
KsWeRvQuXnUG4TWYLEsGNUjkmtrNTEKOrWrw9xYNt9TY1V87IM+JOANJ8pLZbkgA
dZsAWUruxTDcHS7lMgmGvf3TlBL3PyY1nD02m2tY22MdtjYcx+HOD4r1QA2oDGoW
dEMQdCQ2GXZsCn3ZbsmocOzDLB4kvBnIVnpvTjrXue4L8ehbgxWplyyQk6MZ0DU8
zS9fYQ/VTN0cxTOyM+QZXaN7ZX/EWW3bDIGfSr5kneIbYKxMtoG2hWPYV1yMAjQS
D8jrqwR4TJNInx7HxnZTQgjTzU+ew6Ccm1Un9aESw6HsV0AROnQqfwniMM3zZpl7
zqoEtcsvwm5ZOSekQNbpVkygAqgNgaLb4Uou9eDcdFCCkGdFJHMHfOn1h4TalR+C
SHIhJCO5eLbcUoygfxAeec/o1uChMyDBogpL9eEYwcHNs5E2een03senUtYEjsT7
WT9mcYt/vGNrbColLYt3WwzZHJGNjbJDp4tAErF17A99dYa3O6q90F3thCabfOaQ
pSrLcu79lsukIrVvOPcYsMWeaHsGFLrTtTJhn41O0gzvsWJqIdhTKIZTg3e63eBw
3BTwvvCGvYInGEqo6Ow+pxHazwd3Ifi5Y0KcMjDv13y9IoxuqMJ38wOBM05Z3FfT
+q7hE6nyvRi9to9mzg0QbxFSr4Mmbyz2+hQh+in/x9TaUdD+Zu1iugwHY2UNMFcw
tlLN5CSiY5XAVXwIUQn6uuYO7b+FN6RbfQgfXl5MHb9ImsTN9yF5owLh5Q2e1Tsf
ExiAID9tstCItyKRIrTvojKk/TbzKNrLmyMeX5BQptJJPQgwSWyV+9MUWbTEVfAk
2JelljYcgtGcSOBkOsSpErYruQFiX1CVEJVicRtFW0yJA1WsYcvIx7xUX0nboIcU
yL8lVLEUk4QjI+on/YOtKs+o8Wvva2B+87q0WyleaoSmJESs/BFZtdnZl6q7JdvR
ryDr0deiAn/VNPv4UNlXFO7WoKzDWZhCgkLPPoSSWezaFhS7QC5J4UmkpMxNSrLo
VQvElJA+NSYv3NYoBzr7+395IpZG4W+/yukyE/nY9j4ATyf7OSyErDzs8GTSDrIO
kZfRMlebRtNHtR72QsJCFOylxfyJM441VXIbhl0ejh832iiHwJfELEtFq5RXNKvo
6JDIbJfFnMrrV8ZjUfqV+hQ4feAgBij1seXy63RARdwIH3hsaoAB1oq351nEjbL4
h4+C8ZwE9aIIp4cYak0GTPtcvscsfvlGjEGLZH5B7kJhdFA+LRukKmo+5ABF1nHv
HDAgbKhR32mw7WXcQPhAcCRSp1Cw/OgoUwvjexJEyyqyfAS//W8+6apAPRZJasVU
WObvWtM4HmSoXJI87A6/M3OpR61U2Bfapv99CiQpdCIb0DiA48x8ZwGgiRVBYXIR
+9XSHJWdCecLoqRaFT8RsfVrONEEU3NCGWNebMAsN+vS/RVSRpanhoCTIFIosd2H
JjQhBV/w1PjV1cMF6qcbcWJEbIwurjkObVakaOzKhfsH0oIEOPdukDUyR/FAnlTP
I8egUtvYVYiF3zpnvTYg4X7J5HpwXTmH31eBcrlKE4rRH7Di17m7SnV03CUWGiHq
o4mmho3cGZLU3Wc+XsO9+zzz6+K2fXvU5GWZMbDeiHJld/UbzicKzZOE7wy4qNSh
4mnKJ6W4b3HtUu0IKP/4RQuypEIkbFfjy786NH8GzBFHBCoxKlE8L8xFqs3+D1Ky
u/T66494044fIRiuNFzLwImnQncSP3jZHkfRE5XFD/AGgtXloWx13R74jmqZoaLH
faU/BzKn3v9sdTFZ/ksVoAYNg6gZHMCaAR4vFKLC5bFKJ3nxHOyrJ3pWDCokE5FR
m9Zi9YqzPt5FxACrplTScbdaO6Rt38TK/r/Vo/itT39sveDbv3VrabKbauJLUDE1
Eo5emQdhS5GP4YuCII3eK1k8H1pouzkn12oG5o08x8seLORL+PCscqPfL2QjPzyC
9vGkpmS0iIOR7GqUBWoJm/Dhm+MQlQduk0jdk+kmSWxSevCni+fBbtWX5dGhMIXa
xKCpqMNmaFWgAXPA/S/3fPAGZOZYYdSwel7T6/JdwDEECs/hN8PcXhmrethsO+zy
8QCHy5AkqAtbgcwtVZyRM5qCM6zP4DBwpI+WmrwOT6HkI4ZDhpFCd3xX1rigEDPk
HxZhYuP2kgrH4evDYdD/ApgZHq4ZaaOlx6mAqNA3S2P4ptB2IMv+hoFuuoBDW/8I
YeUbMCzEJNKiF7kUbZpshUHOmZoSJKUL9ng6GNgnQsa3wpe/NKc5gJQa0+EdRCtH
dTU9jJfg+U5RZoShHiQpHt0XFYftdV2BKxXTEHCmo9WmjAWiL+cmEqpaVE6dsdFo
KOUZdfpCfZ2wfOse80bqjkGVhk1l+5ckfAsmtUP4+Fu0bEi7gP3eJgXNKjz2kbb9
R+KjeUFKipk2dAZb9huiELf4mT9rauLynOFaAAfSe3u2B6oyLUC0Fr8YuaV4DrO6
et8I6Jqf/mSAYDu08lEzSeR1+ST6e1jOD1TG2hVMPTDd9kJcdhBRSgcG19/DZyDg
g7Z4a9yCKCZpzMEQ1Qujbwj++EgH1wExMes5OSh4E6oW46+QOeuVIwfJI1c+L1qZ
ak21aknstvyyieJwD367HDdHOxBrZSko5LLoBmgNa3VLIF80wp+QbONZybpwrP1g
mv1kuSz2J8mQbV/NB6pmo+t5vX60tAz2IcehuvxZs+SrDt9l2C/ffaHXrT5NqW+p
UMGxzvq6jk4/k94zphD3UMQG88ml9W/4iGihBQyBk2AJkxukSSJUslbgjyTNKwGs
BYak+0Gvwjmremu+hpoTjEaHz2tR//lCCZUfIfDpjNvJXtpldnoY6jgEsmnV38wX
US+K/ANe4wX5Kuco3//ftlKmZ89mosT0iB8RdOkCwpWuKggBmXvSMUocCMW2lic3
2UVG/d5BPhCVzTmt/TKSIJSvuSmbkC1Y9bavRIx2dWPP2CYt3CbGro3vQDL17TQi
A7ywycINRFE1dHg5ZxvWzPnLpX8b4x06k5qaIbPcBE94sNTPd41YEBM1lvj43isu
lbuDcoiGWVRLYTrxPLfn5msOf7LTeHVgWPKlvQkn3Qz0+5JBePiqppgsOtg2NnBj
4P7U1y/h/+R9g362tW4ZcWnM57vRHSpPuPU/kLmuhn90UmRgSNppOyn9Tc8hQ3wK
kyVAEXxpbTwo9u/OR/xHK9oPTaJqa/Aibu6eo69ob79cs8jen7zp7Wf0PvQI9jpQ
zhPoX88hrvVqP2kmw2COj3Lfz0FHPxXbuM5SZmTq56YavJeDRYz0h5TTN88sHhuW
NF36ac69UK77snWESXQW8wk1xBrCk5vtZKIW7TjV+gfWiyq6CsCfmZ1NRkmxU2js
6tWnMSWMxGa42BhQb6br4RDkXLMi8iRkyCdJ6GFuFlucypErMkkwXwUC0/rs25mx
pa/55BF2J7Pm9zIGqUao/VPZ/HtoYLysd/LB920fY2a6JdOJsDuQis55y7WGURe6
NkosqaW2xjo7pm7RHQGU1CA0qqsPjUzvTPycpNNpWq0dZxnFqFVYSZfWRBvA7z2G
dI/U5EvC/TwTLsH44rlGX3X/z0hDo6qTWkfWg445cFHLGVd4YJeF/TpIzFC7nRMT
2x5BK1W0dIXsLKSJb7qc2/lNGAVu9VhMkHWQEwe8lIkNexTKZAwlZ9/x+nHs0LUT
ot4uPmOhcvq6kAAQqyCTpHNUkAgHy0nFPhDbBkeok4Vf+K6sXGIyrKnhLLV+AZMe
4UixzgN+TcxK+TzB2th6uHx2ObYwaIKmlRyOi6sO8WKC0Q4dj8U4BW2D6L3W9L8L
1UKDmeFOBcm7hEr/9haOdTr1QDJ/N4uCh3O7TJYqsT5SZCvLn90ANSUGBHnoShRa
HXtlNOwfzTrMwRxGvuFDeSQrRFleRCUau4nRMDbM1gkKd864tSizepXM0h4dfpxa
3e/wrXBAxrzCVKQfK+7f2qtioC9XBjDyAI4qjdFmhaUI6PD8Jr1Hq8iqeSwzs1Zl
eiZ3z1Chg+QdGFOJd1sTHKxjasqV/nkn1XxnBucgJD3pnJ2EgYnCmS4z+O9dKNJL
HyRq6XLD/l0lMam1bN0cmoLzlUXtVNBHzJzxH8kex7CZXtSPMEGYT6r1EmZrACON
HI4UwRsMXXHfd/Od2azWKVSWEKG4ZLAmgs0EPaJzyFKsmtql8UOvEB0xIolOFeQb
95Dp/OJR/Me1WzHpQK8BnPj8rTsL0hR1SkpPR3ME1y4i0PymGI7voaATyq0d3T75
ZqnUDjf4+AnTCEqg35WkS2vMHbF3TKmrshXaEUtHKty6MTN1WSjK3s6/55Rimbav
IxlwB4SSBhQzuxZHqJRC/aZRFzktqN4rATvHuhjyXFVx/4Tjf6Av0nrJ/EqZ1ap+
00vgT1N93QJOfDlKTwW0u+mLP2U1/Uy6aTQC75IA3+d6XlbYZ5NLOMcTp6ixyiZR
OBsRerCpg2f18IChztBdKGQpdqkrF+V1hqqdVKN+DqdAIJHISB3uvyPC01qqFw/z
15mSYC37t4e7avOTspqezLYhTKtXAtLISRLPDo5B4BBaLqHntrHd+LCKF4rve3Lt
JJVtrICW31+8b0EJnd3zXXRtXajPhqsscMbcgvH8kvdsYmK0zMgcOPFs8SRuDp/h
4i+TedxVIwM/s/61lcejB1/6cj6//BQ3AUlVYdFic3vw2/TB0fGn9tbJOwL8ejQ6
b31PllNahpu9IYaxhkQDAsIlu2Z2EsRgBUQvc83sd9moNyfB0x3BU9yrTvpShLD6
55wJSiZL55o7rzBXAOjOHuju0aiMXIasO51piiCwD3i8RCNjyc0Z6J7BuYgeHGdZ
dHVxEMGo7GXVWC7UyclSz2jMNLGopKcNmwFN2bv7dCqp9GHB9llu1dxH8XmKKH+8
y6wF99CekYqvYdTmL1AgYkgteQQdc8PwSqcexMXGtC+5KJT0cmjlzcMvqYSLE9Pd
BWe1GD2U5byyTnBpoyughU11J5DCU4sPlgG+eV//ijDkq6ucVdqOWKbb42Edzbe9
re7rpriPQ601VKXFFW91a4IXdzaMbnUmzvafUGgYuCm+Gadk6GK5UE3rBKqs0H5s
JsqsB3+T6LibtVOSIgvSJnBgjsq2+l8ODLOBWacn0MhLYygbFImTIuZh+Y03yQOR
2uk75jGAFIWT5AqqscnAuLpBNjlnF6X1g2rrSpPth4nxVgnkkbWF3OTlVR76kv2z
Y5yMlwVNUqkR/ZgNtdevKUrMuUd6vohaZMEuwkAybLCozzDQS2ORRK8OQmoocWR3
tFxnXEoc5FsEVVUVMcQCxfgRdOvWALuXpIy5Ie0coxW7OUhpplDFYrot0dy7N6GS
BDtoT0jEw2BUP+/G02IK0AHUXwls+H5CDZ8vQ6r9GyMbip8SGanhQcesOUpMRGJX
D4kvVF7eeBB1NUz4WBahSlY9Qn/KnQ+dp4MHpTG0TpNrBTKiEOy8uBYEzTH54Tt/
GzwSi4G8ICiXjmkMyWfX37XcUjwwoCksI8kKeIaN6OvV5oPI07ifbO6sTojlgkw8
r0zXab/ocJNpR30w1pDvbMZwUHrfIJyhNrpOcTL6ly0d2KRHalBKnzoSzGu0J8is
0m+LKsF5oREvtAOrnPTnTHkoavvznwIjFNrykyT8oa/8SDMuyxolZzswwqZw1bYw
sK4seG1VURsI6jbFImfTaYyWMhAqcVOJIJlW9b+2glsW3xqZ5Jn7c5MBLsgm5D5m
97QOH2VDYqFbZjon+O3N/3zh5M0oc0Gyc5L7TSJoUPWzFhavpRDlLrmqL5x4nCj1
7izxib/ZQ/iimkHY9I0q0Jx3IMoSYt+MS8KzBSgdwb6YDJHZ1Xvjyzw5ey+0gmiS
vJjaIksiR1U7hvfXqcIFHTzC7vJDk99ElfANa9cymflWFShPCsC50SFkvvfSV5Sd
2lygSW9sTGCOiNaABal2cpB0g5wRSLTe1ZiSPaqF40rHb+E9zIU7Vm0T4FhijArH
trJYeVNDUPxa+XVaUzsIHcd+4McFrFXTe01Jqdl1AhI56A/yqJalvw8X/FfdvPuL
xtdjBrnu95dImZqBJNW3Dw6Mt8tP5PGO7PgxoadN9ns0z3Jurv6PmQPQcw0RWnBV
EkR6gOqQjYUaZC7X5d2vTzePikoUt1RQONBImLHUKzuRuti4hpcafHbpY0CL99si
BJVDfjKf6hhK3z8jKQtMeF4Ti3YbU4Y2cfmEulB4mmcxYbZnDsOwvYSJSBeHg17B
F/5dSIE1tl0gtjA2Jn4Th5LeGxcE/obmPyi4zaCBGNiUJYfGJOms+nJgqaXYXR16
Utae1/P9ZjDBDYUSHLON/yDWDbf7kSR1ET6Nvmqi8WBeucfjjQhQq6JjIw7/ZuVA
GTBxzGiZbfdKUX7bwa1Wje9PWK9BQ9PQJHTbbStSdceBWeLfJeam2HSVyc0oGwQa
XaOGowOqWXhnbXtgRGysoYTTuwiEbGETapsCjMe4hvDLYtKWX4f3yS3+LkIgC9a2
ggPA3Vi09MHdSxLbtGgbZDyxz+iQDa/EnUGJCNhYYEXiVuYJkbmyGWoul3x+CrAs
07Ah567FGStKEe3xpJuLIu09H6urcKN+z+pDpcQiFyAlkZkb4imWGnKBgdaRS4Bc
rOPDluksOOEm2LJWPUnxk2Ih/Ry1jv673sm/Ej4pmmnBZuURcyuo2s0HdXJVq9z8
YyB4gzyEyyhTd0ZBs1C5aeBEVee1Z8tCphjaGVBAit6W9AUYmccfFFJUB2GOv+G7
/51w2BW6JIAdHENdwkfi1b3krM+ncwOm3Lcxeq39aX9fiT7O9NZTbdKmSIfeff8y
mEfE7K1A/0Zz99PxG/mw5MgThHmDEnRzbl1pB1IYR0YyoRYO2TE9AHgCIIglg0n4
TBLw+6Bx4g4XNQjnDmngIdOm4xf3sDXUIu5ZGbZ994kel4u0MCSz5h+wFKu9MusY
HBHOlF26y/TvmqRzQpYvdURc6YAF9+q2oXIeaLzLZ4EI0AGoq1vy5PGasCbwCuzo
eP2t7+mr7G/6i5LsR+hAKW10h6nL4VP579RD9ZHlhAIwSvogL3EMAyQZiI2e/Ge/
P+2bvuSu8yHDffX8ETt24q+xpocyAUPTjL3rNmG0sCL6KLneVzrBBl6wwNmLrzcQ
CgR/7bMK652CtNjKUNQcE1Hq/wDmfgbtwl7NNP+EQGGgp4sHkLjPAyjdbsjEOSxg
FwGZBr54rnYpjPr1BSDvf0yGC/hg2l7AeXp12UPQvDFlEu5zrjX84WXM6/isgsQI
E7v4tTRQvlU0Ngub/wbsgbGfM5jyTE9YLYngv6Zhjup3smlP1Sp1g6BrxvOjEPJq
YVoQeuIgVsSQ5rjqsuR/Al+v/hYpimf1/JPcvCOR2+K08Bvs4jCNCokdJIqIu/61
SLKFEz/RCYqZv4cpeop5LQngK5+FgliTkn7f2rfLjCpYdsHwAfsCLczL0oJUx1FF
ez2qNgCOeZonMQRrT+1VpdRqcssydCs+HgdcxK/xia/ac/rdqOWuF8o5RmMNmnaJ
pIEtyb4gkEwL533BNcNfwzAYSAZAzQdOESMGOJXfmXa8V8JLtnhyaLFEljh5B8Et
J+JjoAeph5zZHjYHPvxj9tj0fs8BaYDz1S3b0V6pF+1DtDHX/LAgRzpQR9rD21cL
oZkIWxnCF9vYrmwmCkTbNPrrOZnegpU+byV5uZFRHc9Mz39uWS9kjk9Q9oBw2Xhb
B2AppDvRJLPGEW/fevLtojGCqzX3kNBZTf/ocX/fT3pfUcKnaOLacZ/MZ3bGtfp2
ntUdM6mf10306HYf1AZwzG9fCkIvBKzz3jLcELeg0qITcYlrv+x53nAxwd3YkV7t
MbOLFvr0i2YwL4xvGFMOe3dBQdqUEscZIlj7oe8cwqqbZUCAl/Vw/IosCN8BYk6/
SGrB7bQ0unSbm+lYn0o4V0kl21j+Hf45tsP6qe/1osQPxRujpvteapDeM8LqPkoL
T9r/xjbRC5OrxlPF03nENVOkpW1qexijCzGXYCBiXG8YN7mloKI/t1zCh8FpMAgi
Msk0R7zwBAcvov2dSCQlggPmrWOqIeuIM4BuGUJEg+K+UnMO/wjMf2VH9iA2rKrJ
QqhsCZO4zIOaFkSRK7s0R9RiVAy+5AuslXCBB9a26iVqu/ItRmtqMY1r4VQNdXBf
6+sRvFD/ObHCx7vY+59KC3N2e3Nzly1Ay+rce9PDn3KSTosU/0MCwK0OhZ8OfC1L
b/Kp0E3aTLJRyQKsNrfml4YiFjmiWvwCtBA+Cp6bOXy0E1N8eBEmVu8NHYLApOOg
dvWW5HjVGjxG+KDQcdWVslcYFjvfuyp74YgujZolMc1nRQx3SALk4aukFFlTLF7/
8grMU6S2M6EsbKxK9IeKpwjmdhlAbAk7JFmotUcBKJN/57k+BGITKXTnprqlX8sD
aFmI7YDNlqtf/tDbOCBR9H/uzeD3bA4upSNBTpqPHfUpMPVyJeUC2qrq0+CPZKll
8rpdz5ig4rg5pn6uilVeSCkBfKtTCSp+jKli6iaCXequrO0xhO9m1cHpNiEDGy6c
3wHFpu5aI5YAcLE5Djxz7nw4l/70JaJSFRjkySzPVFlzKnPwlrCuq/kCtCx48T/G
1EsaIVda/WMOlbHZ11SVoHZu3F0CySLeU3wpasexM9wGdFjEaWDm7af9vtr5o3jP
WZG+L48vrVNCNh5OWo2q3/Q9YMA0vipLtXtb1QJAfHG9XoWNJB6Y/0B0FogUh4Ou
UcRfhVuoSkjRwE+xMidvB9xXfFdqHWKgeYLv+0Hc58LwmF/hn3vYw2ewbhN0gzcm
wTraZKWx1RCBECbkQg+KtyJD178EAWoAtk1jBlE9ek29OiSpUlzjgcZPiLBjwdy6
4mJGlUnygO3E7lAZiI0Vo4U0WeAgPyV2IPvscHVMEVm1UTWy9Z/AMPlvxUB4uwKg
UFLqr+E5rw4riu7oZBSWcWSpL3xr+KI/t/w+Ydg8Jgyp/gDxL9ogSJbZndS89HoV
acV/RY+5vjADD3AqMtMyCfr0KXcKY3VIqdQMPod/joVpwIQoEa+aaotaye4Qgrbi
wKxpYcFFNTD6d1uHadLvNWVMzxaUznVoQZu6Mv6y54cxIxQbEboYavs1SLKqA85s
2wOIQzP37yg5JwIj2bFZba5SEdixFtbWEMK7yNd5bQRY6NnOFfqB28VnH2eYtbhr
S5SXMiRAjS7oVBznjgnO57U3yo2EB3dHMM4XM2PHgaFESjaVaoluN6c7k6agPXOR
U9V85ioYGSPFL4ukJlZCyjCEhJBr1yv3NinI4aYrHHUIw/vpg2Jyo48Hqyafm1nv
vW+bY38hJIgmgTPfFVFHSbn6X3aJRypbTNgbZUFyJhJdQEnz365Njxy3mnkcaLRY
DgGdJDrCgV82cPt6935agvehGjz8e/LCo+4UbzkRbzkC1ycS9xBQzYY3xUwOE+xh
a2aq81A3tvf2bXsRs0aAFoKFBfFwNiMQqr5/SHcT944=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:20 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mcKPnpo3TxJFdIrYIy0PgijWJW8G4wwVbeGG9KVByYNiObUhnyQxAwHDIAcVK+2w
XYQeXtRPecMMPrulzcaGPHXDW14tZfUALNQ/b4tHWKd84wdLjb94sjjIK4juNPGO
wieUMbPPg31TX/+Q5aaOAukQemWYvTePUJGSrzFXlR4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26192)
v0PEVsaG7Qyh76kV+u7VQ0JxI1Kw/zdvy7HUug5VBwEVuKGUPhneHwlCRzkBTtBV
PzNNVZ2j/vIFyfSgtnCUdrcrsolEVMQHDhNPUNCvsp6KwJ9L0KBXzJSTrv2zMvio
yUSTJZsd0rrTtzEbN4UiRswU0QmFmBdghLNNsqduAl9iwg1PbIDXd8z5YX9huzKB
GDzh7i3D6TMtBpP5N+dVtLvifKfwWErGw0Y1WrhabIlCh7YQh5OtED+ElzuYcOQU
WgTd5U2BLOgyO8kougFHN93Ucj91/q4SM/eaX4wUjFOYCn8EFOJWg0o8+frf0GRK
g19aREHMQJLoYZVtBXNJgo4YPRpwSWZg2RV6nJWl8pAdHkEbtOKPYVGHzWSGeh5v
qY01VoTAgJgqRr6JAK0StJOzXUcRrNmtM7V/eImDxe3h/QO5IicDtU5+FsQgMOz9
Mei9eGf9YC/pei4W9UATN9aPlW832XmHWaQo39R05r5HhAv6b6kh19j6ACJaHTDd
o7xgE/36+K3nWYLOjc7HP21F0yQv25b4d3Uu0bVFZo+4ttVlsm6zTKm8D0pWabH+
bMhq9LI0pglIx79CtCTbqhVWw3bPsb0F2ZadPPLi80tzVvQphGV/vpoLf5WhbopE
owQ8TttPT5jAdtXLLVtI0ML8I5w5pYswNrbwKdzmNpwD71Mwv7flf2gfIoA2qTQy
KhmpAC0Rl7CLjqoV6fiA7dgBuag2rizSKycPRRR0FywZzaCSPt1wNb6GQVoc9EAr
dXRhHEBSDC7By+iOz9DBrZTjN6rts0dRTjIPcsSIugEkymBXBdedmPRin7Zfp/5T
n9++T5cs1QWsp8tKt/MRehK4bp6KhqEnoHxYxX/oWGOh79R5jYGF0IVIspvadIx9
aXE1uyhhbOe47/uGwXrHbaDoBGGEV73ZWymrmkmAH6yXqGe/sx0WW5zHDIKRAmrv
9KCEOiPJ+1lRHWojQHCG4GeUJTvd6mbWvME4QGDo49j0/Z2Gi3AJPujwyleJvirL
wjqIQfZRnmEvoZqYs1S0RxI265MxsHWuZ10lptP9mIh8FlNerQLR2oH4xECZts4A
G32zts9SZmgVEKalDMpZAcH4S5DUDDOPd5+1FE8sfqpY0VWL0cfbsoKOMQCRvEiQ
IGI7mkR6sS2H5tGgrEi/BIPC98QFPi+YxhrzqaeYOAWXG8MP/iXZjA4DFP0/i3Ux
NWZvLDH6aHGaAEFBUsJCIPD9DA4yYw5CYkd4okbYo2eFSK5pchSa7tpVvTZI14cr
mQTvpRDRRQUrbLmhDD/s9Nwk8+2QiKqwjKL0ujG1gQA/V5ICsVVKqMiZpOUSSbGG
QbcEg9pQjI6YpRI9wbxiJIMWTx+QHB7cX7S+C3lSu/xG+RX9BU6j7TYduGJxK9Aj
uVBM/3JUJQ2r+0cmNPU5IuSpZz8PV4VXkSBZaer3N8nfw9CnOSERqnU/oYttmqN2
luU2rRTduF6A+wZLtQJkulD72YWRZxM+bIJuWPrF2T939FDGzWj8v8pR7xVGDi4Z
6rmKNku+686d6SAGqIsFwD8VPVr6gwafW3dyBLxPErzZsnCehCZC44KU/ycyMVrE
pDAMfeT8v+RjeFtDGC7QcsxLiBmyMx0DtqrC8mWZlaMxH2/nNyFCkMev8y0OSZe2
G3qeS0usIYW4n7qim2tjyo2j9BAX06eG9VJbaKEkF9fUHHwnQkItZf4NQZ94BSc2
DfISsbhu9KEep9Zb8PaSXKR6KRlj7e/BPGAgCkF56xWoCImHcZD28UWptr4Gs4AX
SDArFwP4kn1FwmiArWdalJg+o6xvx693/LaBu795hzXDenlAoH7N6IC6NvKmb6KC
uTVMgfYYhqZdTKwmbTAnefXqpU/FJFO673O62yvC8Nph+JEYZZ7OmD6jUk2O4pop
FjbLS8pwX9K0KmLyvwblpzSYTWV1vGNf58CaAMJdiAcVtoxo5T3Gt3Nd7ACkqoDi
KP3TownPFDjd6bGNCVwc3mbKPn9gNHJ6ot+yKZVd3H6XEN30GlG0wGjU97ZdALec
gp6Zh8Zi8k2FxKLjjzFzhPu1xhGijw+YFnQ/uI47CHkdDGaD+/vP7N6r/jEz3vZ0
QrZwY7/XzWXrO0tntJ6enjMAG5e8xPHcqZ8OgpoYrHjJpCAXqlHpvMdck7T6APxw
L2Mnl+b70/kvFfn6pcI74NygcVaOnxdhHIBv37wjBUvUeLs6aCgfSDijytELCG2f
5CnzF21XF6tyZlGbL5pXO6XQM6ny7Rz5q9AOoRywOJrZYLZECrZvuEQTqcONYiq6
mxc+P5un+53yGup8r+1wl1SSXLX44tAE4rFtY66QcM5csMJkxg69IZdhmpRoLEdn
X+Zql5m7xQfArqHOYwxyxMO7QsRX9g9Fe0xyjnN5pZEPLJMLAcYZckPP+kXpeij+
wQGwITOh8zzodNNgeYmyfz3McHA3YZbXWKIl/UBLEQAUgWwba75qo67yuIaiCSbf
t4EmZBB2lQt9xHAw8hKhTYN8+TRwAnQs/VkhL11HqdzZkwg1cD5l0otAKSpqt+Yk
wjUNAyxmnYwWvtjMYLNcL4211zVi46plRUO/ya374Rz25o2iyWwj8bNkoa0MJxBx
fJCNnw9Z1xQLAxKBvTXExOQiP/K8N9MaszDcH9/zxU+VMTb9sMPHjoBNN4jyTf7v
z8AhA4hR3VwcJnru/SURdmAxR4XG8V6qNqDgFjgpfiwqIgbLy40DIORVUZQK7pXi
tT4RCHiMdvlvrk5NNd+J6zq8j1OAbpdIklMizzYZJ3T8FN61+gh/YhYO5kdEX9yT
GfVfVj8DjVgxRByx02PbI7EFqbqdNKt2IuB9Q/UVf62yykY6nTlfkaG26tbVjvTe
/WtK2aKQtcT4aCRE+u//cHQ+dAVs70A1hObsPcoOp0XrF5o8dMxAoHG0vy9p00pQ
QLXmAla0ZYf8s7N0j0FFomsasHLJlKZambW+KD/coG2RVWtBeYTmQsuIsM7gfKb/
Cu2Pcsykuy7zYrP+fK2uczyzZ6bq6URkPa7hVB1PibetSPVWoOAEWgX2oiAAmbhD
3IMVASjTMe/QIfzP1PelBrUujZkvGO3kk993dpETcxVSiBHVtK3K/c935sYU7AkI
tcl7pDOePkEIDGobuxeaok6KEnlxhSRYBeAJviwOZnF7Gz9+pFA74KEVNfkXoO06
NWCGkdEcUaIgv7UqR6JMIEX861FADAo8NSvm+RsbvV+7Jbhta5YcE6ACrogn7tx+
Gflkj8lPIFSZet86XF5EdTbvenEGr6ZQSO0P1ONagdqQ4x0fAXqypEjgO8pml/n3
Uwuzpl0VrInaxdJiA3IUSPeuSExPPrAm8tum0CvzbPzblf3kJWGfTHz7ZBJHUmAa
3ZP46FAg1vrsKsnv5uQMMf57C6yhtQwY+oUkk6Yk0GUqf2u++9QjC9rgVsMxR2g3
19Jy2U/t8b2lz8JSqi/GaHeGOZboFazNPhJBBABU2zfD3rOaQO5t1aoB2nC35xZ6
SAqLs6+oXwQMyieLEhErq7cDzu7PrAaz/OjwjI3AOYjzTj//rkyPwyYv+QeBnDST
JHz/2bW7dxvU8R3rEM8Jzr+HV29NrlUw5C/VqNkGxxtb4lqH6KOPHm1EYuawNVu7
Yh1xlCIW3XCCYAT5LIDZfwYpn4LKyMIHKNPaOSIRCVBM2wcQeLT6zjl8Kpg6na+W
p9f7zLP2Zs01EQhnNJHEEWPrxm4jpqZhKjWmewCqzJkbLjQPvH5yGxu6goxRJk+G
ajxvt4j1/yF4VE2YJB7vyawuwCQpt+aJ3y1Vx6Q/+eyLvR16/E0hZlXkGNQVYFcT
BkmA3mIMoh68otY4QvZqBw4604EhlkawlxwUDkael3+DFoe2TS24+W/FDLo0Ys6h
6hKvO4Rd7BPCBZTFAvzySl2LzOii3Q0o+wvBbx3B8G04bDFADIqeJrDz0z/JWXo+
0nnV0TJKi7V1z8IvXVSIU9gWUZ0scknF1w1ZJDtKPnvWhstDz9TVt7ISpEwRwGUd
NLuPW786W0zVJ7n2k+vJm6nQkT0uveoyagSapbIcWSVArXKQCf7EZBWqPBcenbeQ
NaMbnQPjodDZ761L3K1TUihxfmdeQm/h2OzjhcM1LKcG96cMBIZu6i2fYUJdZnww
RlIuxlKLZqsG+zHRzoq36q85OSQ4BDHAI1U2y1DqEipk8DqDZPXBlt2DFhtWZfHW
XL1RVky4wEBZvStmL6Ai20vu6AATm2dLiQveesN0qGY6Q6VKBuNqZpW4EBLGB/1y
pnBwepLPXL6bW40pE2H+2M/Zb6gySU+BqTzO/4zxVbRzhh6/dfssuGvipSUHqxvY
yxdA+uuIh5zYkkhOdVkI3msIPDJ7pFbaLlZfeIQGVGVPTBRFEcbLux+QPEkWQz2m
9cHEPqvo9LHjDYyZJ0hm3hsPGm8dbjXrb7k5SX1lrFa1bBUz3XqWZbZCJuEZJO9L
LsCCYduGKZHG9UMowc4MC/36X360Zfh14weDAPfclMDS9zJFT6A5syRYP7Hzscag
G/r1SqkwXycDugwCvi6bPsGfD4HWSgGlKWw5lZzqgEHg56QFFnvJLhWWcsqNCRWy
qkAEGjaiVcFk4MdpZ+xKsXLlx2hBLR3WLMwgBEti7u8+ngM3HrCj/yKxMPa6hBKb
zRzEmJS6c7gaIHQ8GWfsFlvDOwGxdqWdJhuyKAY+7oPUaSiSXBzPw9l0Aq4zEZmT
xNby1tkBNJT0FhfWnU9tjcwpjI/C1Anux6OGqho3inj3i+o0atecKaQYQGgffSOn
OJzJJX/swB7pfpEwtY7AFCyaZO5oD2Zm02HEoO39GghzfYIBMtmqrnuK3hXnvj/v
nE/WSy8td5mM+7mI5Skfh9J82WnJ/6Jgl9AuAG0KO576VPLjH5OMzIIxhE1xbVfc
A2+5BOVZpof60X0zT5cG8/gwfMk3uAZmHLpB8dTlj5EeHFNUr/rwQIHEzlsY4i3g
ppXSTrCg1I3U8QiCk1KSp0NOzMlagYaJZOLTl+9CJvZEQMzOGYK2hbXIHzOUIYOW
P055N92soiF/uAt5FvcrIX7+ln+Mj7qBQuQWl2JAcbdDtNWfSrnrKbZOriJ1dyW5
sKxdom1zfmobV+DYjt27ELcQRjk8PPh4ORjmEP/zsLpb5VplQIJ+9nMvH06oJDEP
gpoia/q+hwW/khNXTB9SbXVvmlUzUBnZ4m355BpE5SIJ9b9LDC+kdmtXmmV+ioB7
gDbwww7OXV6o5/yFx8i6t+HcquFClyadgjnfOW470UcUFG7guaVSRezPjeBg2JLN
ivZ7rIzJ19eLFb6oMZU/zFSHlrgFRFt8dgqM7QUyv6crbxnZXok4fsXqVm1NJd8U
zWSGl86SGNcPP4Jjj5o+gZqjGmci3iSNrEsT3auxzk7wwxnIIhmhtvxAd//So8cB
qOF7ZhmX1ilCdbYqM6ImTW5yXfCexJdLR/7VVxLW3pOCOdCF3abYwD+UM3lelCyf
h8LQF1yb74cBCfpKkzbes4Ywh5iQFEf1n/Sf3s3e8tV7efozMQxw8mXxVAGB6UkE
ZyfSNRYUIreFFf9Jl0357zhPqQPKR+8WhUEFDRIbS45NMW/mzXps++HndJHRprBw
oKlwdxpTQdLngzHFELS4CA5xOyc82nxyI9T4Tk5AcEkKTiIyc/r3N8N6CiTB4r3W
V2L7S7ldg/mXWwRMIce3jsOKnuz5LC1c/5cx/T0DC5gfGDZDy7WUz4tSazXZ8GaN
c2EeUDjZWzo5cwahV2O2F751Gnf5uLtDDHPBP20pls6/5qeVgdjgg6wW5g3iqfOe
wQbjq3mT2fr6Lp3asvqHDvhnM5gWfC131n8wm6N474UqmK1s0T3CpHNaeltDWU0u
ORnAqdbUtU2rStbgbNnQW3c1iSMreSoHyzUjbs7PoDsKfEe/9WkML7lpTE7FhrNB
aUMDCgXTEqs5cimR95+7Jq/rV0n4hhEV+qFDhVdZDi4VN9Es5DydjwiPOKmESWuf
TshquqEuL/xcN0MIPH1qN2bAksd22PeU46jkT16Imp43IU6OyVrEY6YyAsLIWCnv
jEPcbuY9eAYUHY1q9EnIhknLpD4DOpFf35BEUnYWnjL8tga0MIdGwAUhWKJvD0mW
6IoNn1r9qeIAvTRarre6GGBUsjWkmoE1Xwf4iATLXkjOjyNL1/cQwx0Zasw8HkRS
F7CSX5eTRZewoZ5gLG5bMMxl7FZVi54u9TL4HQjg6divAJ6ADGBL5j7VhjSP3ho2
o5/WrQ+50qmFI4jhcciDve/+hVZafRkEVhTQhNQ5DYnFri6BlfFdo+Ed2FkvpBrt
0Na0+DvsA7d5pfvXlNjP1jiTPtkTcpY48ITHOydgbPF+3JPtVGDXHgolFcw9+3Kx
Z23bT7+EVPBqEkR2c+C4r3yPgPWNzN+B/OzvQQyfLN0f37Yl2j39cGWTKaTwkZU+
XUVp+BVJccQ2bodGMDmRbNEhovNNZ62w6kCdix2pp8jr5MJw9warOZdvR5YC93k2
uMbQPh4doBtZjPya/GaPsiTZL6afcGOediSN+OCvruSSGOB/0fCAwP3nmt35mO9O
w5RbX7gAnSH+4XCcbJsPZXsWjYZyWTawiQ0uYiQ3YvFQDpUAJ40qVyQhnX1frpMV
x3uF00b2Sr5c8R/Cn8CNAee9AdSmYvcykzF5G4arOugov6VPOIyztDCtz6qTl0FB
ej4Ngpfyj9NLkAlZMqJYFBaYIBNzQ7nGBmm7aNLjcUEliCcYJtbW7E6Sqjhfn2PE
5r8e75OJbDFE+ZP1/h76HuXTlxtsc+5h7R/QeXew3aXEw+2o9ojJSRqkYuxxvdwU
WCtSkQ6L3rve8YJx9ypblOcF3G6NuqH16cDHy+rKWFpU/QxyhQkfWaWKwyI3Qtah
PgsZSEjup8oDRapovufTfhAVa/f0LrKYB19hZaTUVMY2bMIKdoHnU2D1eesozTtr
HdDjHEnw604vK5yE4EZJqBamNWmdogNMZeGIuQsFh7usTXOCRq8Go9fSlvW81yu0
Q75pSI6frY/8Ial92Luq+2+2pe7SkXtZnF0+Cgni5LeSv2MzTh5Ov8oLTwHdC0r/
V04EoVAE++CXQCmoXM/T2BXwq0rI5MjMx8OOAIB/d2JY/iOjY/6zMEMfeHRzQ1Vf
kZt7HvdE5C3EqbDJgO/XmIQ1qNAByVVGbaSnVmZnEWItFRG5ORFoYqn1h6/VpMVB
xNHmO9bMeTukmpFNmhdow/rqgYybIJatOCwx5E+nSQUFbNnxTzs5D1hjMyN5zb9u
gbSMSzpyuka0m29auJYmmMv734t+ty5vK2BYlkDGmtW+y/d7KFMsJTyHJyHqIYjM
dBQ2UHnyfHpjqlwIxY5CL02EuBVw9TWieOxpMF4fgQTlsYVf0Za/FvfPyr5SPRPN
CbQBBBjT83eQu/6wY+v7WBmpc+VUt0iUUC6ZVov1YMrc+fZD60Qf2/qi47NL2GgY
zrdbzPkPBY+lrOLMuTa8a40Xd8coCEtOngPZZHD8uSmRDS2bBb2LH16ACjXqXMvi
7MJZD3vFYa2PVwYC9hdF9QyRdsaMtMXxSkpn74Ot/chiizL6sMUTnJiXG3++0LAE
px0PScjtLUjG32eSFWXA8hqiLWNxxrWJ0U7PUEM9sUmKwNSpLvRq5rAofsQmLGr1
HFXT/sZXQg6VE+XWtt0v9Hbv/XTcsDqN+Qe/nzCxuPLOKimOhi8FKcX0VmK7RNMo
vili30ZMpaN88WMoT0EFZ1tNhRhuujN6FHFj1GczqviovL3heL8A53SR2+8G6bYl
kUFKjkbih6WXWTT46A3SVXqDCF5nNLP3lASTPHyBPXCGVXmgGetmAQF3KJfj/UG/
isxWF0F17j4fp8X2KxkszGooFUKQMwiztBDjzVMaaTqFuBc9CAca455zXlOlZ1Yo
vlSFlKkR/vXUVhPYJKTbIqBd++h+ZqHQ83VOgDoZ0tXuIweOwnEWUACOy6BY4lzV
c8kro6reFDYSc5eL8pWV9DmOuQHdzPTdAn7du9NIXH8PbbUHy+ZJD6S4HWfq1ocf
ABW621HLY5lijkbVGpU3U7gbvCNW1Fz9hLRY+bV23AsXEwzNWroOBDukpzAMXxmT
voasooiTtAo8Y+Ya0yj3w/s+gtArAc2n5fAnbHKu38fHF0sbjBCsV1eG26vH1cCC
X//KqxtMEAwV429Y/XDSQxNncFAY6izi39nBvVN0LfbCY+JceG0HI+MQcY4d/lO/
crsXztRxXmrFlUYwCdMBOFhKEpil0AZKzrx2xkDlUsW6TrJQftNms3T3Pg41bKct
1mwEnmp3WdtJqXK2jUJiyaak1CABpwGcOO9rGwHNYLLtRjiToO25L7yYazbiKmRn
ZYzQ4hoomUJzdWOf6Si53khUIxEqb53ne3jGHPSJ9ylIZNAHY9S0cilW8/skK/CM
6W9u8OggEXHFfwSyKBB0M4+kfsXuB7bbslVr6qaMSNdpFAEMQfmSnJj8BKm2YKGz
KvyEJ8Cb8QZnJpwxlyh4jgAN5JdbYlv5yqorieefcHV0XBl/Fv9kaM6WQZ6TCwPU
U2kcgdwhtmm0gU0d/WHPhCAjqTLeQAA0UPDM3D4IZrZOmA2JF9NDY55HsES01DQ3
/UgVdRAZTN8L7T3a9Fra3LaBwZFMKpmAb1ka/En9wwSwFMXumw6EiJTfLJbeED4/
+LMzhdSUIvVc0W7RArVVhUzenBuf8p7/MC0AIQGmEpaUvhEa9ELXJFgpGonWtbeV
+t+pnGQkDLUG/+Bx8YOYcSLW4CE2MLFFDqj9sSMQrvDxM7AQoR/lDCWA2f8Lss5T
D1ezll/qIKaz8gWwFgHwh8NM/zVRqwIwI9+elydBHQzRQbAMjxnNwERXk22hggtx
Q2tHWI+Gmc7VRHdbUdwPuNO6GnMtKG1C4BYoZsIio/3ejQSNGzXuz0lw/grlhZwL
irjbtSb5NnzO4WQXy2pdr9TQxYbC/q0Bpv6NRHBMJxykzX/K32YHtFWp6aY6gBIP
PJwxc4SnAEQujZD4YCaZ6TEgxVrNiB4t+Krer5LlS9utGORoBQq3OZtCsK0h8960
WdEriIALOCpWghzbNvXtPz3LMlGa+/A19jjJhbDJCWAnLeU9EqHbZvyEmk3nersG
lp2jHluOgWnDehnQNuijlzltjgwJv7ErsJoST9tvYTeMpcxgsz0I8/JEiqHnH95s
9TYnR+VQ7nKhs4F371Y56tKoQleYjN7gU1KKhwcw43cKPVaSOgmr9oMRfEmPOZB6
uNBvr34wdqOeEubuDPqeelrCf0/lCkfy6siuldH7vDT3LDS2Lu9q+IlEU2wNSe1+
QzihfCxhLQWcPLVJ894vo72h3L7HP9lvXNgkOlw+sxzvegXmu5eV/FAjMqDavEcp
5R5UlERBwRwWro4fGQYYaHO2+6HKYqZcKlfgV6O2kxkDZ1J0RvxUKVpXVb32/bWe
Vle91V7VRgGzLoh/s0KTpKOSAIkOGmJd2J6FcoXpTAay9zm5YG8fOy5TUeiMQB4E
d9nn2/eG2B9sLQmvHtyolUBNg423wvJr/OtopUiE3hoV4k0chmYydv45rIWBgcn8
cQpfe2tHL2VYpN6INLa5WO725mCFtls5mQK0h8e0+4PwMgm4E6VGU9JMsCQCumOG
DWPbjjnCSj9ezfQ2MEUf0sWDcmEm1OqIb11x0dBr6+xh7f/anqptWOcwfxVWvmd+
Poa5GEC/yyJExjCa8tlc0q7AqVtnQ8VKDRUkp1iTc0m3sEWgRmwbRSMJHFoemlws
qQKONwwCU6TtZWkTRYIOxPsoGGlv8LahvUJM4uRYrvXZmbbDS5AHxUiaRUxwSGMa
FFzV+/qPJpJ3PfiWiU5fNJk5bAdAOgqqKFDX1ixjXo1fyCianYxNr8RqJ/BNEU6W
i2hU/eQTTTQjpkYC90X+xkZCypsv+NTCLczmdv2WPf+aGaPNCfHr8z8RIxsNrZpq
+i4YcHbaOiFVf5Ol65Uaq3dQUPuSDTEDPT9kfxgMhm0LAR8kh8Qc8kZgaw6kvu9U
VzRy+uyc8tgjYYxix9YiRJ6lUGwwZp/fhqJP0xglpDpA5xpd5nHvOP6t+9NXvPk5
SL8LZz0bnvmZQr7W9uJ6YA/e0HrsJyD1dxW2RS6hgLTcDXZxtaftBOVnKPEsvLeH
JXINaO4GMcK3atJhfKnyEiVvIBYEPRcCYqFZogZ4O/hNFKb1vnukApUWRniJszhC
OFHlAUq5V7SDER5MaBO+QgEpGVFdtuvw1DgrYHouu/kOjOXv2k2l91GjqQY8Or3W
U1f6nEwtPD1h6BJgVwdOkwOevi4SWucvwe6nztdnIgDBuBhVElsdlgznkqoRMKQl
x3WERRCxw/Frmr/pU+MNqMnnYCVlc0eFtQaIeafclNvruDakMvfFJEoWKqIoWL76
7EfyIfD7kGilvxYEIA+5Xf7K7eNq6erYEYyECHk2Pqqz5GIX0RYyh+sy0aT4OYMj
ThakfhGDfDpwUDJJRxtwDOgUGI00MwgQwsmqixxgqlDXm2ifDYQquQ1sSHQQnauQ
pxSKUUkaWGvB9uHI40cgu3B8kHnGLn2X3Q/TBRJ+ikLMrq8H+hlzv8aO++2UJxKQ
9yNTSZ9GIs72Bz//odeOEUHSk4W1NY8KCE8aw2YNhKbsedZ3UbtDRJvnEX2aJcON
a4u+3KGT4+4dOPdJ5lP/iPK2hJdSlH/sE36+ecWmnaghQ72Mf5JtdtBpaZCBQEwu
CSwtAvSJ47DzGlEAw4xRd1102pWmWXyd/erJrwpuOLtA9kH8tnfJ1qL1QHFsZ+eT
kp7/cjKTonfeINOrkyElDUwIaEEZxLJ9RDZXFitgeJ7+d+uCMtkezkJMeZ1+LQbI
LDKUI274vL4K/ao0a+eOq2zGzwfr4CGZH0798oDspiD0S9I2GI73bdSMOCBhJ4cI
MlCp5o1scHhtZfLDry4/G3XSf+2SNIj7ih1NV0Ju7+KVKuYoZRMWPzKj6lG7E/Ma
W43FrfU5WD0+m7Wqt6rfACzdyaBOXqgHptBLVaRRDxb6Oe5M1WHBukCP03ksumjC
c4rHdP1jhPFJFiY36tLSosKfhJ0gOypu2NWrklesEE+vy/jqIEyGsFB5NBq1oBbc
iNsMGHwlVzb8nk3dyi/RzMkHTpO9UZB/wMrEtjOaVpgK/e+8BTIBoRcYuUtjsh7y
JvbfEbjKdhPk5jeCn7yXFd6ylstEYUT2xnStMJDvWT3/5gUdEoizlKebpkNnw5it
zLnYl2I3jRCVrH6N4i8pjW+o2A9xSOm4lvPJzum4K8dYhocQLbmQXNzcSKDrkB2F
dE753O1eK3zUqQMIgu70PahatvcTAlI8iqtLUnq2s8u2HL2291ak6BPOJUlzx+mm
/8DEGUumVGlO2CVao0t8dP8zfDRRaP6xlIfddeKaXMXhHcfp9FZv776VAbl/FRqK
oNok1y9AVRA7VRZc74PAKqjJoXAEVSUtBZLAPQhPjK8gXD9m60cSVkh1aDGtw2pw
uia8ZOeq55iOyPXA6flAP/ZsQQN9HpWTYjyKNP6wSXkIcQ59inbuEgxICA8H/+KF
uglCCWm6BVKgwEayLcxJw86MoGAX58FmcT0/DmVfpdjRyC+MPhQIH70RPt8dtC+f
3mn0OTW6wUf99/F1OXQ4vU+QN/MllqIYHVx7NK6cHfbNH65eb4BV0jXKcalkLM7u
iVZjU4y5AMfSM8WS9OpLZIFtJ/yReXbhKQq6OXf8iQ4gsVgpZ/zxzdaBmk34JMyU
B3gvkKAbnzidZEaa+rPA/kIJP82cnncCyhrj7ZsDhvDv9HjwwGBwKXvTPd8KEstw
G7WIN87ecdJ269C0CGjDXhy/SCYpyl2E7+ows5scR50PvxpoB2MdqxE/1oo8Yf1I
C9DbfBjGbTr8uIWGWpRMzXvbeRzyTmOQ9yK+EJeY9buPsYho6gOImJYkejMa4iIi
Rzwyo+cRqoS9EdGksMLNt8laUS51BfJbB+ru57w9LcFNJYNpxrgOW/H4+EownKx4
yWa4xXtiHqZTdlQPPvBY4Gle3YzcGGNngDVaCf7grYbxIZk463qBzIVkoWb2ujcy
gwqzixeM7fFnep+8n2xi+ONDotdbhLnqLreSVCIcfxCrJ5AqWjdF7gMIjGeajC67
jy7747Azzshp3WlexPgwTp/MODGxIHmogTac3eQ2PQlmns8KHnEbPN0GYuTepmnD
DGeTTYAmERiV09KrpuD8cC7PZqc5tjZVLOw1hVkjX06c3RK0cG1Q8ZizN2CLthrd
o6gx475ue8tvZ+WMYQt/QmwAN0u+aujE+nN6IRHWSvRs5R6MImTtubOXcwHlbeY/
XkeSHn97ipblMonyfETR5b8qgWlxaDkrWOCqfSMcis2HJT5DMUgBPbJgE7nLrN8/
FNR+i+NsjNZdT88SdPckCVY/aOMsLD3lv7f5Czb8fAX9I9I2z6hZPQ5VRestYLV0
DWkX8LznGaycqIH2i2UGHQ+g9kwgkyTNpjcMmb0Y69iVj9Qw1kbEWrRKHxcEnjxg
LU8IViS4k1Jmw+CbjFrZtXjF+GtaOGgsj0CUqsjSgeumlKhTonaploTk0qTmVY2W
aD7igSTFLJN3q3PtzMke/JU6am8ScePD0JVq9QvD3tOySNRiKpP7AYoOVsn21Mg4
6s+iVB66vBL36i6dXWynLNIi+C+dvtffEyCLtgWmMNIsD3vdDX52JtKk6e2UN3Ze
e898LUwoOMChVAsHvpI/drUnS/Rl7V2jfnEkXSqkJX3RFONgQrbg3CyNvT9LqMRp
R5WRCO96brrgqHGiPctJbpTdHprzHOFhu/M3g8vYOzl4i9d/Cf6k6fejXysDAEPf
V6nJ35e3NxnKA3WrnHoKg5FD5oomdDx270W64GFYRsyC3kOGjRAmpwRssXFKvlwl
/8hrNFim5d/mRKpw6+6suLDsQnu3TljNRISwqx3F9hxOvKywK+zJrtu6TYTaeyZP
pUByUWj3EAVQPdHrlFhCxpE04sQ2Qo83RfhM7csvhO3MqP4WhT09S5Qi+j9RD+65
6JYgttITJpvLBC+5DJlO7RzgSNbsXuDXCJ7EqSXVy6VmRSqmVE4GAwjamHbgz3uk
vS4Z28ustHiUnb6cWbLxhbSVU4kmDGJj1t8hBY9YL20WwpOSM6cSCcS5WeJ8nQZm
dCeovQZOTmycKkyx7omfazKzGO4eHVNmfh7t6NQbJCR4qUeAAsNDeJ1+hKVSJbPP
0Z+PVnc954Lh2BmiX49R+LBEwba5Nl3Rg2CyWG2Z0aOY6YfI1lTNc7zB35qLLTTM
6pANLrk87feNm3OxelcF2FYWi6b31lVmAFgrvLeQEwijDNXzWwSbLHLbBQdLeNnW
/F2XrmgBKlYFY50s+Ru/LyzQZ8E69R3M+x2IVfxNG0vXmqsUuaaSlbnjYY77FG/Y
L+gy9V5gQtPabUhE+vzVdxNMX9sWAqvNd0QN3sKoHVJ+DlcdRFzFeRs+5GXmtlJa
PVetOejkEteB3A+ut8u3NZLXcmw4WAHwd2odMSRcQ9kr+E/W4cGmuUpK+yjwLx6J
szVYvnf5dVfrBtEl6k16adlMxbvVLKFUX/xRLVtCtv11ko6bye4Hbtec7B4lPR2l
FGlFeNI0vRhEBU0E74637Jr6gL0UVZbevvP8xTx4pxGqfsGEbJ9cPFLpwOTv1Ww1
wm52dQ1FVh1oNP2xvjqIPUOVeSbFqwhAC9/1dTonyqgzJ5LC5KTzB/NgDs7D0qe8
s5LMBnj2PQB35DwAlzn/kquSTFDjQfg73bSSyXGJLSBK1k2ekiIdQg4jdR4JszSO
A9WCpUsPDpIUx23/D0pZUTKlVwrKQPjq5h2swhsuBOv3ymjkqF3elRMsOb9O8kCS
xHkyimSYw4vCtZ/Uy16n17CqtTsRglQ9FARHc29T4yn9ejFkJdP9VgM6GfTx7LQk
3zxEDCTisqFOVEnO/Tjci2ApIslbTG+DfveMp2hevXDtRr1FQREh8TsCLfLwGQTt
hlrrw4Pc9UPHpYl33tiKa2fI4E9oLyrg5xvzXYdtHUWlTjLmcwXd+nh79/PLtBSq
f3jJKVqWRy4g0+DS7PnYRUtLOfn5LwNfLR8qCVqY5605mYSIjuh2v4mQCUaMi0pv
zmrvY2uja03w9bJIt3FBOllltKfh0I3+pjXyFf/VX1NyUfbOfAwmHEsUsbO+bR4d
xooV3vahVe1dp58CXjjS7QWQ844yYsYIVT4Crq92FJZd+G2FwuJyYq/JkEsH6kCw
oIPZAy0o4TIZyDp2G+5gBqEVF0j9GX/U3wN1NfW+UyQZJgm4DIQL2x8ay8bbtRlU
gEmGzMaY6D8UwQJ3hrCTqaWKFro2z96sUG9drHi3mL51cMKzm3Q45SpTteMLM3To
KOatFl+nBFyJjlKV6f92iJwfv8KoZDiFP5i9mSw0qD78wo1QiVbPL2LK2WFdG5o9
OVPHJnp7swd5VeWFICN85SMaEqOuqO3gUPRRH+vn2kEbZ3nN1qr7PmMB8UJK2Ch/
dGqYs++BmzTOlBuyyczuENXhZTJN3R29/dCQOnzc/JZ8Ml8Ov8WvOMy6wWgB6udt
MnccKoCqEDRzP56k+mkAF1Gogl8DjV+XNhmqi1ajVt7v9IfTdmBc6yYkd02WAUAi
uTHQm24GKpMTZptpGPs+5ON3Ma/9nq8hPOp/Tr+ivY1LB5FWYa5IQR84OlON04eT
g0x5wq73ehUpaTERGn119KBjQ7zGcfivJpszEkdYsmp5k9y2GopWZddNtjQ8/1Nk
ZV9VULrCBRzLeZIp5QuHqnO0tMX/I7MyjJkVwsiS9iHtiTl7ugAXBvpXoSp+FExF
64EQYauMBGYcyScZr2nYMTXsypsH7pbiegpTiGj/YHK9GfdPKiIvqo7u88y3qLq/
MjGphCiK8y+XE3P4Ws/LK3Fep6S/rI/5vACVoqHHcybIsgSzmCOUAKqoN6/ng4uD
dZKc4hE4NZOyZRxM47AFhCiLQCoNXpmDHoVRSNAgm9SXNnrF5iBmXelYvbuvun7I
5AJ7UkXZIfc0UDTeFeDeSaxzKuNhGxcrwwyEyke1fmmE70M+aR1AeX15+BMiIPEA
y4geeFpaYD6f5jFscn3ePFSjPoYcwmYffewtSY7wUEjv9Y0mPH7PjBk20m3930ds
6aUJLO95KcKsl/yxteygeuc2IBdvIgXD2wnT/CeW3hEMeC6ddTLoYVdrFE8FhxgG
MVFK0BQ7hDvkRmwIoFY5c1Y0SHNPUa5NLcnrrIDHdsyeA3pehwVoVrJVO5ZkJbsW
lam1SHjNW4+MSQC8b62MyZIcbQMybtYQNbxtVxJ/Ifw3vp/MAfADhtcWDIsVSb6c
90+oRq91+a1zyv07ooy9YZKbWYsaq6QIC1mEwT0wTTBfy/2nVzjD3nqHnCqM1s9y
aygz5Q/N5fZBzaOjjUxrVYBEWtEb7SCuBqRiY91/KkLhasmjlZ3D0Fvcv/s74xhR
0QNn1cgh1Gu11eWlKKkIdwB52020ZViymsL005wbF2VOXpDykyfc+nc73ZV2HT+Q
5z436Pp+gySDCugGz3cYf+4QSIKo9CP/QI7HCaT24Xnuu56PtJ4P01Pcf5xw12MI
CKcjEDmeSp492NdlF27SXYpUThXFDQSgzk8nZAyZV1FuyF6R4A4Nx27VL2rNXNkc
12rWsrtvfUZN97/lFiCrUMPbAbc+Ppn1gs4MW1AL6CXDituygdkQqXs+1yDIRrQ9
piVZtPU0ML1JYR6OwNlqmrhtYop843UYlsbkI766Wm4ZgBrViD0TAhbF/BJEjl/d
6yKBZrDczLh2oUMTc1c255wfq1AD8gIqSTHGCul1ExLbOJDXLFKmn7kXE2PpmnfN
eKwKKcvTIwXY97EImucGWC14pfZJEZZjWY6d9mmnZVBkSPyZS6VudtuwN54qh4qh
aSm79Cl3EN1ClDb7yEO2umqKsys6ENjP1V//xUC6CLX2EBQhfE+wCQD+IgGj+wh6
prUbDDU6CPz0xw/Wh4AQHnRq8qStQ2H1SXCZW26X1lk3VTVioF8R784HMBB9dOY2
Y7MRvEmEwKb0Eh5ngxecyeIw5t5EPB7OkF2cQjxX7eEfdi2/AuuyQmzhmy0Xsb3N
nCWdVzPftQPCfs9B2CYvaSgWE0HGTIOEhqBQw7B7IRsbqTWA7kTHxskiydKLZD6K
uyuIcE9N1uwA4PzRuFwA/R9f+hWglsk2knUn6fgQbRRlAOibIIHLJXsnDNGt5bjH
h8OTgyiR/M7eixJ4lfdaMqstpecPS9vR8MTo0tLJ9IHP1I0hTGqAI1bpLjHX2klV
q9tO5YtyQlZQeEbhueG5crLGw0Z5xAPDJsjeHc3Lum2iqWoJMSTPtD1W5kEK1egf
uQ96X+CPNT2H1/XPycgMBwWSiRHSee+1vW/8FkT8DtnwMzE2jqroz1W4jgQ0f0dp
geGvwT00lXSVjxe6k6A2j9fE7Z1OltpDaFZ0CtWKlJebXAIBlG4wl8su8/ZzbNdK
GK1qezuDT5HQZfNRuNlLpAH3P1XPt/QLjMRu8MqmFVaZbIrUq/p4Jpa+zaTcY9Ej
FF4JFrRkutmH029zgfHhivajsOnzacdE0NwNaoAC3q/V+UTvqs+HWxmHSgS+1KMi
xNGcOmMs1TMP4IaGoUWGJNXn+KAVXGwStF/47XCD0NUdArFMUesxft51gZ2p5jgg
TEM+uq6UuBZ33VHapMvx5xV8AffRz3oTKTn4442yaCftxBbvLkP+nvLQyEvLbbOL
nSu/nBkYhIHM7PUsUWfMuzno109ulnPMTT7X7fOhrwWknF5uO1sAO6e+FcZ0/NHk
y7t+R0AgBkk1JxK0KUAHe3JKKurBqAJ7KdruXxBGngfPcFDpKhkr7E2fmnGodkzq
C27dopngmbGs4L1M4lXaRvjBClsai++xgZwUtJaKTNPmXnAo8rSmk01dvDWpBN7j
2r35bM/cok2BhRH9B50bnx0v+XP2TZ1LMOTwzVInp4TCH7PtYrLKFFFv4UtapGin
9FVWTVq3+5wQ+sJtD0prZ9nASfS1PvDzTBFWxDediLlyh25vYNTyISowUce87JYW
JGXDeCCsiqAuUwPaNXTTr4MMHxSciXTpkfi6HWUBdSHOp8qFiJo2tSv/Unaus12c
kDR4x4lFU1/jry/BWKZCGR2dZJ+nJ4WASXwog48bObnKhjc8DkqEoKpk8/wYlGX9
+aPcwcnAGIpx4H2mNX4X6ua/ReLEW34ULa32u7OZxe+Lp+TwC3C09TNy5UxkxCoy
wAnYwa0Tfposa//95eOZWNaB3oZMNE3K0yN+ZsGPIWXRUzIpN67qU5NGaBNBxUCR
nknCjVFWZqixS4yimeXsQwXxOo9dcxOF1CeaNOPmCJyPGoXAsMYXQiEzTVEdVAx8
DqVDVjbDfY5yBCBn6X2oQj74opop9lcYPWZJhfpq/Cj4A2LePmVuN9BTX6Sxt16S
cD2vx8LdB2Mq2UKGulYQP2AGJ9Xbrdpy+XqXcZpE04Cn2Y2uo8tlP0xorlTWbjXU
Y5lYJ2fC+5BSogUfDh8nlF/3sXvanv9uQUiN8iiLZewVRQEU8SmxQGgsdyWM9//D
mcUQsAXCxmA26AgjcK/bng8VJPTMFomXU0AbyirFeD8mEGiPmM5/yLRIeRAQgvnh
6hzGOzcTDLvd6nNdQmHke8Eu1gmNHIEx61NEAr3cmgzCXquNzfsp55rKr1j9rOON
5LTyUlK8IvKXOUnJUrqc2W7LLSQnhs0D6ygmX8T05ze3WT6RchPL7oDSff2r1F72
j/sEL+NtWgNxrVSfhUcZMj7FDpucRlk8NPNDmxPeeW5ezxHhskSP8IxfcxgCYiOs
dFGNdqMjk0Ma2Vx4QvxQywNI9a6K2LGjdLVWsajAi/GYRQu0UiavavkV0yInb4hT
VQsmNKHIlL5Ca7fgYA2eJqBZTUXr5bQY1rbHDlZPZUruEFL7CpNfOIfGxie9uCsx
nYfYbcXLoO3JFZV1/7Qc5ueWM4dbLjdywYd3gw3BGhtNzkIjXMiM82YKdyEiiqky
UYfaYqNO+U1sjFmuewx95DhhqmLDIG/KpltfaMD14KbbYnd45k+l4v5FbZ2/7i6k
Oem4tWabRltvNTNnuAPCOaDuO+zlncsJpZPEgVs4V2UjC/8ZPnhRUVGvIRX/osG7
f1T5QYPFm0t73KvRVXXZc82Vna96GL9FJsLX4WxOlffnvhVIFh2v57D7rxC4UfQq
fs7WpdXSP6egsAvDx2jGSotqsnVE3Ybr9D5fxYmj9t7/WM/I2YcjQCvnDyYeNte0
mbALMf3MWSCQqERxp7tg57Za4feO982OWXX9mOCWNb0AKMtWtp8ztOKJp1rGF9GO
zumYkPL+45glqIRakabYie3/YWf1HkQFKKvM+cSoK+ydxwlzGYO46ZynJg7GhO2t
NFODC+y+xJmwVYGR2v4FRSi+RdDMbsc9ZG6uloCrs57LOcr+kzB9xu9oVuiI4fAt
h6T2z6n4l4V+3N1xpME8PO5kgYzAtpsHtzlTp2mC7oNPv+r9IGgoBy9gaYW5gxUc
ToIOf+kWp26UuMjaB/09ESisAJOEzFY8eL93sAFHLl5ueCSSdbVMFkjIo//RL55W
DGS4TvgylKEoGBjGMHPoeJ0lWi3MAeN30ekt+/s449NEFPrI9RG2mMn20aEm2t66
OLilYvAWkQiSHFGitBQ0NPpIQ3FABaWgKdvW2tP6tXm8tsr+R2NNwTUB+HgOicNd
npNuJk2XgMis/zsJJtPSVODgLOK9uHYjYPoOlkR0qG0n3+eNhwhdZkbSNs+FJvQr
+2dPC9vpNL3hK0+SaJlZumIClI07hpSNUaFMyDs6i3mS2BA5Mt1Ngr6iON2ZIPlS
ouExsoMoqQQ6uZwZjHNFA7Zjn6G9SJNiQ5nWMs+jyKqQ7zylX0D3ebfgJLzdsRPw
Gefehx1bfMmQw70SMKToJ3iGlxioL9R/Wdgtlsk8JXoN8aKyJjwdhUfWhiL6DtkG
jrMGr6K0zQnZRQABDDf0xEEDgJSoycTJ47xmu34nGXtnPM8RMZC33+H//SJ4yZnh
HZ9iTk3XsMCYTcLCcTojLCA2P5ZK5VGEqQ47gBnSFRuwK5GsI8OocW0svn1FyK+H
YLvQeFnok4G+G6bkDiF3XhACS0Dc3EMpR1AHrLB/44pXexkhSygQCq25wF2cyCU/
nMSAS6AYf58FUFPWgoeOIVCeXMq3LjrVd0rvPaqGJv4cQC9x9e3H9agZfh0eIG2G
+m3e+0S6BUgTgOVXVc99CCQXbonSXMTUVnv0OYrv9pXySPyF43DwjU89RvYw2tjZ
3zK3CCxbrUIxEAmNKEk4/sL2aP0bki0SilHA+JOOox+q29BY4oHFmEqQi6UHkmHV
QQqY/4hhzrrkwHweQA/PYZc2CPkzsCcH817w9r6Y74cEqb9+6xRgLRKw5fipfXAP
P076p+1Num7/cqTJfSHy/uHgTnPLh6tsUCUMDEk/rXeKF/36JfsJqaaLp8whgq13
Mdpce5/uiYsG5Wl8AvNaJ0rMzP8UYx4M8Lm88Uo3SJdbBW5iM8Zw/+g0WJ6CALRH
WsEHJUFOZVVBKmR/tXnf+IkFD5RsPr7ITEiN7/96b8vw7rCTEcNIa3kFqV6ZDNQT
X4ggmWgc27o6Dk+ZKnumA3fl3YxEhCmbHJqtjeS52cB54g4Zwn76NPbBj7bUdiFy
37/49QfBgqr6emqlzy7WCMMKObqXbBoLyM0ax3PqL5U8ekSJ1/D/U0poaMWBNm4i
qOr5GyFBos0ze0nqXIviO3dvoZN4Zb/O2h51t7ibL0G/9rj1ZR1lFC0ecqnNJ/KY
WD0kgs8rVZzltIDaRlCVD768eNafTQRLyrAcAEB4OlbrThtVXV6+CZifb01CizNr
1lghjXSr97illyj/9xxUTK/Q2oi+FQndWg4AyA0fMihuY44Mw3WgS628HWLyLS/O
63HMcdtzQvrfyoJXtHI96a7lW+9dQ9q0El1sd/BbCJjJHNQuIfLRFA+4pzf/4ztD
Wz1R95BhQfcANUFvzk/AdAwWC0kk/qwfXKyms8afE58BOjnJ2ZPorkOus3mDGIyc
zPdCyo4kGUEHrE3FuqWWDo/M+myWMuhoIZk2AGHaG6qidiG6WKnHXttPqVgAuQt+
lNQJLcc2RZpUC9mqiux+rdaRJ3hP0+UhaRWyD6LWmoPb6QyDpxrsaANYNJZ1sgjt
p0TbzjE5Vzfi1XIzvpymSag63+ab6DyYuksCs5mHgkK2D92Zmnw7A5Q6LKnSL/hN
gdCYqwVnn3ZCEGqG5U4ryUTGJmrvw507k2s++QBJ0TBei7P+ULy/b/DxgafkDt1Q
kwZRGfDBJhuCTVrhuKKsT/ry2AIAU/l3kvVGPWrRufcI1NorfF5gc5oLHa3Pu8BS
8mO74X2kLZh3amrygSyVk/LUtWnmLhwFI8Uo5lTZ9OHuAYRAwG2Hlbub4FQXu+XQ
/B9HwHng+zq+cEAWmsUi2/IGd2aDM3gt/kK9YpQAQWc7Ji7iPbh5N8glGFoSotD7
xUJn6xyrs/vqc2nP0K5qJUzDzJ2CRB4rTfAF7/AE2pNgxBZk/C24kGTDlLJr/7MO
yIXggnBsPMYYvu83bi8b5DsidYD2BbMip/eDjv1EMKUMQKRhpOACTl7VbNVidAlW
mCIlwHEFgYdEE5gqdZI+6N6zexDyessdRNrnwUKBVsnv87030b9Vd9ZA49ssbFIP
k/b2FbdkB+yM1EC1nU21J69n+ClVmiP/Z/bNktFdNM4udBVKBOLvBnMvHrRwssaG
2l+7uSWs1NYFrVe+tUBZ/ZUNrCxFfFV0zugXmekPLIro+wzaxIZVn2lEGXGvDOF1
tg1ZHLnbS+I97xXk7TZ1YWFowECbmXsWCkkfe3p7o69gF4EMThGLqF+YlObIFVG0
ujnjZaR67I9Q208hZKvGgZyLJJpEEIl30VZVt3jfOuDOVxQzbxPoJPZAQWvXwZHN
iPVCz7jWavp9Z9efBVHcuPNBqKl8pfor7TOsXDUFMkUeHTzJnXYT/6z3vZ20C/0E
0UCK5CF4alyw3B9gIp6xH2R6cKhAcozvI+9/vGybaIOKnMaTI2wfW176yFeV+SVH
/b/WdohNpn961+aJP5SjN1IeTj0nnRBONJC2BfZDcD67tYZr+WANLQOQNuUGeYdc
XPTXlo78/rBQqGOKeG2GV74DRAYRts2kIK186PU82jfuYldZPiejga061ZnSNGNq
vgt20QR58fB8MbXgelivWXb/0likj9tLXI4gKQXaVj6EF/nnTfstHa0bq1hiB/fH
jdeMCYQ/gAlSuwjW+h5ZjdOOLE8RiYX4fvOiebovgX2QXM8bkXrDUlopuT0rPU3x
/2WgWix5AIxcbsQ/0fArF0279muyLlP1giSkwU54IXnlvG21xVT/VVXs54pNXrYs
sp5J9WmciPCYTTlBnORjBhYVfYmq4trozecgipyH+rp4r5mAr8ZY3WdEKAlg0b/3
j0SeMWustQCXZhFlwm5L52UgLJtgkVnba0UOSCF3Au5XCzrt4S/a0jYfc8qWSqef
ukjJejrVGFoiF9hK5P/l3J70OsDd5j3RaNwTWPig9gyG2UgYX1hDBVkvucMKxqkt
JAlhCi8ssHMRhtJBoAs0m+wMvWLEsVeXKrxF/grSZ9m9nD0UPQRKGOOip1PheEJR
xMDhsf6/MjVIFceF47UmT3trJyr4q2QSJPu2GDV5v79h9ADjNMCu6M/vdTztvBce
VRSReaacnDYa1BGjEJE+kHXvAKpMXKYnmc5TxSd+Kb85Gz5i6fdWTOXN+rJJ/Vld
3hK45qADYfFSdNlsrdinL0bKJOd4BebUd67hZdQSO4q/qSSd2pZxP+VjrAwzBws2
jy+Th/otbkS36V8NMIXq7Px/uJI10JqoaX4kYafFK+5liqAYb1y2UfaXcihy9rGU
+sCWJWn/3yX4AhlfvLdtwTusXlY0Hv2x0/fOSZHFUaJcTCuLIlBCuCaikkWeRVKD
+FeNUEWBjd8kSgUZ1lR1lXGwAzGyRLs3Sj8C2UZbssVbyXtAtRk2IPPn8cnc2c+r
9O/5Apwhw7eEWSMLQvPuDr/DX3pMz1t5BfdEbFExFjSiYIpaiZNq5vB41JWKCVgV
nzV4C+KWlNcPLYZRS8jSqHikmE/M0fH5xkSFnirfnDiFgsUkuWKuzSuyX8/kB1PM
pHNmnqhIiSp9BYV8UHRdNHze3dXZLF8Iip19XyaUIV2KaXMLodHJJRqh4I2fCKMr
8/wkvFY20lbKka9liUc7jFwk7xSBQ5f7Ue89IuP9dJv4UnYTYMqrmJq1ZcJkYL2j
FtgT/Mhm+aQcj5yxuqc7S5BOMB8FOo7IS+G6XLQOkvd00Tv/ZOtUn1YJXgV33xlh
NWYeF3AHe+TQdnQQ/yJp3ib73628Wj/3O/iPmFoKJDPovpNIjjiqEYETrQ8vzNb+
LQonXKkRKzi3jSmufd6oRSS5BHqM2bPNWXgDSKTRTbO+19GHIMmnlN0Arq2b0eoX
ndY9b3atKxR74ByCP0e9URNcOTVl050UT+aT+nKZ4oZnwOfBUw+vgLWT7JHHZdRB
xqi65FvJw0eodOb4w/d2GSgw9JEfzRDHlELdMeQAeSEn07cFRYbRNKqCJVXNbOzn
J2nzWHV5e8NMZcPr4/XBFnIxp1wMovucIed8r9q4ULfuA0j57F5A/oLPaIzzSmh4
w+9TkYSq5EEcxjjZimrBgRjyzqDDSsQBupWiG2YVf+wgkrGa+CFCILyaGR89Zmsw
DJ9ruEZaNWy7j0Wp1+5axsTRY65dUrpp0M64NlBWmKO1maYP+1W3DBKFeaq8Ajaf
5FYdQnv7xWf022OT00fipgrsYoQGblUnUa54FfCprmlzsjAG1z9Hzk1BIXHIByiU
yVhaSyqkIiRmSCGfPtvOjmxWxVFlCp7pczDw/q8tqcMVfWMEOFT8j0Mhej6rxZEf
1KBPz6aXNz04WIfBb9a7KBzDZWb7mgVSyOwZMeCI+Z15ynVsqUnv7pPHcqPgK/i8
vTo70gmMdL0c63vM4dtzvDPjNO9HStV75ySaCpyJ/yfyfs/48kO8Hr42DqfbTGn9
8tpCEKTf1Tt5jEq9aCwXvdW+yKgvuI8YjrdlnVws0PGMqAYF1G5FBfneC7+dsjRu
+zGkiAAuVrI2xlny4M51Wo1I3vw6YxHDjILHGMLUlBX9bWMCXw5UnAaSKYD7mksg
3UMkiJx1y71eqnUyfEidT9lcXSQD4mOuH/2xFuVGtg/s1Kytrni4bQc5sYeE6mpA
IHom9WysZ7ioD0fScSTK6ZjIF+QU0PyoGd0+wcTouLhKEnblCkbMqrjsqSbS/OSE
FFC8zlBYNvejpWtm8dpmJXJFvFydP4cYAf4lPSCafasiiMUwllqoVpXEbIw8v1Et
fjhBUPjiCZiR6TIZZjdRYb4VbQfTSLS+mATyIWgufZHlRjirNZmQpgsRRwhD4E0C
LCR7i3b0Q6g8v12sJGWs+fSZ4B8mldfmAKCxXdK5CEp7LK1bbMB2HW7bm/rzj8j9
FnYxN324lJEKsHNBM7nqT4qU3c6IMK7AqndtEyXOqcoe4/wOY7jUkvwg6sx+/NKz
miJ7Ap0MTPjQL4FrSGaVptG7IPD4xeU4b+Yzz50kSSwlxdc5sLBtjknzwdIp5BYg
7uJsaaVqs+VZB1rLMzW9FrQ0PKjfMeKsPJ5ZtKsNviMc9Mk7y3K2Obmh5t+puOsB
9dQIe8f4DOL5oDbVDzCUSfX+cl9ADgb6ymJIkyhPCFuhydpNEPoJDYs5rQL9M0vQ
C/BvkEKhkckvJf0Yyh+NzjpifV0WrFdzOfNwyey+a02ZBss5d6xAK2NubzIOlWrw
cWpYUIltYq6W3atLdX/9UA/4ZcOMnKwa6lDDBEZpdZMkV/H5JPhhxZJv0jbg2H/x
B+RMoOz1GuIDQg3qJEJbQbe6Y9NkfauAeoh+TFVCC/WAl542PdrUUrGjwmg1d2dP
fNT8zoQQf/rHdVyzLZLZfXuhzuQNeU5cj6cfeq7mu+oq7G5pg3UWoTmApxnLdfE5
/cV9QvPih7q7Ljrez9J+HMpQgwGq/pZLsgqsyQImLswhtVVr/doAKvZVBALGfPbQ
0r7CGxFQCeAHzpPySWnE+p+Uo4GjnbCRXtN76c3w+5T30wHWcU6jOXv/LAFnKLU2
iquxo4e03X/Fr2ZwlB9ixcyS1gjZVzz1HAQp+VaPvrQ57N3tLWX8h14JIGY5Yrn4
iJMctWBghPID+GEKmdyTutDWmkHwMe1cGJ6tfKk/lEjksrgmoJkDM7Ias1rOKgtK
HuE58QiDXi+FvV8zDBRA6sdhYeZ0VDrGPyc8gFFNptGWQGl9bbcmS/Zgw030BTMB
hZ4mLP1MLyysEoSZhVp8MAQQRYbzGGbN2O9HxuTRaHoAWHpW/mx3VzsRzRVrrYey
RQn4tli/M15JwfD9HejJ0KpEz4GzPQ74Wl6HrskJG+kh6i2+4IRDeI6vAbBVCW2v
ayY1ZdDvkggBQiTuCTUBVPZ82f/fxFoNYnMdH0CbBrH0LCRjD0gs6c9rK3jwZKTr
rbwUDQbkek7SvSyMBcHxQwtRTe3lmugCy7E1/pLQ7MYwnED3DeuSHh27lHASvPVA
WxHDMtnLD3/DIcWXClMHONUhsZprxSbLFE/evD8lJAfgRyYdicfrLOsH9CqjJpbj
VkB3+XtQNkvuwkcaDTUQG92oK5zrjxaBLvMIzCKkVTsN4UTuSqhvUxIUVCOip2no
sLREIQs1hTux2vsXB5Tu14fgGmqN8K9qMtt0CwWGsG/BhxBgz1JwZhgRKLlcI40A
A1sOIopVP4olQqv5U+lDsruR4b2N7MCWUX/cWj65mwltJCDHe0ad90BiziLO4eKF
noFrLV0JMYP7thNOHU2nT4AUjehqV8IS5MK0Pk3hAKwggaqzyf7ZjXSZ3sHM/xYu
Qt3lGiGNkZTbL5PRUlk1DAUdj2paeN+Ij5SCR73G/+kUXHsUmJxTxnM8nQlMf6bj
nffbLVBOH+H/Rb4IkuUfI4VLkeQctd9jejk0j+u8w571sp7VzIgCr0g1YZ9nFaZU
jpF+06hyoxGINMKF3ivQKx0Ra0y4dED/kNbtoOEDdwOHdSagpXmBaULAOhqFnFzj
RPGyOolC4GJOQgJb66hQlmn7OEZw0o0eJsCx7ikM1r72wGl7rXLxyIDgQuuzjyj1
qTGlEEU14EP2011CwxlH/GZn0pYmXAFLa2PXHa5WWcXszFHJL1WAUOY/9d9MRaY7
ZjP+YAQ5aoTNDfNZj9jDyYZcLpjgWkqhTUzkzPKelFSl6CwIXnYnvuq7ObuLA16W
3tISOLfgKJex4WEFaC934YEUSU82kym/dS74jPKkl+j6OigH4U4w/jHC1seSkOcf
RrrYZfCNhyxo1XkkFxmU1XqYgzwtO+hGaoaefHYQEu1fWPN1jgMRmoVKRQUUagr5
+uvhxLcfPFY/LUZsDw4IA3cVJ/2c9+vteyPJndCfnsN6CEcanT/c7l28LAQFSRv5
OylDmgXpXrf9S5aIwM+kj8IAO5I24sxA7ZvLjARnpxGxyEIcJ+nMkRpMyXPNQEgr
VZKeC0AYvMeEbh3GMr5qcSB8gaRD6aXdPIG8yw38/E6kTbCH5r3k4DFRg9tlg3uU
sGoaFJkoCongv1QttaAvnJsOerito9IYrAAPRA+ZYqmp4ChMp/Sige2BcYCG7KfS
73xBPB6ouGz5czWJBfP0F3axr0GtccfrX6T0P9uXWl4CKWY/zsfP9Q/87YNSNzBo
NBtXyfiwpk7uRB8LJ+ALdJLhyRex69dupmz8knFkgbeHQS5/KqTEK/gxiUsDGxzn
/7W2jmnhXYDvStIZlwmiyEDAOzZeTZ5mCsAdjm7+VJFP9MHZFrDnMz1J4XhfyBVE
UrD0sKZAypYfBBvbuHVkM7Rq0budzZ8nswU8W7TzQKs487sWZOhVxuzQV2V2ggIr
+qJlImfOHQgGljlx3wUvEm7dRWXyVEPDaO9fEZOoT50HVJikYj6gz8ZXHGjci09k
uR2dPYgP/99YMxaMmeofIIInivj/EwlpQUntTp16XOlW/tJhEGqGJZGRn6y1odlw
Q8tmXPl15emRyw9shKZcZvhFys0XlYsjILgSX+IzvvoKiIkq+ARFLkPGe2iejMv3
uumsRs0pEhpKnKc3/4egAVlVV9JzxIeuCUSEWs9Wqcte14UylW0qhAx74S0qnIoH
ffOyPGT4H5lqDJJ7X6jDqoILeBIBgU47RvgfP1/RKdqQMgxoo7U9GLWl8IqYp/KV
IYm6QVUSf4s2Nbu67HZK0/ypz+GVOCIaMN1cVkIKHPHB5RFOpgJxfxc4qIuMlZzY
GOkPsdg1ADCQZFnL2y4BI40Gk7woW4YTtToX/Wk0eUP/X7CWVb0QzFWHNgvMf/MT
JX3rEE61HHVou6VkREU/79S+2rmxYMyH9U4QiqG6WDF5XHwA4fBH6Ysz1/PHb4Xw
lV6c/i1SVLrE7xaba8+raX2m/MERD/SLDjtGz67AxFBi0HVuq00X2x3OLDEcM50l
O/TCPc5wj/T6lIsKOcZd4sbmVygORDCdizezRT+94fobkhcxrUt2gW+VSm4GtuvW
b0ttlMLxUql1ZsvwsRIge9HfeBzkDk/cFuqvxnFSUJWQEQqBjZ/d/sdCbBBSFQWl
5+mGnLJuUoZtFcyl9uUVPs45s/IKR0GYZsSGT9f9I9M1TOKTyeGC3H0tp/oknUMu
AFkKKsd7T7UtZgvXYgM3LkoiXk/oZLVulVJ9MzT95OxU/hxk6C0Qqe+hwE3UGVIq
xtyW2MFPkUf+9HWRU5S8JMGyQ4L3zIBsUD/xpfF7qs63Up9ewSNaruVYUxzlSVxK
r5nD5v/VVW+t2RXg/G2GFBpaeyjb4c+WqyhycFwPq8QDdTfa+JQ2JkTzUX5CxfZf
euOWXY+nLelKgBfJJGhMYKuYcKUCxp1QSug42iRN9Fq7+DY/Bf9uh5lx6TaJFYQE
CWlKeApygwD8nrcqGDZBgQGVp3hkVCYNJCYJm7c5blKNCADe/rM38gtgQ5GhBUYd
aQdgWwAyk1mA3PKxycVpOHQEoFDRgiLlFhC9mxoeuwHQCs+dtNLkiPENl2XI6yxI
H2ugNoj12FQaQ32eCryNGiZ83GxV7llOJ5m8YBa0QE0D65frWGRavE16Zy3KzEtA
VQuO29eJdTEqOaXseTGMXlsLTAu7v59R59RBc7YCiqyyOKLgvucJC5SA7gVOp8um
bN4GHHJw+PcyGZYY57WLGpm+gavtvq3LUNj5hePI4livJWqLFt18bMMuSnQ0C+BM
2aDczdLO0aNuMOfaxrAqAXPovHWC30KGaXH9+CY/qfBO1oW1xslmUVXk9ZXnwq7M
Exn3tRjOvUCbJEdM4OestAFY/MFH6jsOHhVjt3LNQOkhZ0h4wy3Ol9CwohflTfbh
/MzFLvfQo7NrlUeO8FEyvgiFLUbE8hZcHMjJsrGlaYahHP8Ta/aGEfVWoPxtu61w
XB0YBu4blk/CMguMtAtcw+WNF2+RXicWbzG+0mjulPMmUNjXb/9TNeM4208GSJbp
BAS1RpWEWJ1csk/VTUN8/Vm4hwOr9P7t6yjL5eTQNStByeAuVl2CfSU9EFJrlvG3
fXPFa5OE7LI12ErOTcDvzsUtPOQrbjeIHWrI82aRBo8e/I+1dXNK8Os3+RErCaP/
fvPtxNB8PjepmyD2GWnT/cTx1sNX3hOygJXfpRXaRkvLR/XqQmGxKPMxQFKjZClc
gOCCV7phb57a5DBUoeRc37UTAj3djBfRjQZZOnZ83yz9LkFjV6auqFHtOM+U9PDe
H0qLIPLFMlrBNAV8SmZMl+iOnU7zBYzDkdVqNCMKcm0dmNBqX3AwWu5SHMTgwqbF
eG2558XtfIvfMSt+lF6tXHmNVpmJWy5fnfUfydmtFl9uF8lzzV+VCJ+YinRksdaL
0l7AcObo+qXNE2DVoNr5tPRLK8t14It53yWU3c3/7NQ0RI6eY14pfQJW8hO7blb2
DNWxvbJ7tHz1ob5jwrzlOvBaUsI69/+Ay2lwBI4bamSj7/xuJzXzvCOelIVrjdsP
j499D7vPQqZDEFrGdPuRBKD+WWCSiN2gzpqA6/O90Zc1AE15cWAkfsVU8HjkUAwu
kjQ11Phk72XQUg3gLgjscWgC9SefAg160RabczECU0BhN7/SwawsyuXWaCIFhScX
RMpMyHzhGrh0ko5liuyWN3YC0VWJGMh/MUs9oF4I/LmyV0XfgZDSGGWaOqkd8mQv
YaLA/AjLGqqIh3eg9xvfmygQNwmyf7DIE6EiAUuBuAQXnmawanr7jWkyo/II61Jz
z6Q4cGxnG995YOACanzfw2UaeKwV6JWmB4lzLwKeR6Up7Fj9UJBA+W/W6Vs/aVQf
6YCqpyKTWad1nylh9wkTstCmN58yNAsRvG6NOiLRxNMa4K9bNrCTgifiYVlhbZkY
RZP6bjNdiqG2LSiBB1FMshP7phXBFTIeRjXLL1+ASzZ1/BvPGLTA7BztdJnWY+ul
D9gMoh+JbPGKHZbrL5u1daR62CRD5QPa1vUnHAn0aikiTz88lQIbxCdfjkhjFogG
fov51T61k/xzNrJo/OKbs6yq4kpkdiivtu3rUkaVSwP1HYJ4mTXTw11RJfkTRja6
kVk/f9IGiqQJwlVYV+dphoTwAm7Tjd30Gmt2qRzj9TxTGie3I3yDRyxRNXt25Q+d
/lBI28uE4Q31dGipOmAo52RH1l3G2sGxR7LvnBcNfGJShVxLNDbnbPr1vYXNyEmC
EBRvvddfnZw/JpMH3k0892pHQb1800mejZMq1He4lk5eaxoWrXD/Uc9ETfh9jGHs
xRPrxoCoXzLFy4DKgoFOqcWQdkem4KKWV3jUy7b+R5v7WT26So3UdsYzutDqJpwc
Y/x1fxzyOgWQT93nRhgq0dcoCby6NO5XQ+Cc2DgN6JFBV0EzwLYBopmBSZOw6uVZ
KCcjoq5MmeW8FjajarzeVKXiR96debdHu9+sgIAKlvxkQ4tCmLrcdcKf5+23uLat
WVDbeq1xKQxhjxQO8jhzawTcsPGQBMQWAEU7e56Q/RBSWMSZcYt8SmBMHWWutw8k
eK2pr4KvtHSBOy+7kXRRscYZ6i3PHGD/RPh94WRidePXwdwC2vTLyMaOdMb4PrjR
2LNnaQlJ2R+/1HWu3MutuOXawKbCthq2FMS1Ccz/xpZCeuv13W4XK3bBsCUjjLXW
0QCXm5r7YoeoYngxYxhuW9Rcpuwp5dQliMaQ0GqyOYBiRZajiO+E+6jKPVj3l8Qd
j8Gkm+ZrufnrQhbFUNYCSbdPtW/+sx2d/qJH1FVjhdNLY7uUsY90/PQFEdm+v7WL
8OwnJBRm+uYR1iRd6K8OgSk3X9TZklgk6hBMciSZYgrKzMTKA3G9/etouLoAt/bJ
d8dsBm8Lle4Ea08wBaanxFwbHVJB3bDhytAkmXdnnRo5unt/ZJCoy5qGyf5N8JTl
7vmmUrMxcEA2AhiWZo1o3cS+wDdwxMLed+eM0sT2f7iLHeqY5uIQ1WOggN1jQGl+
S/+09HeoRhAnGAw5xqHUoOM+ez7D0wdO7To8SkiucXkDcuhBvju1vNdFtmlo30T6
IkJkpKuyUL3pk723O0jSDN0EohKaR4+wjKFbZ6M1RJJ1oRPDGDRBcRyv3I2+Z/FL
ecLrl9XXlrruJR1MdyBoDNAfMyW8IhM7ew4lL61V4xAG4WW7/qCPWqa0yCtRRilV
neLLOapmePVt1ZMUo2Yt1AY+dWFoKBrD+SkQeXuoA0tXuSbutjcPSknWmJG5pIS7
XbmEJOkEg6bXhPIcy59001COaEgGKnvo0Enz+siWnuH73PYn/RU9k5mZ5y+AxZ1Y
iCMwaJU0pcDnQyD6JnvSubnNiPUGyoGkpMaA++5OBF+6dbSDnwgY2ejNAmKkiYzX
F40rlY1I2WVdnPF7RrbjVvL+GyOW2rDex2+5WPgiYKNYGRIF1MtGHUZAT+Ym4R73
HTru99oi7IW6EBoAXydDjnV3yvgMNcDgEjiltQXclhilh3MLkOtEL2vJ3cS/JA82
+xigP2WG4TUx1/QeTQXJyRsQ/7Jy/7R+cEvt+P0buq/zg4db1lul/+dLCGOAJQqJ
ir9lgXKKBCbUmS3dWpHu+xPVjGft3/mjCUYjCbCQ3cVs41KR6Qf0zZU+Bic88M7F
VRYFy6MXzzE9KURIt9XN2r1yGmSOsNqcFg7QtpVC3eaBOTV2JABi3Knk4FcDNz49
CQ7xlsA59S9ztLMdZzHyHCD0JGlb8KBTE9fOrnJDFJTwKXzE1ObT6cc3LZ0GLLJT
U80aP8qms9Jo2dfXG809U9pe1rliqtmoL5/Lh2necL+1ZYOxW5vER6JEtyACeJ2I
PwWRNrHeF/RVQ2l87vo1NN3hywwSWJertj3TsntJpQCr1SEIWTYasE1lSlU3IjBn
JZ4Mfwp9TgNHf6UKVWgyY7ofHp6LAnsKpYmx3kGMBR/2pFfqdL+xs7t/QfXc5auC
nfrue1rDAD+JnJkWdQvJNK1CeOeLnBWmyhjX3V1gyFOLztuLAl2hjPdiFcgXdznP
bOVvjwXbxkf6mQiJjAZ2JAgEj+n8PNfMTBUtGgwXqitj1OZ9tmn01aAtlWD5MDBK
ibGJKJk20Wz7eqq/vmEMiWw4aWgd6cWpKb3oSHIIoxB00YPvYTBsmY4NZaI9kzKc
5Mwo5LvlU+jRxWPdiYh2+xOOuJB/y2jyX8OfapqlzbgUZReWNVUfJLytXfqGzm9+
NHf9upND5ROAi1zL7lJCN9JbhiaNUfgRrknFx4UIGCpnoSmTGF7BBU76Fz2z/NW2
EoH4aokAEvXUJMPKOMPfgYOyVgdlJL0xAnTGVcFTiQhik/aUVZYIs3tmWtfmXNPn
pnf4jCJ3mqrxaEvjTNGi+R0gwAwfPGlk3SfxibuvGhe4FNOcXFGJHpVJgm/zR7tL
KWhMiAi/HvLoUL5bf4n2BHArm9FBWwhD9kd7sUcIVof3E7v+vMYYmTNlNtHBr0lW
4IdS5aly7mRxjw/AV/ZzHBBmXTyaKd8Q8VZuhC7R57Vc4sGSkJz3Nxhu4lTUcmp+
UkdXMehsbv2xyV+ZzuNieJCkMr7AYbHpbEc1yZHwER5xe5tlj5u+PhLvzWW4H05F
OVBHxnVphQ0GiuDzqdgeHgXD0gHGaVwCOcUD0A834phmV6VY/4BTpfFUh+QgjKlg
8DGTpTnM4J5PJqLJk6045U+C9YCA3dHLUHBAW15N+jNLL6y1Umz5QLbp36eiZGDv
dVm6p1DaSMP0qBzwhfcvdLgaoaYF+tHKXsgPgv/mcRpDdss7bbSbBFgolGi1AUul
P9cPqnxTCNRB7A66hjf10u8/d/42fhI87BwvztAYAH7tuPdIxEBzQ0rapRCYF5go
+qN87MUH9wIVIw+G+jtkNx2b1peUquMY93A25dIIaWU04WKHOixDZyPzmAqlWcml
PyazTZLHFR5Am+eRcigJrQkUc98+s3ZuyzPfpcaA/z7LI12aW9yi0ZQzQaoiXy72
4qEk169iGL/NWPR5FWaT6kiAt6bS2sf+yJwtt2AAEZf81UmTdqGC/Vb3w1VkMvp4
V+afiZEM/x5mPpwwRclJIP4xeK+rtDtKCCUyKgkMf5G7A78R/QRbjfDAtgL7T7gg
E/N1adrPXNO6U1n+1BzCy45JO+Hn0MKBkgl+TnO32CVC3+J00oISjVQab3kAL7Ab
yoELYsVstFDjb3l4j2Pt5PpttX11o5zZPyHXo+/gS1/JCL22j3y639KNv4INlInk
wFZkiTBpf/ad+jm/7Qc2UUlFuBwxGeD1wF9G9J4ENtGc05B7M3Wg9YPOQ3T+jzPE
ShqsMJqY5UhEQ2394+un4ROlMK4VX3mkmiL+86NpqDbXZq6cZy1R4IDwXOYMUIPI
AKomU4VO4R9QgUH8mEIo6iRMVXO1LYZQT2Z/MGitR9dAlgYigF+mA3Pg/eVKhKhe
dU2O8A+5vaU8ZqK58r6lSRRqR0rnv7OouxSlefIPB9r/iSyNAbv54cQ7jZtCIR7P
ced3GDXwA9t0jcSa5+Qy9XU0QLYW8eulsi8BqXO0Rv7tplZPvXnX0c10X0FP/1SY
b+pcMYJFUzzjOZsrjkBMeSxtArBkvo6nzUJst+Nf82lXOJnF/1U0pl/q9VcEJ6oW
7ouknUQOOlQQkCnAD6oUY8U7n9L3gv5zqX6VV4Skfn/V+VXlwoq5LKvRqxjfAy9R
s5y/La7giCNnosTfA7XWfaWUAk1OtRT7W+WSPt5kSP+zFbitmTJgrEH0nnbabl3c
EfE93tyaeUG1kdYwwsOF7jyY+9SOsCC3Faf8+DTr/A/rVbxLwxsahxqkmakZTS1+
Gownn/gex4/gfU39wcK3yVnr6NVFvKaInu7p5+5zR1yCAiGFygDmZ/EVOum/PSd9
iS3IB+vV1zBfNZo+t/jsUfZn00HIrFWYcGabAtNZOljqLFgGV7sxVP2INaZQhMb6
+Wtwn7ZHE0wU2XT9uLdvq6fpI0wPX4HNPIsG21J1R/YiUQNgs4mP9egzE8j3Njk5
kqsId/qINrfRbs5AeyL7l6OR33abWuH5tMoccVRYSerM9ODWYY/rjzCdG0+sKlpk
Vcj3ulS4YTw1aBYuvfaWrP9+RmbCHtAOQOZVwElxAAcKa0OX37URNe4b3iuC5tD0
Koy3eYdEFZbX21VtVCEmE6dDpP4XrO2bAXxUhFFDRqWrsQr33XAi3YGm8S+L926g
IrrtLUI2fJz1+1FPfByinO71RSzN5OvArv9s66fieCc4OjUUYyEqIWdCPFOHryHe
tGkpGrm95gcJP5iepYvfj0jAi0kVhONfC3lD0r9xcIeoojJEHdB2/C2Eaowllm76
Eid9feCBoEfXRcZVhh3abn4aeLN5ekvqA0iDLqT97DXfny77wJkA9zlKoHUqTHEQ
NSVha/ZC4XDDzlPUGwwIPS6PkehF91kW4Y6lLVgSlEBChvSi5vGYPulG76trH+kU
T+J/qwkXzKS2q8OcB7gWsNKnZT6o4Mb1vi22T9WwbCrNDyFoDiZ3CjZSjJ91SXUU
goRixnjWvyxB5UwA7HyIOeFdg4nrIqkq0cu2PddNzq2Cmzw74xRZvL/3TxjlSOLB
mwrkhZkRYg3drYdzBNLSvC7v/kODOdF+5E5ioyRjC4MlckIEEtwOXmxLN2J6SQ7N
Qso2ny8UbBxP5haH75zNPI41fgdWIsq5BE0fhwtn/3J2KcbhWXJ8BceJJi8s8IhA
UvWROQ4r/hKAY5ckFq1Cx4tGvYXZ7V4WKOAz9gvo+vJ32FnOQwoPhzpDW5h90uW7
lYHQ1epWEmL+Thp2JZL5ob3aSeOzk4m8zl+QyI6lCFgeu3Bb/rLhbTY0q8zstn63
DhlGqBpMC7QlkGnJa5t5hsxqFeUrDrnw1t67YllJna6+ME8iW9CRu7gUCPCcyDBG
4G3yWsC5U4/3wkr6BpZUU79EYWfQVRysP+HJnDbNxhLnORUVBFfgZuYg43XYnT++
S/KiBRbNSWBNsac0o3oiibcNs5pj7ZUJLAk1cHhZ66aTImOy4he3jjWc44bVP2Kk
tCr7VkPeG4qcbaYmJ5hDFJHwUoX1BOeI6o9oGzoGIQj0CYS5UbTF+LtSL24s4ChJ
nG9MaEipjzJsrC78g0AzKhvdLDIb7ncPgP2cRMJba2s1WqM2wFlxGVyT/tjk92O4
pyEBeNa2Jn+Vc2FX4wBCs39Kt6WrdVjZbUxByvhL+KERyH80ya1PV7SGeW/Gk0k2
6S5bOgPRNWhY6yQzLHkTYtkJpFzAGFoCOCQ0wZeZvy8Ki5Iu9Vv2ufR2iazTuMfl
IptF4eusRGi4LxHG1u1PJ6cR/l/B9UkNXCq7LU3l24shHo115iiriNnLkMGEkYeN
vYgRtFiyzewLwDRGJzx53ormUJ6PGUAD6jcHiTddSCiF+cEqY6e1SRc/oDVulGzx
/c2avcwZH+5slxeAliFUxyuRNrVTC4/CHTWn8URlH5AcMibyslq6jZ4zodb7YNmp
GuP9ew3WPxLPxopKZS6AlAEQa9TW9E/kkjkFF+MzYsfxrmC4TOjymrFKz7AI9f0K
XQ/2QWcHunUJMYglQ//WmqivpBtY6sn+Easw0ppwQ3GnDfB2cez6btZxVSQ4HJ1o
dVI9KK9CDt4TkqMyTorZkGmZQ9HfgQVFtK6jrwkvS0oi62aZp6z3KxPr2qg8zNq3
SnMIZjFg8YSTqCHcZNI4iKSk6fQS5IIThAQXd0sbboK6fKLd1EO+ag/NtHM/8fTN
eSEytfh3Z02Iu9dEXmVOKEiQ79FO9TltyVZYDBbfiovR73B7pQcc+qZzEI8/ACL/
hU+9EB2JT5b9TRTSYuAQQzyv7QoAFspIH9VhfhhuEtt53AyPqfwvTeUbh3CU+fEX
mZcAZ+fv1z+s4raamenTRGqUPTLcAG2+LzvwVkHR99jjcgwsngP5kB2j3ZTCb67X
O/Kx5ydgx18V6gHXvNwDGC+slONgTo+Vlug37W33V7L1oYPQhewCrOlnYovB7n+L
Cyg2UVVFpymsMr88hJBUBMjGJh9oUcHNhUiE84Onkq6vSiMGqpDu3kn6zzpvZK7m
cPZ19B8kpk5dN0lNDSi68K9mywrTCB6tyhL9k/oDSOGoxgU+hit8HE153Wc92bX1
nPcecLloeYMhh+JZ5xG+SxIXiUEXWhYfJxUtSQK1jePpgB9h4wXL2fCpeab+ut3E
vl0Z/bVUkxjUZjL8kjCaaHcGD3cepkWHy4yiLbyVWar2I7OIqUaBwx9SuJC251eo
EqyI3BDMF7RhXiF0oiHIZ3JR3iafi3n4Rzqgfh3YmeCDimhBXLX/UNo2tyr+GtL6
bPS8o4RLfvWCs7fk2KsmWvD/Kt6shV13ROma4ssTSjo=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:43 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O1sPgSzD3l6T8nTTMWk+vn7q7tf3SPKcnnnAbmUA9heV840ol8P7k0o0q9dgv1uH
MmzkmQEv29knQ9MSXOGs/hkzxVNcwfaN8B6KufS5HCFuADDASB/GWjkUcBQMB77+
jNmTZrWnRtvscIWEleoHZmoEDI4BtK9WohZHJsLyxmA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5552)
WGnO+SqPbMSgt2/UvX23hc97ahFmw3WSaIWubYaBHyQk1WkJRRE4eE/S5fdu2HKx
a175bc4lLGIr/UQ7iF1W5HbC8F8Ry82fNbIPkPWIyiqdBEiTHiubBvZGapjNC0ry
ZR2XzQKOLHYl1gYqtfYFHBZz3ejtMW15bNr9CBK9XkE1zA7GbrtIZylioo4kSG2C
sNK7Slc67FDmDvnvl7hMPTBIxMYI52tqqBW+EcXc57023VbyT87dUryan2ZHMcfU
/JfENhc96fLl36YZA8Ydn3lBHPgF3gfadlBcjSGs5cjSUdQXzVXn3xahRAjTH7KV
uyBq+bf85t0qq0hHHobiPB7Jo2/9xn53QEXienGxMg4ss8kwB0SYgst1WZq7zM3/
HB60PCL85zYpUAVg7LVrCgvudTGhmYGezBUGJ8vf5cEJMVqkkQyUtZImtpJE8DU8
As70SGKzLz/1TC1uVsQo5msSQeP08XKyVGyfh/IN3aOPO6BsRIxo4ZBn2XoeTU26
0nMqRWt/JaqZ/8ZhfWEht1FoWN91TduQ9pvSNfvhhGlI2mcl56aF5tEqGkfw4Up/
ufXmbBw4+N79kQyoarabgm1SAsi89KUPWVsBxceMJU983I+cg5f7mwfTnAl8Xcvm
JstpCOuQep86oBYG5ot9A8s6per/Kauj4yXKTp+HVhrQNmAew+Z/JP8R/HBCGHte
ZKNFuPZOxVPAkdVU2e64D/zHnYGK3+3No2ftQ3HEjmdD6JcJIRAOuT2zfPZwxn2L
QZFJAcS6vGN9cs0iF/Qe+os89nmpe7Z1ceJw8ooJQUVml8iUgrJIn75RxyneWN2S
S5AwfASmQ1HUan/+I6nfbRI7SIsejTQSpH2kTBecDqjw7terIM/d87tZDacNUHIh
S6inXboy9DLCPYwJqqAA/mkbgpmkQtjSghyYheqjIuXZ5pOx1mrpm53ITOuwaeAN
PAgZ+60C7JfWmXeymoZLuJkElAcNOvSA4VCK53JwM1MB14zLghwja/nmLfCeUB23
7HkD4R1/68LGbYX7jgMg/tM7C0M/Sw3ahcBXW3nnuwDQvZy4VxdasSsN9M15+9bg
RgjtFprjiI7cY51qY7it2hT9VNblGXFmyV2Uq0EBZKsAkk5hpYzr3jlBhIP3+Qnq
B4SVZO2vXNyJotdkDg7uxcyKcdOlENiv5+/AADjKx7hKuH37F0LnOo5I2EgU11n/
sGXNnMkCMX49gMOsbGZHQXMyJC1Boq9W1pDRKnP+E9FAcFY/tTmIizc/4btPVWQn
cZ8KEnsDRMA4NeWk0l8x1hdttPge5c19vV3DdWq7k5cbR5MafmVkNIy5syfzTr9n
A1H5P3QbOyaqe8c/Bc1nzIIoxJLZjs7u+D6a5QwXKL393g1LhAb//AQ9Gs4aDxZK
du+gec0gVTmB8IJltrVdPo/kNk1+p/SRkUh93Fww3nCpUDN7arbZlfaZb0CnvZ8e
Z6MSK3S2WaAGHNDVcGxoYeinNqZzY6iPOOjEGxsBBOip9pVwpe5fedN+naAIjX9z
3E8e+aIZr7SvblBQHr3ISUk5zD+JvB2Fx+iFXwvAhK7eZRp4SUl7TiCILoxQeEHX
ZrB4co0GGjTs2JrQuOyUJPuMnE0I3KELoAJaVkH+GKgiPeynxa0GdMDTH1rZRjYw
1Nbp54rLenZWa2osEmsKLejWooj/OYlJ1xt1ie0XOXxCngf37M2+27B9nwXSMLI5
+1ihGBZ2vVqD1sQ3K4WK32ymAFP1ghHKobXwtjYgxcbPpAJOnRK2AfIjl4w3fAFk
sLE5rkCXw8wJ/Ii7lYQ9vQgdg0OavzmUjqjMPSutDI/a3z4OXatVQBnmcS8GHugW
5fz026+/1jUhLYbamsrMneeOjUT2zlSZqWsfxIcSsGQNuSaOoxfwP0mUgDAfViXh
8anAbkLVvFcNyQ3GfKkqVP447ueP38rTTEMBMkIwG9LkQg2wuYZn+NGJOEKj2gSS
wyZbAmEysGrwH4MWeapM5r1+sRRgcgPcFQpbgDv2cl5UHUf7dRmwxjRPja+n2QoF
IoI6ARkwEE8LegOvoS+hdKJCAATXoOjNtZhNed0uVYEpRG60fhz94vme1uF9f5eE
srLlnDLUGNLY0FvlaK6os/yjJLR90yNimrCyn8AFm4EDOD9wcBKzgR2embqv3yBl
ODpLBWLP1j4Q8KNrcLo+8kOdT1vH3zdrfT+9yLddyeMW6m8KAfyklWxj0kJG4NdT
ORSzDpPeYs5dRIjuFV3cxl4LuDDebdQAym2fXuAtRmPWPi42ITmRyxKPrasTYFuL
ppP4H6/6mpr9H3+mdx2ewYt1uhxwBwVUdUOiUT57pYBPdCUOOxsJEoqEehJmAPfI
E63sAE0cTXElRzsEp4lt4gAo9rfxbsztMNDv97enALU2mzgTBKLzMzWfHpG7Bl5x
R4M31Lh4neltoQijYMZe/pLMCCp96nfQMLk6N/7St5Rn0aqlt5Lks3Or7J9yOhJ2
d0smy5RflCVdi/NFrHa3oTk6zwdBfDAZxQLqn+MT7xPk45XZayhzZfS6JeJYTKMl
WRueh8wWFeCHN9UK7J7W8SjzunZ2t6pCDO7CgT2r3L/DS5b/QIhOADU7SypKBbUC
nB1t5R4cOIurrWfRxDF5YfPs2ZGHdrIyKmvMZ12IMZvQohkK6TUz9JkulpVQ5Fib
DiiQy7/J++ZxvvtWEGvWi4Sv+BqFMW2DV/xZys5v5V4InjQL6G3X/740cwgV1H9F
4h+O34Q9DzwV6daM4XKx47HpnuPZlNMvCMMOQMplFE6UfOI+4ymjg+L95V9C2rpf
T5YRe29T+O65CR2rn9lzTtR7fLRQgD6hDOXzrEipS6cZzorQDBlk9wsyzNbAF++z
qMBt89FeZz5EeXsUwIyjul6eoKnWvi81l+LOqiAtY8/zWqR2gy23qG6mgAGjF4tX
dwVyAh9W8wmGd5ikPWWS4JqhBe9BDgnSoruRRW3bbI135tGP6ROld96DwS1woO7j
MOt/ggj3Kxb7hpdMYp2Ev/8OAFOT4W2h45n1T3TT3I6UQJPsUqarqThPME8qi/3T
rW7UP269KyYV1ohgwDs1twA+AKvlN9hBxaoBkeO1mrs5NbqUWmRxWKtdvRXGpk23
wYWSgg6rVzhfvjQleGcXoSXYJPjBVXdClQY8luWqtIdaJbZA8VPp5PJq8Wv6Hpav
itgrC9v+E1pDPqYeupTUioTdwR1b+SiOWDeR2fF9no3CHjJLzp3UVrJEd5V2JNY7
/5ooWaYzKFoWybxnINLACAte3EOjL6Jb6JoS6bkOXDU1NtG5qGO96JVDO7D17Bxr
68dvnSMa9BpFKUVrPS4UlHdY7BppbVLIbfrOQR/QGeZpa+GBevd73/Oi2rzDr4w3
FhcdjniPAZCxbjFyQ4adY5ILjl7k5djS+twRekejJmafQejOBV8Dr9Jv4L2bAidp
1gCvba5rJ8emDjrm6VbxSukEJaf0XBXJGMNbjiFLmPFFEGqBJVNcMwgL65N2mOsW
SgLzt8+Bqu3+tt+GrnGDmhIt6ITiuaHYOPQlAxQ3Y6dc6FBToCcWQ6CWLi2/3UkR
eiY1TePAKOoaxSKbhD7daKtA1Ww8/DwgtpJSF7WJivTb/qGiO0mH90C5LFHwjHeS
d5f2gnP+rOLFhPwaqzf5cMNJEiLX1oC5sodRAC5c1tEr+WuMKVl7FVU+4JNUcMoh
nu/tYnPwHW5ECb8ylZX6GNcwzgsApSCrM5SM46EMLn5D0HXNKzM4ntVR+qExrA7t
YSkcohUl1HuuHxg4creavMjQ/Bk6IaIaphdz8td8l6569/lq1PbiAkibwnNbNVt9
zXmogosuK6p8QEhRRwyX6JmQLPzaRcHnruGa/Iiehku5YY49J0HaEEtseLsc7+N6
kz10frazrBPKgsRHe7HYEvQj7OJsAG94IqsabSJTBIfv3Fl4ZFvoYFY4YSBShytL
NnevdUqx3k71pDfyxFXSpXpk1VIQDDXj+2D0NQLq1fxkUI06QScT/BJr9CS9nmv/
HNMXtB56JD31Fn3z6JAtuN7uwzhXTe5XVFnMhBUqxHfk/kt12+iiVr07jG5Sb3wa
2zE9hKrLECsbK+eyoEg7YrieC9lfXyvydqBy9EnHqho32KbouSB/jCXN8f/t3xhU
kLvlC7CPOodT1fsw9o1HRdtMG534b+70JrhO2k52V2iW5QitlnFbw3/eX31nwh3y
2PZwJb9sBF2rB63JFb8To7Q4QPvmLBc6ZtDr+Nrs8wfalAh2dPAp14HDz8EnH4Kr
F2riRKtIuGrN+PchMXUzFQQK7k/OPlaMg9cBJ34beW55P0faMZc124ZzRHRnVQh/
nZ5QpbBW4GBg/P3xMqLY0C63/jikssCwsFjP44vbORRUxbGjjGx9fWVos+7o46RI
6PAgkVwr8tmArNCnrLC7mFOrG0FpBfgVVYue4KE/8loe54oX+S+cLyN8rXs6/M+n
khmRMcGpHOiFEdP4PKTB104AbPewYEJkC+Oxp0OnSI0GgXc0Y6PwpKYO0Oj4UvZz
sjSCPHT4UY/aw5+aSqmsga24LrwOhFjRD7eFULBYADdH3CubPi85iyAP8bQOp1ES
J+/12mfimH5U3dvxKI/10udilPhsQ1+/Mkj7YSJ1LZkQP5om/aYnrySV7ikmT6al
CRqYvCUmZpKXxS8AywcYEiprQYKVNGtICeMnDuRSYw9kNca2OA5cMyWmo1QLrec/
kyLnYFicXT19hbCC03rPlprUW7nckXVFKMEuF/K8lIesJPKzBFRsFC9kCmLlepwa
1Nm8n+Z/EI0xjYZJ8utUyj2FVFDE7bw7A3ErRu6ySMLkKXhTakpjcDYKrrv1mU0Z
qb6hlwaEyq2nvx/G27cDEqLUiXb00wFKzX6Hb8eymWXDeB1/zapDbdj6zscb/mMx
GKhK0l4W4XKNyYYmsWj7aqdfc81Kgz5L5Bbj/Z2eZtYnaPBsr1VrUSaxlwpH92e8
fmHZYXkyP/w+NhC2yBklPDogoST4Jf7gJIi6zndi1xYozsGW7wbAq8yXrOBW/KtE
TEKBvgcOvJuzTaBt6slhOc9O8PrCrO9L/a5cql83ykyH4si9Rwu6Z4JBzoXZeWPw
RYFRVjnQQ9DPHfvWh5WPcknAxjzM5cbR0hN9y5Rl2Lf1WbnS1pBc4GWjiB9wWs86
wR6ArRseBleXf63pNPKGIq6C6WJZvGdXWpiMWyyYUc8/ZDAZNdeSv9RY7TBvshJL
GRevsWCPwoqTjSZ4kOsNFTIu7O/3p+K/peycsSRFSpYOQu5e096IYbzjr1AVAQ2X
nnRMFadRp21vjS3LgJ/MduGvz+LEhylzR0qsNrMKgHLn4fQKPIJWdI7h1SMUShs1
djcgeorVZqyBgwr7fNqUxJnaQxClx1ixcymCx6LWJ7xfd3OS0PSvvSOlltgqawO6
zxqjVLyR1U98S4t0fB5OiKX6+wDGWcKvgvxtLjXI9HubtU6qdVy/zUxZTXBH1CGP
lcWx3lSaEmtyhl37wMhRYRS0QU6ywu4EFHkvu1DY0vlh+1iUgj1yPiRWkhhR0jgF
oKlIFH9crLRGHY6vY5yGzLOVNw7cAXaFSa+Wiafyd0ZZ86OU7cnBI6KeZbkNLFHu
Afpt1FASXq3Gau+6Z+FzLf4d9WOaUarh8V8zu2Cowq08OrKynd+bibm1pIvvSLjN
BAoyyp8jj+6k1ANYBPRPq+EIfEBKkaSoHsIhMS5WBIZIKMFEvaksi7VDAJ8JMlua
mUWRF8W06KZZxBmTYwZvn0oADMOmZ13Z9mOcQ3ulSghEWUwYb7n/lonisKrAA1CP
ily6Iyae+alKrA6z4a6xyFd/geCnj7eXyjZuCW6YGlwFsUNmu5wQw5i8FZ+NN3oE
iALrsFPldQdwluq2ZpU36hu+tRQz7bgGfzhyH5+yLKkkpqy9mrTRDCknGl4JIB4Q
//HURm69Me78vpUj3gZzGKzquX3R3S1tpfPkKC9sTGQxXYwpRRjtdCgHubcMKsdo
g/w2RtpKKVxFjswsJX2h0tN/g+qTyF8Q/WI1dS4pulj4P0zvJXIyagSp1luQzS2Z
lIW+gpEO7zKwq8BQcLB4z9pK5sTVcHsWxT6ccpt3KaSPYx1xLYXOrZH3WQrlZvKb
CCqMjGS/l3OvtwMZvFvSfaAdc2Exwj1A5zbFObkDPlz/fx2F1ZznyKB3rTSLe3xx
LlZVxaCRXQ7flAAao6c++g7oitC/uBA9JweP1AAl9hEvLAYY/GCcAWl8/IW6EBAr
3PaI61TPYL/qiw3nKvCa7rYBs8aggPHdIMzCkzUACpvzT49n2oP3WJmhjsAFdIS0
CGmpc1ZFUjANcsB/068945YSkdc8PEkXB8AEUOdrB/hRYfC1kq410XCM6iWW7BOo
t9aoz97LjUfG9xSLo+dfVYsxTx8AdZj4g+MpjDw5LkVZrlf9UT2kvaqNG/uDTi6B
rHfLGB7vaa0btclAb/hvNagrVfmugV97WyR7kHA9vk5x3yAMErEya+UIooB6UaaK
Wi0OIjcuFwCrq16ip7/9pm+UU3lPtJ9sWd1MtJBIQU8anrIfdnYGGQWGnc9TzgOm
LwIYXzWYWhlVIcTO7EwFpCUxOamBCP2IGDo29qgpZe94T522rvqoNVFbDR7uDmrh
zfXx+VikttH/SrfdLKZYadq2LZGVGpMdnsVxNc6ugaiyjGsrgFQ6yop9l9RSI0rA
XrwuSF6FaSJlMx6Yz5ATq5Gc0IW+tIUpVMJxYwAyNFiKifkQ+Mq48L5RLkXLESW5
8USUkSQ4gks6z1VWjkCaNr/JTvUdD+M1Do0fhyFgnhsEggFFIk/UaU7yBtptnZ7F
xR4ZXIhivMH7YSH9GAR45aYtQkQvGB24PpfdeXvN/e9/oCZheOe2r+4t0d9IZV+o
ATeE3VmzvudOsjL1R+Zk2kzqFgMzqYPn05Iwe3uQdmdWM2TanzHShMf8NT5gYWeB
VRs6sFORQxnoHPgRjpUkmPq34JxsXhqzNSq4cG1vBCc+7aVZN8h7BXPJlTbLl3Ak
FFgHVucVxTKA+YWunOpDd/tAZV6MgaMI5AaKuuVBmaswnSBNFWmnHVjAQqvuIl/d
7SBRfR9YpeeKY5x2tibPqyUKdQkdrW6+1sHc4kT3lW2KhMcUSKowWc2dEz/b7BUW
MTYy5V/qJhZHKiPhvnqPsy+Pci1016IhKOQi/GB9a/OPjffLh5typxspXNoEyV4h
NUYU427EEhcGHc5EWf84STKTR6mEOeS6DnRF3c/xszWL6uAcz/QnYbF/7gXXuL6X
tf+Ov3flYnxpPCP3Mqa0INB98CNxDvJLgYzVUWtN7mz8ZQppyjP5f4YgDvoLhFhQ
vQQx7q1vPvQh3yROrXzhm6L1KS5///ulckWRUfEmMpI=
`pragma protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO��@���	��m���SC���{R�e�T��Na�:K��֕%<Qk�o\ѯ8�Y����ˣD[��b*�z}���I��i���D���L�||��0&n'&=`AT�����֛����w��R�$�R)l���k`�jH�`+}�w
݂`fo�8�	=C���=���3ޠ���`�3	���+iD׿#d6�?�yQ�:��a��*I��^�V ����H�3j��oQ,px�Pq����s�NIQZǗ��^#�������x4S����AkແE�QQ1ڹ�4�x:�6
�6��*�MbI#�e���V�l5#nE�rU)H�{�r��&l��
Eְ�m�!ѭ.�3Fp�րPx=k��Y��<���^�7S�:E]\}c�
��=�l�����
_���Q���Wvc�����ܪ��x4�P�v�����&���E%�6���G1��`�{������(��X���,у3N	�+�|n���؀E��˓��+�,��LH�D��DogU)I����}�k�&3�(�z���r6.�},�6�$�#�b���e-<�}*C%��{�/cn'D��m�	<^IJVR���HN^9H��J�-w!���K*%@�:>���f����9T��2�Մ��8��B]��1���P@aHWO�|�'֝�	7+*��o"�5]B��.��y��\�#�t���
�c}�,0�1�f����[I��a����EZ���������o,z�{��@Z��_�t/c/��7Gr��EW��%6#�Z�K�t�w�8�ܼRXi	#��&[8�IZ��
ZݘWi�P���bΕ��!E���<�h�8���Y#7���$^)os|Hp�-��(���(?���?���[Ns�����z��T>S��3����)�,C��F�lf�TU���B2<q���d!]G��	�P����O�������T����DL$���W�WiU܃=x;�'�i�af6�Vka���ZH��:��\KL��;VU5���5��N7m��Ɉ���
���}���<q����I��GH%�5�A^���0�GL������Fm?<w��K�����u��';�x[ά���
Ϥh~���w�(������'H���[�5Y6ۘ�JJw�Q�ul6'�$���P�A<�-n�	��m�jÑ ��/�w$ �\���z�T@��q��Y]���ە��\���,Ru��Ds�'��k�==Z��:f�}����}v��:���½��![��3�s !��F���(����z������{L�ŞR��!��m����J�$��1�d�+`W)��mUM8���ۋ�uf�\ȶ�:\�?ֽ�XMW l����|VP�r�ׁ��v{�j��B3r�᧪�!%Q_kCު�_�M���I�R�.I�W�/�M��I���w�J�B�w�&��wֹ~��g�ࡀ��L]�Ne����g��E{D!w����K#՞-�����5;e���dY���PkAؠr�e��2��n<T
�x_\֛�W	0�>��BH�H��z�0��(��2�m55j��a��@�*_Xq7�-}@��P��E���='�g���V�D�7�I�u��j��;���k@��
@d����D X-�����W2�"��\� �4"1Ln��'��T|�a�� Ġr!�Fɯ�� �eL>&հp�����y��V
y���|�!���[��;�I6䧧X�=Y���%M�#D��	8UYd��{�!-,�&W'F�*|D �Y2��?��R��@�l��2�%0@7Nn� 6����Q��AS<z���R������aQ~GT�U��X8��ϓg�Fo{\���{~ڊ+y���'5k1���ڗ#�C�	���*���]��IEj1x&��#&(E�PB=���S��R`�}����d1Yk�L�Z��z�����/���7�~G����I�g��[�y����*�˕g����o��0��LE4�Ĺ���R�,:�3���#t�A��:�d���	�G�����].� +Q�o���QK��%�ܿ+,`cY��*MRyج�9�:��Y�ҭ<ivJ ���'~·���M��[�J�1J�˴I��#�ͭIk0q�a*#5�\�3�Tq�@��M��?7�����.a���Ȍ# q�VˍJ��-��;A��?el���EG��_ժ�Y��Eh/��b^P�)U��@.��f�b�2*Ҁ�f����u���9bx	7�C�?����������v�K\tD���m��6�9SڣY` ��;G{c��OZ�k�D��R�z�<+�w
��͠�j6�-K;uK=j���"���Z��PՃ��9G��#^F#�9�k�	S}��2�x@���,�;�P.�M���A���N!C�$�%ec���$�鋟��eKHB��䊺S�v����*#� T�3om<�ɻ���۸�<O�ZuK65�g���Y����),��*�U�b��q��c~��V��eoDo)wm�%����<��'녔�'�b�~B�`*R��tꢖ��p�M?�.-�D�����'$�R��M/e#y̹ު�ͺ6<Dm�j:dFX��58�$�y��7�+����ۂ�_[-�г�N���"FX�H�w+�v(� ��8�J�V��N�w\X�a�t@J�lj���.�k~�Q����.���%�"7���о͞��
Q�Z�|%R��	T�uK
1㍻��K�����֤|�-�񚤵�u!<!��	`�!��U�M�4	���
&<>��c�E¦p�W5ⴞ/e�7��7�G�g���z��(O��Ѝd)f��s�BҐB��|Ӎ�g@���~��zq��|�漄h�/ɉV!�EsK@պ[�؉r���Jh�ڳ�e'�^$ŕ�Dd����LO�k�%~�u�޺���]��Bs4��r�2�\��+8�J�kJ�?R^[���2NP��-�Z���Kژ����w:�Y�c�f�޳��u�
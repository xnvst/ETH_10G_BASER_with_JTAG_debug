// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:34 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z5tJfYfSdgpyaNuc0rhbRGU+Syhdd4mfej9EYyx4AS3Av8BUv+inpgplruhB5mjj
xoZBvF8zuIQzTaqgqoMp55YUPjc8iKW/iP4iwM0hR1c6Ro+QBekcWcdGzOjOQ8nB
6QYGUByDgP3H8jJJ9g3yPkUFC3RvHhuW+r3VcHf7Erc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18496)
1KXVNVfGusEkhsmUOH1RtuWOYwc+FPUUhHvjadMAj9zaEgglC+SRUqKeUDUmAtOJ
R4zRuauhM2EdioaNtROUtRH7J8HCE+WN68JHT+xauspY0vi19/U+iirhkeI6fV4k
8H83PoZw/kEgrOREh5aZhWx1IaSCzRQzdO+DKvJKpY/aXdUQrhNXpYtmQ4Pj4/NW
ERkzEA2Ow1FFuoI+Qnylg8FHegH4PCcHWrrv2hFYQA4uJJ41ykIjHWOLVNYud07k
slYsF3meruXEJ06bXJ8K5/k5DWgOZHqR7d7TiUfp4+0X6DCgCjURCB2j3fppU8Oh
YFjXLkRFWIpVfiBFnrauqlpJ1Od0gXCpNNQpDsv5PNO73LfqL6b0wkS0ECrH3kfn
i43ZOHHP9XfRg4ki9f2BToBZjwOdB/rytIt0XfhJKQjvZ6SbODxfUV9eW36xAROq
kfkERGPeQFtZc/rAgR69Oa2ZdohL/PhACqGSYskVhIUHstNm8VBOtH5GZwcAN01i
VuZG2GPGjHpRGH3YXZWzvIPPpRShYWRtjuXIVlQdnJhFo22YpstTY6nMYlDyDfiu
Mnnmj5p24zT8vRIkTyM9rZjX/Ej41KwmI80yw1wsiSB8t7v3RAcEmlG9F8ZVE+vz
TaxK2kT0t0LTLMecxI4ntFc6weujqNzX1KOVVVDB90g4ZAle9Kd+MNdOIPy+Hvb1
lGQrZwrzpbCx19Pac2DTJh3YDm4cmwXxxeFVYiemLF2ZovyOTQRUrBKiiM3Ha7q9
BcMMOP9Li18YQJxw0IxG3szdep0Gm947GUmXvfAWsHS/XYRX1fQodRzGWWv3q0bO
jKwJHlUqfOJLTiCPzkIXtRwsfAicvilTbR2e4Tl+o/DWGPnQXTeHGw/en3d14DW+
jPWCnd1cm6z4p32g+6ZYCVS4QnbntIK1uGIOYjYVq2495njRbp5TAmXTVMmVJjMU
/Nn9wkeMM4uj1WRnvKWLTtURSz5t78og5289pbpHNZf0MGGm20Q6K1EGLnxcPP1N
tWZKG02Q/mGS1J2oxOfq/9lfTTBNSsFmSp9FZ/7Jtq39faxHDX1ivJJr3Tltu7GB
qBMA3ZrOgkhfMr5e56FLLKoYHpzL+C02LVJkawSQlp11/wGAuMQlvgvALlDcGOIf
PWUUhlNtsEbF3cBtmODQA1xcpEa93NzLinBSOjX6gJlaJVS/dIwwCixtrDWKtu9U
1lbXwIJvYk228proY9DcY2A3E3w7c0yfcyzLIFgQ+//u0cbJuYGraF8jgFyO7hvg
XC9G5JH5k8sTdn52NkvABNE8mINE1SoVK4dK70MyCSr4WGymiF033sOzhDR938tG
BGAmF15zGFEnHOPI9yISkBBrHZ7c//woHntUbMRNMrY7Ad3I+czWBUd78VZDrp68
0jpJb/RaT3NVlN0Si3WG6DU2K4GESZdQuInOiiuvCyrw+XcpW0uKxt+65JD0Qgq2
9lBBsBkR8HT1oD9ImxGtwTpAh1VV2vtqesa1Ezaa2aESYwZYkCMY4K4ueDXk/bvy
ToY2FnpbBN/uwyGxJ8DPUh77mE1Zh1HRA6TcHl7pOuv7RLZz4thXodpWVqDMD5gS
f5NEbwgX/XHID7BfIPh2kRvf3TaWs/O0tAvgiiIrKKbU0YEW04Ls3t7CBcgtzEvZ
uFjM3UV11b3OkTZsMAlBz0ayqjIGuaVDCG9GOHOsbl2rWXY63jLqvk0r+uG9KQ5E
dnXs4Vdg4IZM1lZVABZIZhp+VIYnjhCoYMiaFPz7srJnL1811huW7671KWukcRJJ
t3MtR5KWw/xNHZKUVjge/FqbXyTE38LK3FB8jGYcbQIhvhl0cmcjMa3hroR7YSco
Ki/hQkL9c78Q+4aI03UQ+xlK/g/FtceJCyBgwgFAZzDvbf0pizvnKl1+YcD+10sf
1kOJnGBFk4qtVI6SArJ9Wq2gUKlbGa/didQ+vXkT1W8gVrMcYGg1YKpwGIm8NJ/E
dJ01H0o7bvSxX92IiMxoIwh62bzS+YYL0RLMQRfKmKb7sO1CIRhj7BuzvxId2xPV
boi/v0sRX/mP9/gAcqwyOpZGIANipy3o2Kl4iLt/v1etIy48hh3uVByZdQRUuk2U
Xl+Tb+QTsbA+DOFA0yofxKzgLr4MVxW4lKAQoNr/CLgR9+ZvCdtBK3XJlogGhyhZ
+RheQlrw2WR8GfNlud1X+pLwbv0AqhlEeA7jmiYvwQ+eUMbgTdTIuYp3mhHNT/VK
53Sit8Mce3ZXBB5YA5ELgUMwGWCTJ0Q9cLrbi6wq+PT3JlajkWgbyIgJjK3Uu6JZ
DnqTvE7Ur7wiRoZbAakRtzT7zYfQ8pkCLU9kIC4QpbT6cAxxdDAxJFpeysmNT6HE
J0GLTnzPLAiazuvyHAh8Vjf1WpL1JZqpsws5phfb5RUz1cfBujw3A24Pe2fviXYB
4d9pRNw0qosp6FFesvgELaHu/P7nsXyfXrtO5qGKs7TH/TvQJvEbFnY/SoOusWFm
ixrQbBxQnwiCee2lWsWxYCnF2tbe9sXTX22DFRFSUWShrymMcVcT0AiYybLuvJPr
rrEA7Isnncg6sr6v+UQ9XmkLGIM9bHF4u2ghbeERr/7qzJEMadojGoFJKcHJKow5
huNfi8hGUEvCkWAcfRDPk6ZHl/D9R5rS7HNO9nrYFjIkQ869aaD5PQ3vkZNttftU
jmt+rkTzbcJEQQmHNvuqITA7mnDfMEdieixAjxNMqyfo3v5dGgYRKytByHBOq5Kg
hOa6JFhh0vn4DrkeDcJX4cCCp/3z6CB4vtXX/nko18spBOLwaYYH22gRKHMuDJkE
NBMBKuQCL8Q2f0baSLg0FS6XGFIs0ByhRPVPJI9ftuFyi0NJ3NlsFRWNow3Z2BTH
mDRWK9/DSWV3twwzANYjm90jqJMzQsnQYg3ObrM348xLasFfU26uBZkRnoUoUIUD
ZrDsin7hMwqq6H2FNkUfIMPyFRhfIOTOqGN31UI39uMVYrPQ25e+q7r5jKKpZFFP
QTPxFkdnmhEmOtmm2Pauy4LAGXjfUvAIxrj+QVOlARsqvog+cSEocDbIvbTnC4wZ
/Ig+jk6kr/mr2lujIdqWb5Ow2b+KyNlOuLO6wt6LwuMCl46TK91vNYOdFDvwkxnI
FpDYGstf3nVbJ4DOlJlgKu3TqmidpC5R3hHfnHDIoV6qsrmrbkbguBgM7ku4tww9
hRE11/1JqAwGrwpjMzGiJ2ThEpGKEeNKNa1kB5s/n22HABtYJr9H2TShAmHTaa6y
forJk8CB8lji73yP8jXs31UJ2fwca0U+l4Az7S6vUFJZ9fTzln0tUV8aRz0n/8p+
YItG5V9SZcTdcLjhf/4rZ3cwVxs1J8QtG0i6O3PS4y8I1sSO1E2rAkAEeSR08FbY
z/gMS9AaZqWn56SlLNn+PixYW++6rCinLwzXAVTQ8ZTfb32pKMpNjbTWPyPNVVdl
AsLbd3HKdZg5are4ZB0Ug+wOTOMjNc9WqewWQz6EbBHwThaU+hnt2mOUgaLQVait
EW0nQT3dbFzVkQpTwye4OAfh4KyKas8kPmYTIrxNr36kVLO+DzWotb/ADzpp6lnv
CR3NrjqN4hpQpQkNhGYUpJGBQheIj3GDHac+h2zTCk2B7NSfP+X/OcFez+++8Zqi
gFoN5VOqqcG/SzQjvDNaQsJS/ilHBXWbNAeldQeZzK7EMdMTrd1vzKM54Qk8OpUP
12eVgYvkd6jtju3QDHRU6KutS4Rrf9z1Tkf8WaKWOLEx6MmSzSRTd0e54EuJJj+i
mAKNcfITzwE/5ffRzt7mDyCeN8m1HBJFcnhEUwndt9WhuRfBK0FWLt1AvD2b5RjR
eRm+nBTuJm69azNv+JnhOOa8cyUn/4dGcosvbTVEjZaD9p/P1hJc4rsqQiNiZbM/
bcVMna9gOcOuLkPUL6QKpScADFPdXOqUtc+NzIM/Y31WotBrixHAOvYXsYZatox+
ZzEJ9cHfy+h3yxTjweoNFnvn7BEgGbHyaIrMKJuPYAE7f9ALSrb+jiP0WeF+Gxp9
M/9nqHJ3L+szuygnHczVfzjqJ1/3m6jxM3JHR0/3fK0eVLXhREMopdoV0qM9/kKB
Tykh9p5VaicAqyXwRLPG+nw4CoTE5rPdGJHdJXh59Uz8jvD8+nW56j7OgYspC3VE
WmfeyJSVLtYQnlhiwmKyHU5lQH6Dw7xFJqMjtxque8OIUKa3tD73LEP9k3mVo01M
VxShE4z55QdwMD8FLDYxHcuJeenwJ2rH8e+/PVu2oHG3h60tNNufxufdLilnl6/t
li/uOlcMeva9pDPWbE+zCInznttDvBV2hihYPlt4SckMWhWhPquccZ35ZblpSky7
UsWaGETiqQBjO7v7gd9LsrpelVDO83jrrEk5zOaRCuQh75S2jkLv3OY7B9GfUzAJ
tuGpVyDodDD5a0bUAFB0RHYmPzizQfjJ7Delx0bLoQGWdv0ez9A85EPaAdONJxse
xkEDWW692lnvYzvTPpcOp0KvAYRyKNGncwyw1qzJ2GdR05GN3k34fXa9WgEd6IcB
DZV0xGGPXTAsKI4tH5PiNSdCJxxdkdwn6SfCS+Tl2WQc8i1ga5IQ47bPov/Yzuz9
fA9WQhQpGuaCAHAcS1U8+o5Rz6/m8hRdlvB7N9qm33TJdGJlw9X+yZl1DSzdylu0
x8B4k2ZbwlRt2gnR28HyJYX8VY4cqxTB/zi5YoBdss4OJoX2h5iAUCFpLlXIRxZQ
FWKoAxI/0rDZOkrkvhTS9Ydl5/q+lB6ImwgAFZj3gJoQ48ccl4ZNHK9bv4t4E6yC
W8DPLCYYyMlwBghZEpZzVN0csOIieHyvzmuZ9/Q1xSi4y9TmgjU9VZe+4uObaMjB
ItokIh9ZEjBuReHdmSDHnAZ18bNnH+gg5CpKut3b8slzy/ItPuVj8auK6r4Cgtww
awGvYOJtejavNcbXOhqPQbsDjn00WakV4hZpf/Dh8KRFPHNLWXc/OAsS5+G4frPk
xJ5+iNEcnQ+GSjimmyrR6f4LZry3BIeVCf/TnPSBqfUjg2iq1oRBju1N+XEqnEVy
rKdfDkrnatavNcEOQOE/eBs3t+8RBjD1dbwVVxXWjl7LyhA1kYWTHSTFHhoh7AZL
IiAl1GaXvgtD/QYGsMwiXpwJYl8+o37gWkVHBHqC1BdddsYSiprlyW+57fcXzKcw
M+OvtvlfRidEhNZtmM7SkItvQvdASecTyCwZxzZQLzJiaVNjCLQuf3clEWSoSSPX
tXH7NWobALLKT+BfL19+0rnRbo1UQdAzVYOpm9qZ4yf+zlCN/A3hJPIRYgSbdHqf
hBcb4uHfeFWtZStnXdYm/B1b688DyTDzWW5W9pZGrBAR/TKpQsRL6S43BRMw37yt
fMnj+2JZmgP/4XHjC2XEZ/iFiBRyCWRNMyB8oEbD1MJz33UH++Jwmh/UtotCe9/Z
7D+niJ0ksz/9M1IL2UXcT/3rPUG+bx/lNaI9rXJ9PeLRSTnvnGJMGrXsCNNG/bw8
Qve0T7n8WUtKq8lIlA4LHTJrQP7Lx/9+Bv6xlgFdrntQWso3YpkbxZf5pKb0x673
0qNbZzdduFj8cRqhbsV/O49tzyRXVO+tKpIW/VvCLEO8PNslF73J1CfygCxkiP3E
lBfFScF08MAsczr1L8Zh+8eNZRLKy7z2s30CqukW8w+BREjmVK+ZXJaEb7ZEmOka
c0dH5oijVQty0JFmUXsUWUitift3Jt4t9l15SIBKDzLVNKRqqos99cm4iGxMJ1Qp
Ei1RoVJJVpXretYMwNmRwOckR0Y2ojzpAkiQcGRG08qqvezgg30f21vnyE2hFoes
9VaUdUk+qfOGmGOCVBUGg+bxwuL9XwA3zMImzEV/smRrs3o79NBDK/vD/8zb49jz
8g3MGG6ryz2rCsh0wXE0/wJwr0eoqYmLTU5L0fIwSv0cuztir56nI+531kCiBgbU
Wv698Vrrn35i9+7KdFQOepv/BZt4QekXrYpLM4EvVh+7tPl7Phr94ZLwOUfWOPwJ
1SDbv6XmimivXV4vVmYu/usdNHODf8spFVcXK6Fhd7g/FBu7N6nwApwMPOuKaSzj
UeINpMYnycqJRMvj3oKN2QJrUMcCmG+bpYELo9w0zJy52d2sGY7w6/fkew9pNuA7
KOUt1ZvIcRZXaD1n/sePihTrzGQ5RLnvhKajhQjjGAm0ql88ghbNO//RrZZziQ1Q
wrQrAdL/wFPONkquV1pq9vKLYCCVqnuTks5weu+/Cu9NilTUN0P1GHodtbjs7qD4
n3X/v1ZgB7KeOV09p8Hjn9MCjoBNZQVP148LDWTai01G4BgDFrj+cVpBdVQPAQUq
/gSETPVCJVAAwo/NCEplC+brb1am1/4yjeqhillfIH3PKSADNcZKHQS+B4dfelSh
NZVGP0R3g0kc5Oa5PNnfHEsYALvxrcyZazKaLKc1Qg+daS5gRTTJtF7w9zSG+ysG
X6wdqZE9HGqZIPGfnxTzWNMmFa69BerIP6pV2Lp+j6+1s+KzRAil1poids1xHUma
GcuWWVDzOYm6tYSOwcf1MHyKum5WvAaE73IZfadIQjJVVubNIW8DC63KQJqTqisu
ZvzpiHfcFzhN6BRJO7oIkZ2pxPq3WUH65Q/GOFW6iMkeLuoZtBVIgx2MhzQxmX2Z
mVBXJZMcjBoYQ2BsEadJ87NMshtLXgz4D+3MgpEGQaj0OmTEWpqTvPFxlbI0cgUa
eZEDwAoiyvjtAzo6SoHOTGmUGa0g8xjU7uN+IcIN2X2Yo0rpkvnYSMzzGbT8RYtZ
5zBhRa4XFvypNwfrsUap/cqCScNCQenm+YBvuUXy6B9AoKaxFEXmhrZGwunOX2Bz
g8A+nTtj5ZeRG5yBfAgl9ls+rHPUXgU52Dt9b0tnu5e5Rp6738vhpS2M4cioReV4
xDhkZJR5hr5chemR6Ufe9p4S0UPd8lWaG8x2+p65tsw1Lf40GzBEMh7OhAVBzIUL
s4kmKqDu9qASMueuuDYp7LKCENvmYeZ+eMDlvEOjHRAvzbdi9Ro1oR0ewW0bKDgD
w47kN5M0VJZAFF1S3gIEdeMoQv3gOiyZEJYkY6gKvp4Dz9sMZYzztBOJuaVqYeiK
Pzr9hVmAfHjEz9CQiA4B6NlwLSqOflNCe/IyxWSCRiKVobxCcSTXm3tpscbzQFur
rWv0jWj6WpjyNgTbc+ouZgAp9+rNDspUaIE0qZNNHh19SigK6YAV384deNJdfki1
+0ZeNPEPy+adLvYALpU1HVg4idMXwg5129my8x9a1CUlPDu2NHxx/EwJu3FZzJ2H
EBZC8MCIpLDWXykxAoycuxlJimzaeL8mpAQvWZnwhW6hhPQ7akv9x5EBXYemNIqb
8hwl0GSLsFiqnf7aZ/YnQPL/uDdrg+zkNqK3yl/ey5so29M30mMYkzmWT55MXGIi
qDV2pAwPdqLkefzfqrUdjZ7vhOSGfXHyyPp6DB32wub7i2rBbY5LWZmtxlOq62rp
Wqpn60L04mEcyklj/0oFjwNWeNxI0KtI64+nPzgimFs+p5sk00pVKRnnlAeZQGOO
XnIV4kBJkL89PCchZvK4hKJSwEgW8JZJGXMBGn+3ksfq2Ob7FXOCxL6sVljExMJ9
+72GIlCn0Msm2SLv7fK8awoE8bpsV4DTEEMVSzYooWV4YsaKTUozh30/F4yG4fCb
VyDCFCZkpF97T7a11YWGNP0ZDwb7iYZR/lX5n6bvY24SudjSSSyODn9Mn8OAPuz9
7+CUw6un2XNUrgmY7f01LnHLJlbVCyKWC/ZS7SEa4Qt7oy3iYil44EHP1cAqNwT1
8a8K+G1VeNJES0aAzovgEJXE9BHpNn30cGhwWiYIFjU7s5ZSj/BbUmtUEne8xer3
zKhr0JnhRtzPg+Lnj3A+VJPBeqidOI4QkYrVJF3bMnxaJ3cTNI8UqfWP60sN71Bq
B5u40HV8qJwY3A0yGrXuX0f5Pae14VslaHm4/TzUkL2to+oHXZu3BczrERpqbGYW
N2BFdFyi11k+ap4C/TFIYAJ2bdMQGl09mwZSZk94Po6vSGphka+e1zmJ+ADQugfv
YKyoM+aN9/9aoJh2NPXIXNb9RM8RjruRNZWQc4uKIax0VTP0N2TJ+edpHG/pKnaS
QC8P+ABMyREKDwR24nSEzgB8BLDjqUR4V8Sdm7AuVpDEdzhzKwqMAutT3xpq6P5m
wqpMJ/hiA0kMYJF9vtIgHj6E7CT0u7JMCpRSFgNDLVgdOApe+fNuLAV7HZKKKb+h
0vJBqzonvmWVB2uDrqcNi8O4fvkyDHJ8pLEV4NzYCM1D4YM/nTq3V3gl/Z5iIeiK
bLo9K6kfDiA/J1FPnDGqJLAP5Fhh0WOZBTFY3E2MlV6TQ4jO0LLvKHVUvRNEm7xu
+rHVmMvTPgs1xCydrpClP4VDCAcARNE8Y4rwV3rqWCqxJ8QxGKHZ1lpkTprGw5ZH
3EZB7HpufJa58CSwZ9BfhNS3yMhGCWeNnUe1IS04COa5vCbeXX+e3u24b4qYMi5o
Qtp9eNi84syLmIg0LEBOz7F9vHtjm+TR4pgnB0uKz5A70SC4ecfTghoHTuByYg20
IN96zr+xQVSJbUGp5JndoVDW//heVRU5VHHGfVk94rThCOYYwkHs1auZXGkt5a7w
EMTmAhreqdu7BGdlbPNHvACL64+de1dmx+AYnDY65AyWcO8Hl/t8jURnK3EyQaGI
koYI49riSYUtdj0hTn5Q9SmGAhk/ihJX9d0fadX5g7gXtk0JeVvYbObKJuVDUPkx
JmErqrQ/RyKnHDIWDKF/lqWsvdJgldmbDDkOsMFVym8qiOR6x4b6MTU6TxIg4FdO
qI2/zYWk468WPGWCzpWBXWSV5CHIJK5Ca8L+R+/TBWSnHarrJ9OU53c2xMBGb0+y
amcsqUTW+vdmqSP0z8be48dYOyJTtLf+29cgpasj3h5KuX2HZRprVVoasXlHBZn4
eKYpLLjROW7s+E2NzOQC4wFrX27RTiMKLB2eTAxsJv5yjkRQ7R1+j2n2+6CNZOEC
94O3NolJTdECYhIpjjqiJz7sV0uj+LI4pcDM1DGRdHca/oJK0tljFMnleZ12jc0s
zuy5DhzGLRODLzDczISallwJk2G0agdRhgqiDspccR/x1ppbQCZ/FEwin3VS7OGi
ib2Bu44+WmwEQH17mLOuuA2CESSwWzI4LvqXNSNGCT2FQQ6dfeIH2IWdd5s+PeuC
P3ct7Enqc5G9pRvmC9rU+ZaIXS9lYUm6jZTEA2+ccuHMjd1+D74yIf0pzN6W4Nnb
7l/n4w5QMDqwPal3aZMsR5UIBWzyCwUzs5fWMrPBJ4KppgCD3HnbilCdjzn0iqjY
/2GsG5n+LLGPLYKDbMrIb9PkWNBgCaSuEaH0+CQx3ghtDHK79duBCajnNoByZGes
KKjg/zBUbwaR9l6ltmQomF2oTO/8XIx2SjihFmh9OPslMMIIUWc2t4F3W/Y2iCp/
iIOBudnFMSSoXfIknE0YNieOHFrT54UvE0BeQgsgUo0wUidto5BNpadL1S1LjJye
sNbqdkNfam4XZfgEzQczMhFMJJNwYSnl53UqW1YC2LuhHX13d2yiVyBmzVtsTC1/
McfcjjxKYsHtW6EN31H3F0yyM5wWaoXlawwv3HK/94QdjARGjtWxtJiXvMeLch4K
P35QtV8ZSnmcS/ci3qKIC9KTedCvcCeoD8Ezbg1P+Y2+K0fXR6+hqKtWH0FvXp9Z
3twy/EUmV5HXGnxx9gaY2IAMmH3EKiI6F5covFjpMF+seFE2Jsh3Gs2TsP5S9xkn
uwr98R06zoZ9l/EWaBzyYXdJqKHGNW8wxYw2+uTUFeN3eo4RDfcJbjb8L+H+WGrs
6TL56Jbbeqm6blttmLmRejaF3tdAxRGgT9DrHMPc+hbNTYJy3XFQwZ7DaUkNlNyo
S9Pbns+p6WNCapyz4zdg8++43cBivTjSM4Hag5kU/rRGdygrfS38UCZNAFEc6r2A
G0SDIh++HwAS6FPqb5IcWw5lTPoE6btBdUvQFxLHtwKki+QE/eTr/VSgZ5ppUHd2
3MWu12ZYbiK1VIK7kpiUcuikdVROEOdafUqWvM1BqbWwExekxhMdi862OANmsh6Y
wT+JG06vvfcDgXLNWCYu//d+KpPQ5jdX3ARuGQ8E5whDBX2Gl5gmKbIf7Msm8UI4
HTMzS1k2ozpqtOXJEGHgaHdbXKoYkBBhAJQZxQ0YMMcBR+e17r4lfrleEfB5j7BG
gUthAzWAvUdW9fk209ZeYwJ1qAvDEE9+CmnqUUeO5h4pi2LumooLL2umXWSZmIb6
u41DxEedWVM4DuIcoREbXdZH0WS3mWXXy0dVa4qh5L0fQb245lSpEwnmWPU6iGOv
lHSmaHuBXBU9RmqT29tzxUYjPlQKcm6j4YBrvaJNsBXf2pqHkefKmUiFK2n3154p
k/26DfqSV3CvjLHGDDk3mRrhMyCKxV2wHQ9lyi1O0lfblHKHLoafdr6ZYTvKwNju
WUNkZXhF9/EhZgJPeyc1uvVEoV8bS4bUyXRwKf7RULuR49Pc0zPhin+NB7qUEO19
DXdIAGUURup2wjLoZ4wFRO5307nLQMTNnvtYUp+NNXipej/vXAqCkMmbRcWKkuKA
vmlAiTXARTlRDav4Jg4ze97g//+1vEBigVRYK5ZPzriVMWTZHuzO48tkYaQc+Sdx
kaA63Rwr4/AfPj1L4vj/bXozVm4bmFL/I8keOwKgqkCBa3UhqGB7Vt6vLHBUbq7H
Egz0DzUgYXU2+OEegpJmt+57fCP0Tsg62vL2S/TFUbwytXP2pedzut9k81PWKXPp
536qyCuldY2m9n6Tw11tqROvFOIFG3o+shn6Dtl2gHTTusR/QyD98dVrAaOuOHJq
Epd0DV/kIM06Ukg9Y3mKFfWoGTcKzXvejYg6pPQmXY8vKBZUMd3CcctLhXcG3hBV
83MRg1aa4rYTFaAh/6EjjKkMpUcpuOvx5z8Qe0g6k6CN1/kh0cRcmeZcIGTXwzxC
7Azh6yF4f0266Yw13QED4fD0HcITDOgSePdHBN/ujhzuPdSci9Ln0xbOSOgIPkRp
7sUv3mdnMIZIc7Ri+RtmJMO5/vOMJUQ4JqUhjJAdL5X72kvc4GetyI11n9+szl0b
/ZtmIL3x1KwVvziW2x6+cbRkOFvrQDyRxb8hPjQ/Z26szVhxPyg8aOdFAfM4tqTz
/kZQbCHaEKE6parzVu9kRJE9ca+b13Jb4iZjmX9PUX655k3hRHVXHBLjOVqUsU8r
ZonCBrmUy+XqOPNdIzvkO//JrkZqyWTiSbHbJG8x3D1KUhjG23Xo+Ffjm1J7uiAS
rEm446ZMFBnP0u26+kWibqbL92+vFqYBKtBLRCV35gXyvMJQ1Ikpxsx3nd3PV3zp
CWOb5MSCR8zmFcp97xBgkHNHzJULEPZsbWqeH76kSk8TWmvNKtBozCwR0lcQdig8
Hakp79EFPpAVYXHqMcC5862hEhQDy+kd4zMdNiM+Ua3+JI213SiJj01nnDi0OFi9
B3DJtUNHuPAoSAf8e7foqzMImjzo4Z4KcYVOykIoeVeoVlN2PqfRBjE16DGnAu4t
ygnhwHOaPR3eZwiC08G4PEaBqe8LngUX8wkK9ekEZw9gmwDlWiXyLWslOJwqnF7y
LWilgl7mUOsOTmYLf1eXJ1ATQ7ML8MJIk4CBqyR3HeQWOcmy34DhOsRU5VqhpyA6
EBfp9uSFtH86Cj50UlynEVhr/YenpNR8d9aNLRTo3EBHpBQDiKYOISMzOWxscr3N
bXiin+/PcvlQ+TwHuPUKb4eVmG0fV646NahamC6kfK6dwXVrlQujATlG4E9n+P5R
K0GhEFSrYEpN+KheKbHkFMpDNGa5IprGqzWnmiYIc7apCJM61KIEIfhtGeElSoZ+
t5JxjLekFMMuutAkzTy2riopRuT2+QL5vLv9KF+V60E+AKIbei2ng7/JvsPN+5IA
3Ua1zf3koRf+H85c1uJ+r8uLJLE/YJKkJySjozLVE9OVqqPTcJXvDUrglYiigcIW
HK6WeipjtiBoG6SvWyM9BTFfJv5+mNLYL48234mtStPxZTJxbigOQ+NIcEm7mYGE
fONTQCQ8vgKHo/RdiFEL6JwYyJaHakGTpyzTaEGI5rT+B3yUgDUDgG6dkUg443H6
SqHFKQQQnmBymQRw1mFpRMUj47bpoxFbHyqNEgJ2n2wSYRBoEOOJtIhn/pRjwUIg
7r5UJK4qiP+s/LKXTAOS5+dcxFPZ7rT9R24T2d26DLMW5HkFC45VifO3p0uDdNfz
Opvul3z7QuOJBB3aEV65dm85tI699X55DlxiVv4Vng0MkGHGwRYfYrpFbg6W0ABN
/e5AMGhr2qLYFkE+mdoi+kZQ243iXghJ2ao5x0JG+L3zbWaR2tHwykpEENbNWiXZ
Nopoqvz+qg/Jr0mLj8LBUGZryZ8+Eo+ZkUjKSqxPpdCLPyUbavt8jXXb4o0DFJ8Q
WkP3eSvaObg4DGBWUv6GzDx9mHsDZ8QFkFi9lp2m5mjJmliOGCakcsDcc/SHAhM5
e0saZX/A7A/2E3JMD8rVjbwDQzeWbN50a/1UnAoz0cfs4gSyhvpJECrm/ps8MK3p
ZUe7j5nVtZ7xPrQyDqFxnw9TL+J4TAR/dTMANABP+37uDwlVuXsWpQ+VhJmlBDl4
pElqFQ+GHmlp/POiytZTsjfExljbQAp2Chesui4nhp0A+HYLMu+NeWW5fSwxoRR6
kq94FyUD43qw9Pdsv20SqyZfOafq+bq576Bz9kRMN4MN0JvsTGIKhwxwQstaEj0y
J8n4s9K6YYKWi+adHPeV8U0zXx6b76o/gKL7n44YrJgV9cPe99dcDqjMtiyrHjhK
DVoemjJO111TYhgyHSf0AIcF9AGkrZeNT9c7EhQYpERaufYgO5NdSbMgNd/W8kCh
BujcfBi6w+4l6geEZ0BlakrvFRZzvk3ZvSoVO6TKUi68gge9po0rsGRgPHmTxCXU
LBInh+mJPLr3S+BDM4Wtngc6v5BswoHeZbOomn6813NI4+UwoROGdhO7Yk00ce+X
hVHr2+zQvJREHPjzqphej041+cRpFY3xAKfEu4fG/1P33v0Fuvgh+joL8iSUwXOI
c1JWN2OfIpOE1LBdTmPylBgOsc2OFSWMyGand9RVdQQqQ01o9oYUO/vqqQY1uaUP
2Mi31dFPPHX5rsZc7e0F0sxP4qIoQWM79tmnPmrSzIBBjjKDTo4y7bbPvQO7B/S3
YezweyVFWz/CzlNaI6HwKNu07FWCZtgBd42MTBRDbOGoHoUJIpjDijGSsUnEhlJr
k7R8LtI1wDuE9QuL0F1D4eGMRTV+64RnPgbcg1x8WKZV0xirtNPufN52p2mKgNfV
1NWLXK3E3yJdKvsV4IMFGw7aqQxrEKsEGo7DJuzFBQzV640ppQpdI8LPvlyiwxyk
Gqs3X4miDi8trPQ+TvxgPQy+3ALhLs9p2ZcUUWX36ZDy8PHjbHLkKY6nCcPIch0j
mW4XgbRsYdFhyck4IPLEaGG1ANn5fR+PegNH3C6etz33UYGdQ0h1QBifeLXv3Bne
P8JwWb9djeF8E8vlTviu+ASAc2UDzjP02dNLnzKd4aIREck9XNC0+Arjm7sZLdLU
NwQzoTpo0IY3GDHG1TiZkru0zRUCvDkklN5tnISHCfWoyPmaG8ez472wTDmXQMCU
d0UdgV4GY6f6pAc8MqJK3GHJ2pRWqnEsqcJMD02w0w35bmp9ihF7nVtB9wsT65PB
nj8QDZy3ViMxVAkTSXzn8NxMrH+PARahXn0WOxvwPy2W260aL1uw867tgEMMD2IB
6Cpc2TyNSVPN5gMPo59oF8J6ueU7Gns9Jm8sYNUFEFD4f0p3tY2T36tSFfdl4QWB
2gM5FvaDr/ma0JYBtf1Oz4Xu1w5pKpZhB2XDrQtakYhhkz4Jm8BUSR1lH6rhvfTj
aGNU+76gonbRCOHhyWETT2f+u4mTL6pfV6th+fGdAuCejHPbVINtYgaWJUEs5C0b
z8ZemvPQ5qGd/iXf5qxLq3NZQoAjqIBb2wnUQEEblRnSz4+cj/iPRPo0J5kCTG9Q
I5G0LbGEalq3QWm4JbRr6NRiNA9+TesP/Zg2wD/1CLePK03Y8eJxsvy2R5CHj1ia
q0/cFxd/o2AVdmVmoTOB1yDQLPrQF72t2pmSRP5X76hcQfVnrnbMjBr26k+NUpXh
Az9+mBgNKfrWIYuKIujh16yzn1+vtV3Vld7L91uCFyyPrUOyXEUp6AZ7td8IpqNR
/SwVsuURcjz9WAgXgYcolyfSVmvdMtyqSF/xdRHQRper6Kh9gh+fzF2sQBY/nK0a
7idryatK6zxS2paIEuABAML4NuT2btCmBvy4OiiNY5r/a6PKNqulMM+/rbaYX0Bz
SRSHNeVqVwpIZV4fMEZkKUoa0Xr0dF0x355pZkekkubOioC7DmJds0v06m3VWz3p
dblpGRJO8PAe4932RZuFPOZjwZ169tg9fsOH30P+r44hg0NBiYoiGmzVzZcHcMph
kVYnD+tQ93zUBrF3mpVdmMEH4cMIuvksI9dgJtKNQtFBrKyI9ZGqMo+Xht1LKsuY
U1GqrYguSbP3XAbCRBSdhjTmtfJuP2CAAJOrEzBCUsp4upzIOSnJZBRMUslDplme
zXDkiqSTd3pzi53qw9o18xLx7ciWerQadW3t1lolDrj9/sNdpblFHc0eQ51Qfa1C
2Gt8HRWxvepoEcY+4cn87WnSuyzADpHXfl3Fqwq06l3veauIuZWjKyymaR1iOqLz
Sd3t69187SJ/H0hjVGBzUfH0hV4vv+ev+Dy43jqlTcZnwlPBxbDpOd8JAd5WMt5B
F999eJusc5bu+O/Plc9yPXuafDzbS5eUzKyTZAWxFVaGY7CRVFkpsJYnV9IMijjY
ts0hBEmYV45RqDrxRpsr2NZ3TdI0z6fu6ZrrrgySmMLoLBqAbbSHBSdK8fxNKTxq
nh567VTtK3myOaH65kDUbQYOI2eskW+EhftMWCFybkrdd6c1gIWDGikQ4GV9dZnM
+IElGoWbA4QHT9f7pyy+BMXhTb1svLe6/1ou+rsqoAPub+pMDz3zKisZngi498Lx
R9njn6tEJ7SkVnchy1EoN8cTwgrxSEf8Q0QpLOF+cxDVIm7DXssvpAITuUkFcEHc
/9e+ckarm15+78MwHySS//1ctXytqYNxje0SRmMVPbq7J2DmjraidS7P7n4rKdLz
ZpxkH83GDrgnHbz3LL72gYscYAHqCHO0l1I+enN2dGC7LVfziLlsDNKJXVAZez7u
shgtKcGS9kTDXvOO8fzAQ+yZ/JFkz3HFArOt8sBiWRyFc8sg+ilhb66q6wWYuxDp
+/x+KgoEB37rPCIQt/gpgCO2m77IEfkPyMqVxYHCiBIA0+t6VkrlVgwv/Hq6jryR
wJ1TUwMknF6quSVd3ogmKZUpoVf/wk8fBgszxAZ/PgtbCthK9W2xsoL+yjS5/sFK
UlFf8SWYOkaSuagxyuooWTrxAsCuCC1AfvF3OqgfzJoUjbvacAv56FhsG8iCZfCo
ChnxVtg/lQyH5aXKUWHnsAg8ns8az3yq+Es+vVA7dRFJ4GmB5dHTUozFj+LZO1Ui
3o0mOVkUzGmTwlzRo2d4fqLhuF10SJYo+zuFkOp5hoqEWgCvxVNw+SCVGb7AuEVT
ten9Ft7XV4xpslewZaQzP0gOG/q4xCzWeCnxYPoJ//OBrirbqDjjbkudHUifEPYS
cPyYpVs6QbB8qbsJVEVccRLC3X9AdyDR3GhFHtTyNCom4ExiLuPvhE7GOF4Jyrl1
Gp9nEvcY9KzFGhobMf1k99rMFe0+Fq7Kmh+d2cspYUXeByWwKl9Oj9cO8BKjJr0y
kHFbueqSa42hr6wHvP+D2qPkaEFG8EFWls+wy6ijeAv+pxjmGLvTHFHRrF8hM1KY
Zw+b9/P+hvU5u0H76SzxE3NoqtxgBhBodjPcRJgQ2aQYo9zCRTbTJOJ5CVvw+a81
Pljd8sZDy7CWok+DxxvN/nrLq7RK2x4hdVfP5zpm5j4Y6Ret5BAJqyuL3oblGp/p
xiRnWVXqp4DSXhOXLe4VOlYfTO6wF2yEp+DOS6twlRWb8JOPSExBRRLlBb8d8xC1
LmLHwJzKonYSYXwaQipZaRaXmioCqtUF1VvLuiNKgMMXcS/ymWEeULjYaCMLcM0G
qfpfYu8wtFv7gUjGbnr5t6EksKvrGOhC4Efu8rdEOjmtu7ANhKh6dTI74l6LFuiu
8EXqIimbUPRmhBfXubsDeIlJW2QdAictq+GlKRY56GXYHWHvYikAnpOpx4kBDfa7
BpPcPJZTrIhHeY/i1b8SBhsltqIxtGnBgaMxq9sr8FoZncwxuy9rMO0Z+gNRpiMP
R6/pVGl2iL0H78IVacnZQN+fqwp9IcqaoAiAQHASlYd+jBL0C3Ep23VUx/Q8msTu
4rVwziKWawKID8tNvA405fIz3x8xVP7MJSEL/5w27pJXJNNsQuOwgTjdzUGFQ9z4
Ett+k3IwjolUSY/lMgy7YO6WPswRXRWCktCWVb9VDsEL2jVqlDONk8n87emhX0Mq
/EyBBqm3uK7MFo1EXlxER4rCEvXSY8zebW5xqq3l6LMX4hyrOJq/mcE4dXIyAYV3
vCWIKDzrPxVWNGej8DG8hFji6+bkya027DJ2WJsrRg4k2okvCH2ZmINRb/gChxyZ
ERs8SJAnsu2Vte7vwCo4c8+O88lUhi1ZJh7FV31uawMWNoYkFn0oz8B/1iD8au58
Jg0o6YUPJukuBrFOdR1GRobA1eFWhx1ArhGr/3Q9kfcPphUI47gtIMUyEyu4z2ma
DGAUeecTNsYYc9TaOAPbxTYY0nryJjzzX+TUq0WgxDFDLoN7jz2iHZwNOw6hqSPm
g7dawSau5qtWjamu915lErE3ERTg/QpCIu/ZWZmIKhKX89Ms2zHDrCiMc2KgJV3K
MaGcY6zYK13xMyuYV5GTWSyAgc68EgtL1wzjwcl5AI05Scvejc26mCzroNCVjpMw
AD2Hsk77QML8hDEqVe+wYnXkAL6aU9o1sFHwn7FclaMG3gD2pLc7IG2CPjtnfpE9
3a/KkHzHYR7VM9fD4ZbAs06GW78oPo76WlNPe21kH6T3SclVL6WsM369WmOLpRgy
wHxu8oAnDoGsTD9HH4S0G7V7aXWYFVdYz2y1MvxtLqc0rEsuZbfQN+p2YWFpQZW8
VU6/dt8st3vlSGE+TZFoSB9WRrOvN+R7Wh2D+M9fG49fCFcvndHLQr6L/AB7Dw26
oPPhO6wXeU9/Ef4tdRz5bg5f2+Mn19h5OVTVU/TnzVoKTsgxvKeO+iTV1rQAkf7o
JV16i2o7wnWJXkJjBFNJDlfzTlncEmba46Te9N4wTVIxhAa4TIVUb+5+MHZRBMjI
WUVQmYIpVD2wvKFmZ3qR9SVt4PVlyP0RxhidOQvTzxlL/rzild3wmEUlroS38zh6
D0GyVmTtxMt0+qcNQlWnIYb1X7I+cXNYaO5hgVy9yDgsR+cIur5jBOKY0WgdLEHx
+qcVGC5Qd290ePxPr7njxYBZsiRBg+6jPpkJfKC8XCfq0O/OzUYYnBIwE7pwllzc
6YnCs0sDHcRdZpyvi+SB6B1RtuHQTJyX1PfuJnHcMY6HdAC8yx1DMdjvV0FFgQ33
pv6KTaAqf9llvV38UYn3seOjIFOBhIcIym2Dgo70OQYRpdagPNvP3L4O2ZfL6S7a
h8pkpHY68iFVXnVOOHv6/nsFkSPiQ2YgvjAtTO/FCtBrvO4qCohr653QESvEemuA
xOhgEHsKE96NC2mOIKZMsy4c8ef1pNhQiyyH/sHo7tBQJ0Bo25ekKUEmGW9h5Idg
fifBqVGVHTupPja3xYlbLrE6q7I+VvDgmHMe0i4URRR69fmCpHo6x6uxe9kxoXXe
O0bJ4PvDEmYBH4Bsj5TMj4/xDUukHMMLVkMBl3knh4Ca9IACzevco5A9LmxIFWC6
b/zNtmnR9MUsRkk/FsDlbdQb+Siv0N1oiSGsi31FqANKCpv8uF4bMrgZRdWy1gYO
rpOzaXpjE6naTGOH6NIjVoYYcZ4XeYCjZYKvW5ZnLUuVI41tZj9GYOaS5IU3rfjH
8ohzG0gy5dIWpA2uzM/758u65UKmN8vRCYoAmkzVLS2u7fU/lETgwR82nNdI15cw
OGKWxM7SM97CetyQ1R81Dv+cTZ4b6TEPHQPX8ScKywBasXw6LUetcXJWz9M7oTrl
SdixCG1DK7iJYmlREoMpTMz1gNoQ/3tdDgFKO9VH09D09L1tw5fc6+ExmniY3exL
NnOIo0WECnbaHCCcsQoTYJrewex4d3z3nDnjjR/3HD++cfgwDRHkzWeJxs214AZR
mMQIm/wHKLh+Ukz2m+PgZXcUKhhVQH/ob0VNuIrALPBUfca0YJKS9ymaqJ5861vy
B7TUL1nkehX24Y0nAByfo0DgT6O43utq4dKATYf41ezaDYJaLfdMwbcHZtuHGJlz
Z3h8d+vJPFvqHrJVK+Fc3NJAHp3hDncaOWy5jc6PhLnVAMP6LNpGrbv2C4rFs+R/
HTiwu7rGKTYggRgHsIQF5+mjnIacKE/Ckz3V9G9ZyZ11VoyENxzg7mOZ62OdOMf4
6P2eLxrjQt06HfnPzgcy8yrh2BbWgyiijdYuX9Z501ha7QKa64xlnBoPjiPNlOY0
EKuLx6uRVhCe1UMlizMab3lLb/NlqFMFgmVsz6TgkDpyRYNa8R5LldoSWsXIrjYg
cYq19fyCvnz3KxtsK5Wk1jPgEgLz1dY79ZfLueYfqZXqG9Ylsf/1Hk6uvjpIjHAH
YAm3R6Z0AegPgRyBQ6sCbbHQBn4Y9VX69TJYbpelPL/1FqCk7/bzWrJ6U7IjjA0r
rZvMq1DRPFNrNQFORywcNvPYl4L+L+4wpOFOySNTq4Ptbjfa4a/TvabMVbYp44nx
fLJnt2Mfi+SoTZ1bYW0wlv0Twc4xcL6EINkeByp/LbBUIku/zk0bd/tvEMDwQyAE
l8wCCJSo6WfRk29yXt3U2ySxbcggSp0JgLddHMn3nkAXsfCliLGq5Ta6J8AUjCbW
KZKVs5Vg5EBj7t9k54kssemG/2Iax0vppoqTdjaFHIS1cuX/DXb/oXA73eY0pLj9
uC+SwZfj2cuOqeOD4vfp3zgBEpmOixoxVBeXrInPQmGeFNmnO3vaYcuGZECK+0Jh
jvJEn/Sv/8y/i5RX6P7TdHelz27SEP1NdBWd3ufxb2D/R5ko7FHHo1tcjMR6/Vl3
2NmCVVeJ14dd8ZzCCRI+3kpifzaQgauyVOJDq1UvbpeBAnbPxKtkwhzep2aOGBm4
3qjjdq8b1dCUSh2Z1922xV6w/wfkXa8/08M+Alp8pEfzg6TSDtd1dtO8Gjr8WVgI
HULqukTtKRkpKuLAvkbfP82nM6gZK7jpegE52k1xl4VcG04bkPwwp2MmtO3gQh4L
YpTcipCpUwP9C6QnkNIyDTttxRdfOiPaNtKYk3vRnRutNx6JW7PB3zDIQVV3kn6D
IEPfVy9yH6ldQYGL9WFD2csHfzvSMIXX0VuMqhisVtobA9yEZLaMHX14Mf42enGN
vpXnKhbPGEtfTB1En5ELuUk7lxrsHwmkLH1sNxSzLyORUi5RVoxSfCk581TIvBj0
aq4KTkl455XLDR2Z0IUL4YurTXs+inFqXznJo9F4oOnXpHRp5NFfPyI71WqBn+R1
5ARJKidAnuDzGJ43xt0SpO3VTKuk01AOYqRyvpZaXKAWQvW2HQyA3qtfvTqe5Bdf
PB5rSsy2YhFYzXOV62bN2yNsHIhfLFaBUQCD1tMF62P2Il9/xyN/MZSkjiEwlQ1s
xwmxwITgjJ9YwbOWLF5pS+3YNvOZfrPGXcChlsJ3NfWA7gtgnqf/71of8qEp2ggU
LOwNwF9UDhHMg+2t6POPOACzkARxYgw1TqSeisSi/UCq9uEgw9TcjVw+mqzlKIHL
Zs7IQIpsljJ3lxlNDR4y2nDo3R8peIXnb4K81ZgyS/tsKOhldLamuYk2sZSlxegn
whNk/Gpx7gVHCtK3YR6bT1L2eUA6ZDK7g5yCwyDDS7FsHP6iUTGiStqpokbmWAyT
KE9Y8iov8qgDrtPJ9zP14MGReJsjjyU0Qm1fhZLGUjNEcJLebmFQ8YGK8Xuhp2EK
3zhMlRME60QVk9+9knAS5tp3EVwb3gOc8t3H52IUygcf7+PHn0CgJMI4o/hCslyc
gvu0diblkDmbrVY8++NulMLV4ewMaBYWaAl67Ts3CbyBoHLyj8/oI9jR/pGm94jm
97sT5BsQP8z/0Nmyo4AoOqbxxROzh9Ub2sgsW1MwEDhyonlZtsvTrtFVVbDpyJbk
3xP9+Rsxm4vNOoUZ5gmA9A4kJwt2zsNUpN1UloUGeS1PEO24GKHekZp/JJgPf4ww
UHxWA9ckdH8yft4S/mF9wrdj34d5KfjDh3Q8tEzJdzQUL4Ph5DvNgqiegmf7sT6N
Tc5pk1CQp4elPTAZC6eVEs6bOrPBnKMGTsQk870iQhmJZU4vwets6GAaw8ERax5Q
N5nv/d6vzV+wdSSTeDUqT53DRJMs/xYvTfdUg9n1FMG9Ly6UJj+o0uXzKotVzMlb
DYPa0Aikk/PBm05VJAncB2+go6MOP/DBCwgyJdeiRaiAMDQWQEGIKfZYzpQEhT92
jnZcsf+mZql/a2YDzLX+TXt7GY73KSEa4V/YhIVMpYoEfwK5nqAlwzv3ssvl+q7q
wovDngWJVyBXxKtSN1EqGGLZQdKKfoRiIh5VLpO2fZwJvlBY7dEcro++PwMEsQjn
uvP8AP3A5eakgMPIbh1kTTSi15mAGEsJAO0MeL6WjDpTRAYjSMy+WmG5oRxGcZni
24YsF00YNhdgLH1B/egsxD3LfAtCGlcOOerAmXDXu8ry5FPJ58DgxiYx1D5PdSkv
/VFcymB1O4rXTF6HoitKbmHgCvAthREgsPMZTG636mxzhN3JEzl4M/1tG3MpK1Sb
Ipy7MA3uk2A13Rhhqc+OjsFfjjnsMP85DEXLNAVwas+Zz9353LkHBGn3VHEY/kX0
NRNA4A542xVNQNi3BP6pdIkwXiU/8+pTtJH3tW+GZJwR0bpi0ynOOR3qBXI+sIeU
xfVoo14RiTikuxO2A//HZEcTnFHe5A1i9o63SFpkgK2a9TiOPJXBQS7bc23juWxF
+mZ2DQmuC2hfADCVWIqBcAaOFLdZ9rVEBln1vgPLuvB05goYGpFsYRTuxVpb6rfq
O6jeXclbUO0cY/cQh9xt6GrTmj/RD5JD/BmKdvYBwlczdHA9gECSHQudYs3u7rXm
glG7QvBymoIQw6KlAm2z6JgWw50JsmFWw16VVtg/hzD3t8ugjRymh0EdxfS4yPhZ
W4BT9wgcmrMJp7VySIhEtdqLdKOasmwCYenQYUwxLQmjEwWZtWIGuLzMIL4W4fCW
OUs0k8OViOoayYY+Sv1FEcJ7kFdy/jtqP6R2GmSNpDiYoUUdVhVgPwtOgfKXhpPD
b6TxdYjuXd/YfQP5bjdIHQ8zGsKdXedAG6hdZS8tSKqYG/IughwQFP+nefv58v8g
mrifcjleGwNPG0R6p91z3AmpLwubBUeUIJIonqE1PsL1vVqWV7d7rInadBkvapMo
HKRk5dWCPtevZ9AH2e6DUT3HDmxPv+nK27wE1kY1MMrywCtKnq3Kvnh3yBKyI9Cq
7Ov/V336karvDGHUGezu3rwK7AvzJo7bLVygncRk3Zq28FlLf30qcZCJdDl9fq15
Hi7OA6RDt71+bFNwzWI+e4k7CPKE/v62Iijk9OJqcAm01R7fQ5Dkc84hdkQFZqZC
/mJkX96yda52tXj0QsBKJ7m20PyA2BKtkKrjbX+ocF3WMg9Hj1ziUxjuH4y/BuRl
RT62+fMnalGkqXIrVhX4UjYdB7LtnJeH7g65GfrnjdNzfKfTdb9bySvt4e9FzgTo
SUbiCOtfgbPU0wSby24aHBe6P2WWktN9sMYBIeFqAyKGzVoro2budpTqwbbkAQCk
XbmlUP45F+uKI2YdqtnhjJFvO+wXdDXyQC71RkHR4yvtmVhJ/LZKvxLAwYor+glR
cX4NNxqn0uY5sguYCG+ruC7i2FO3jhjuiLhzY5Frpi+lLMWjI5q/VVHNkc8PUVVW
Gg7XDYf0KsXwZtadrs/EiQovl2POAmF+ElHUuYljT7qb9Kux2qjLuZ+S6JNc7ir5
IVcCC8M16h9KE9WKzssJB9t/68jXWlSnHjMx//yzmDhUrSDwTBY/Jc+0iFaRU0ZE
QScXrsqyEi+GW6M/5ez79NjDOanom9jZSo/J+Sp8ZN9kFgaXvfquF1SU2cY4IPU8
C7R/kakTuVAc6wtbLDHnh3Xfx16X+T4xtA+yiBDtJpZYDBb1Rf0/AQInKvKPHG6B
DLLSCCpgd4dBZZ71Fglv/SknJpD5We8sNxvr2aG1xQC9/IM1IIXgD53mSxAdWmSB
PORWCOyjmPIRqoGzj/IZ8jVJ1LM9afVnOx5i47q9Te5B+mIkMgs5CTtVR000C2FK
PJRfABvkjmHicjCavirf+jKJYi8U4TvMxddnM5YuO6xvQma/k5xcnviok8YZXGk2
E2E6cvEpmNRvadut3sePaoRMtTNXJKx4jNvPrQUNnCu9IfohZ4j78VO975BrmHJF
+ZejvsyF4FvfyY47prw0MtowDv6mViL28fFRuZOxzieQrKpT8v32EIDvSyusk2lx
TODIdW46YsFY1pl1VXiqrVbQYGe0AznWHakrczLs5OnRdF6FNC332HKek8tC5aqb
JIA4i8sQPmLPNPitaxQ7tqGxEb/PESh7lOqPmJONRqaZBHd1JAsH0hJsve7/aS8g
WiOG8CUQcnhfTu+7q6YEdUxbqoN4y+eycqTk4rrJfZzI7zxZ8e5Bz+xvxAkH26b1
zLK2Ugz4ID+wvKRyh9ECigAM6xas18n7jXjwryoBrUvey0X3Fq6FFbEgaQ71qzk/
33rxU8KSIt/p2xLxpNyaO2sI3VxoyD3ozUxMyLESPeN9PTvZWRPE+l+xHBjD0wvj
FaMtMRhGl2ZWdOh/K8To4GmyZMVFERfn/E4/Qj8PJnaL5hPrucxFhNhfFJjb942c
dbB5iJFp+6E8egYCmk6YFNYTabPky1Y8wGWenezllW+whDXFmU49xHfaWzBuUMGb
2A64x9HnWxwBEUUh4L0q+0L5kNO+7N1S79c3Py012M3zIz8weIURrMZ4nTiylqeW
CX12Tqp4pAH2Aqvf+T3GDAHRJrj4OwHyJPwk9EDN00eyYIERgxDQYY0mK1mxj+xB
a9lfumiEVR/ThXU4Xuj41HGMst2vvi2tUl5nDRMigdNGAGEjf/NyEAYQJTixx1cC
veemCDMmCOicOp2cqqUPpiQ8mAiOg/vcs9FnKioH0H9hM0GGCxbMDf7pDjz3FO99
1PyyPpSlWvL6Ti1zlZp0di61y0SopPz7qSR09N8ur0TW5zm0ndlZGS89hjhgVTmV
kQfHseQXmVAscR5AjDVkn+NfSd2zzksINzuKetuqzLmeGn11xKChkBIXYG4fcRvg
Kysfx1ET+ihC8q5mvF1IZWw0ZOfOlL5MJ98MyLQpWvxRNn5HW0TcxAyg1wlMlkOg
WdLSeDdnweHBOZpfiU2TA7iD4gluUNvqIoJnMbt/xOhPRnBrH3YtN9cuE9OTl9f+
fLMi91NV0sINl3soHDnBxPj3RO0XzdkunFTkp4f1ue1n6fXmS4Qx3xNuFg4+LAfc
sNizqXCy6007cAL//Y/zRhhNqbhQnrZbCrpEKYG1gFlIumCFIMaYy02yivcjSaH9
Ek4V+7JmEdHsiByT9ZM7cSEk8J42ZE6sIoB6U2okOU3O3owPezj+K1bJbixov496
mjIG69YtoMOdJOh+R39GH0VIIFmcVCJZWbhgb0h/I6dGc0Bnuj4P5MDt1t69Moow
oQphroX6OR4mwFZj5XF+bkxGiFw8c31fQLECpTeFBkwZsGrEqxeMY1tJKCq6xVfe
Rf7rDGBPBuxzePhNhbQ3zNcetiT1rX4Ks24kxAV/J11rb2BfjtVlUHjUPqObKcGj
MEtUuQF/C7k3rgE7w4/8FXim2922EYpG4IQ6h6O4OdrXHSdjYty0Ee/9UIICydi4
bOnze2AWOUmReVkdEkjItPquq8hyRGQvm9JxqOG9dbzb5iFQAZJ58mfwQdP/tqh8
CS12JuhvjvbEPGdI0tq/LE8m83P2iCa4ILKz/u+CYi9j18qsz6IiyHAd9Qz4sDQh
ucFKosrFFgQhpnyHUU5LN1sLCGR/saAZ9lkx7WAMTJMFMYFonrMnGsG5cDycYxiU
AuwqggEgco2rV5ol/OblKHffecZA0Vn4syuNBs2+aKMb9Dpt9bkDWL9iTOv35End
RX7BswoY88/gjIosNj0ILn2fCQYauA+9I8Feu2qXLLuX6LRjKqIGfyxjdsbFkic7
TRVcx8HdqbZ82XPIPP2ngIPzE0LDTM+fDcQW53LNsPun370xh+FmH5KR+XTyFqID
tK8VspSa3+Pl9jjO2HHZ+bt7dsuMhMrN/C4h5pf+lG9rFsHLKau8kMrfDE/sq+em
Gz5/cEV8Q9fwiHuOPZt+NI84Z0WARF36QOEfSYlzbl+089uik10HE/9fZfIQTlXz
WZvEryISW9O5FnVu4aqFrA==
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:32 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h1C0zLrw2XuZRhVQZEGiFC5BiRGcp+JHhvLtocXrNBeQc2rs5DnGxFoTEvGWFWOb
/RDpoLDg/DqBJ36tVqapYvJlElQMuCXygKDop+qTLsZLcrmBOnDNIrYMz7mAi/mE
VRo6d7F4L99M9lhkUXu0462O8sbX0dxFPdqd6wig2rA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7840)
Al7tt3FsYG3MDjTf9UaHXHE4l13j2rfbRx+fQ7vyHw6iTKQMXLKI7IKH1yoI2rme
qZwFQJ9FyQqEG77ecSFyGqCeFzz28HA+UKX4m+59J1pjYRqMhh4OKkNaqaksT/Gy
Cu/S+AZYrT0SlaVlDUnEHSf7k5sw8pa9I1ola1tUG+MlbGr9kRVDmINe1jqVempE
LNv06Ick259gKibmZ55N8AKbeZ5kdP9Evm81ggmumC4c0a6gtFRuOYXILJviG6O7
le5Rag9NZjyf1v0MGgIsEO1ykVToREeGK8Knf69ck3j4KZcN+Zf9EBYvNtBqn6m7
4bO15G+qmUl5JXS83RYxCZ9gd1DsO+oCaC1lu+JRRqePCvz1bm7Xi4vp0xCUZZfw
P8rKnAfqDzkfVB+r50KjfxnIuRI+cgx6TM3tFo592CefXmjJN1pnP/e59knwUAsb
falMoK+sd77PAyLBNJmr6o87LmQD+v0iF5tIQZcSVVhPSsuKjKwNkY4fNrGKkxw6
YQB9SD/UoRiyvQF92eNZSKDEfa5siN4vIghpMl6lUrli78YHA88D32szAbyxRETr
69PBtxu+s5e4xPlm/Eph1g41JzB5H2v5GP1h0xxfscBB1XIeU/SmABPbubQev53u
lTcxkuOXfdALAnX8m4/RVkRunGrXS88EVd0f57eest9suE1sAHWuhPEwDKiVvxBN
c7ykGkwKGDM52uH6jv1FSvGHQg55PkYXdYsAOQBloD0PiFrrJfHlThK+fIqN0vv4
xbCS2pnj5VhjvpS4435bGBkC+SgcElNzvc957uRz3A9d5VStXCo0+dHFHVKmLtAs
wucaUkOHMJ9izReMIUuEph4lXBZjUMOHBPS9VuI3r/bLe+FbtNkqEDsk3eP0O+UP
ET3c06n82vutHM4uuEtVV6TfKcQSJCG4mRbMYF4/aWwL7oU5FDxZQFoT6D4S3iO+
KIJi66nvHw4Dy4a9GFDvfwEdU51QXTi8l/87PhuQoQpdyoLd6GRuCuN+55tLjiQl
QprmR3lSUHY+4sD98LPkJFR2rZ8FNmLeJzO5tiJTkNTukwqPjbcBw9sDPmUZH3Ip
y76vzLBFUZUPmKJ1Lu7WKSgBNlU8XWadUJzTtXuzwJK18E0NwU2mikENrDfD4G1j
30RVu5agPzdh4b77yUUWs8FSH9B87lTXsKl12lAis5TvpPCXPQpDLe4n0YFtvWUX
gnkjUlFkH/DmVEC4pMpokYiOsEsjplDJxhokfOEFE3mcGWFvqIs/oBefG+h4VQj0
ZyISN1q3TRppAWxeNDR0RaV0mpZy2VY9nsCS2H7/7BCR12GdVXoZY4zkH1qyzi6l
c7wyymw4Hlojk+SIRoIzQ1TeZB5icuByB09233uYZJAwDLMnHXhN0UnPw9xPtaLz
+i1LiKHvt9ayifz2QC1wrlp0IkRFlBOJdP1hM9QhwmdpqNuwNViCWE7xiCHdj4Hw
fwuElLV27C4POz3zAUuNVB8Gaf6HQb+CM8n8G4IN2JG8H6uVINkLShOY8nmm3mh1
nagPXGpBHqNcexbQIWTbEO5a6pJ2wYnGWryi8M2bA4SWOH5jvqs3tZcvjGB720as
7WvCJkux5qjTaajAXy3ZMdCWETSMw9emDodBt7DUKpLFz64UayG/CsF5yGyrW2N8
gkOe4w6wEAxjhZ7PCyDXWws2oAvqvchgvqcdkPz5axfdaRbzK9bSWdSOKv0q+5n1
4M+yVepkZTLbtQq7CqW94CwztOHJYfup/2vewU5Kejs6/48DZAdIu4yp6Vf08oJV
xDXOrAnPox7P0O6IIxFRF7EHUphj/1ReoWdXwm/2i2awbtI1em3QpVyyii0e9ahw
PGsw0XgHsWBrIWdxpCaZQvdXkrhFE9bN18qc7ZNQDMD8iVSJ/KhPqE/Kf8iFsOrH
3Avz6HWfS6n53LEWbbAVNS8Fjiv49PHw5h3FN3ipTDgKOKfVZZNTtLt5MlW+0oaY
7FaxlNw0s23mgVumFNAb4xxp1xqfK+7u67oNBZjdZCDJs7XCXDb2dDj4Cc9FaCwg
AH6MwzylO+OFj/i8999iK2m02d7LvlpWpZAldguYoJ/GF4p73nWIfbaLiDnAlXmp
Wti02pcr2vXKCjrKY8t4CH05w1vFqq7mp26iJKfKuiYQ/pqZqMJpCirxLuxSa6jt
5Od/cDJBRO9QgJqCDXv6R7VdjugXG3BNtdvoEDanjweFA+RYZy+TCFFFAtqVHSxX
45tVrHrpSBzZZpCMwzaKgUNJwcNL2rfizuiVaj/yKMJTPsR3BV6rAZKbROckcJop
ilm9t1NrPeOoXqlJDMyicFhg1yaEJlquzPmlFKhW8Ks1lNMlbVwnOgGFQu89l3eW
vOQZvYZK6OtJUv0IwcGnAl+NgQf6zfbIDVJqlLpmkBUNu8GDiye8hgQLIT84hgJe
b3ljrIM2pkFE+zJys/AuSD9TZ7AJ+2lBZPbGzQByYqxPn+j/4C0nGv2q76IjRYEt
IvCl9xTJ7fi6MmZF24IK5CCytFvCKRSsV+Ia1i/hJyh7QGBPal2rusylv84oP0m2
mdx5fJqAUR9FRniGXyTw3APqnBQMP6A7sGzncOHf5oSZdrMu0lWHMMTQPus49fni
MJqb6o6X9dF+OU2MfnRWYaQsKrR7HgAUdvmhMDD+NIxvJldAM8mIbYLuoqoaDnRg
w+5yUu8guZy730L65UM8p5Exsl+50ZXsfIFtArGSF3DVjLf90t2olNBcorcrCVpm
RheQ5KQq7d8Oq+E4lht0wqos3EK+nPXcrm2/45fYxBXBZmFlqrxMYEd1jORFIrEy
I5cvIU6kP9EoikjB27gt0DwHALliL7YGpu82VJ56W38lcGRcI7uu2M9r0oCFwJmi
f9SfffrO6Dy5zzRIS5KaTzcq0c+EM7KX+fUa1DTlztbnrFtL0WlbbdyHJ3fAAWTY
ruMflDt4OMH1quoNNzZBpUc1qMr/gdT/CBNzJPssHkO16H1LFEsFcV4CpO7ugqVY
ooVpYTjYCVooTK45epWJl91Imr4iyakkO4PbIHz68ZDrbp7Wi6OyRgKT8KNq/XUl
xGSv4sC5nxNL64EJsskXikDIx6c/psYoumNiv6Hphj7pi7ACd4gisNn9drtuI/Lg
Pi2fWC6QeU2TwF/waVjKjWwWfTGlGtFQkxYHK9yF7tnXwy1vyjsHix1KFF/mZ2tP
lBCRI4HeB6qb8tmnC3XH0gNOIYZzJZU6FZOHeVYXOjXFC/TL2qY+1fhNJR0nqjY0
yNnd3n0vp/SZjcCRI4mIqSO+WkBi6MS2EyA3cum8BaYQvHx1Dk5hQ5tQpfhJqkT+
wx3u8MdnD0WoRhtO6ZOdgXN9g3YG2Dj2KWqV13pjbammUzasuBzo+NPLukEvVO9A
a6oYVVb9lW/vCjyY/uGDooeh64Z/2xDFht7Hif/R1ANScQAFiaTIQX8ViIHa8mGL
xMsm9febXx+E3QD6xclvm92BLzCtllgdXGfVJPEXOHejsA+UcPpQlyssPQ178kQp
Tn5SSg6b6nc51CfyIZbbb4sC+9UiDYHymA4sZXHcvgi46Rg+C92pcAGEZ6jeMHzl
LQlW/4dW1+AjwH5xi1/IwD02zV6lrLafUUEyy8QDgVXpEhp9Gr3HZ+wkBhFJc8NX
fHpxo8ra6ZykONaIg93NUW0W5TSZ+BE69f99tdab2Gs9cCpyzPTWGc1snzn9SMPh
YKOjjmeMpoNSoXg6NhiRTNLqLtUNI4c+PSRS/RkhElF6kPA7BhV1/R6fy8oK1aRb
OlIvod2MxF8wsa63H1tnfOTfSG8LI+RhIHaSZh1JjGjv6ehg//CTJYqqtmC9n9lP
4BjvxVq7ObEDqn7O5lmQlMYC8jAHxVewSbKAEvGW+fL/3TBXG8x4bHwH70N1HZiu
ArFSRwF5STGNR503JTLujfAwdmQVwF+YYckxTZgfcWby7HdVGnfH8LExzln4xi+c
CUwf8PcZizzWQT0P9o8aUr5sOq/gJSM+9+kqa1osUVBCRGvPRX2yctUBODqxw+66
dz/rfHVpkT0P8qV3RNMzIiPVeSrTfFEeSysOiVolP84zVoZCjWEttoGM18zfeS7a
1jMZfXS0JEDKRZzZL5FjAE9VTvDGMkWXFs9oCqmvbm46UqOitbAZlGqTzj2nEYyb
ER+PUYLuwyW1nE1ET739/5n4FXDcWXqGWxjw958rth7dhp9AkDoPiZ1DZ6o0+fXJ
anOjuaLuVqDtbGY1VbVC+y215fOkJJh0sg7L3cSZhISDnfnj2j3cu3594uF2JIg7
reDGNk8E0/JTwBGPO99pvxd4YFMMDbAokOy+4teZIFfkIBP+CHZGX0ubroy1NB9q
DoyuA+9BZqFs7YDC6d1pbN6E/wU0ZXmH93FhojDn80ZginimulOMNvJPFyGPpgCk
i1d9qdL5LKFDXRCOjbkMx/PuPL5f649wuaOGdW2Tg9uhS4th40W10w/pI/DbSwd4
b6LkAirY/tP9l2dUaKnsNUW6X3A/LrvuEl+I/1PT4Hv7b8aBGDklpeUpOwTp+BQ5
E1DAGJ8p3dz/lWyYHICMAdr86xb9zHTbhz2tkpjHn+e/dvoxEugv2u0LPFzThlJS
cMI/iQBbJJtW48zLwf+73oGLtywz5PvSVBbCRo1Qjmzjm2xibMqcwjTJAqiGexch
1axquSHLOp7CR3fDq0MXORNK/5c3i5QAM85qRU+4FliytIFyPzcvNUE6lB4HNERo
9BXLtuHQuWB5MUurviv9o91mTgu4EXmFldS+mfgYDO/6WvrWgbT62sxUHCaUU4Zq
90CGfCJKQ34PAQhqhHsBe+YJWQhXMT4KobJAk2UE6zaE//+q2XVizhQKmGVmJh4B
9q/dPxOmY8aHbBr0hIf7gC4KqthnK+YjZVkeQFhWhDT/FS0xMxnb+SLVq75c0Cz6
vluFDOuqalWaIW7eyvUgpWHzLJmkX8X3smPlwOTzm3vTXsC5Lpm90asyd9vUh5Y0
FEWUVLdJSqqbuYi++bxDeSebcUc2X26YDRDgbiML6netwJ53RlEXzy5aTo4w2YoI
qf/IDGJ1z1alPpongOjKW9zuHnZ/hvnFRxdUNl1OhouCE+WsFWjXMzZFzo35Th7Z
BM9zREbRozn5r9d/y5gbGJAWhzqgSjHrwQDeSLID+0VzZJ/H5eSiBnZLOFMmxNfz
E9W8oELw8jUn1uxM2x0Df0+kNKWzu93gwxcexwOXgRqd7gBERhY3te2ItHK+PNhg
eygPGVDM484UQuP6x+ZjWJx5t6ptKHxPjopCqujcZv4wZaMl/iuGWt0NvdhtHy/v
/eTIslHjWumCXKvNW4X3udCCT6AU4osPFeNeAfOFUS+sO2UTKHU30gNr3wmg6kQ1
9IjnQihluyaE4MHD0Crp6ZMBoSeO7tk6A3RVdIbGBdiLa5agna5Ywmruy2RjnF30
qB+8OyY3zlldUNsaVzxUDbM/P+ACiSKIpZs14BJxg7Q9QLVVfysoby2u72CxnqMp
vn1xOe+55N9lvuFQNgGn73sLvYFAwQvCkBXK//bIYfQ4TYrBgYV6KUJY4v52CmHJ
FQ9W2/ntTZ3HLEjbCoPiNDqRMiqpE3gQ9Jc68HXa2l6p47rpEhw2c/KAuH6sszyj
rCo4ca9XR7Fo3ghY0+BFa6Zm/Lvdos9Oq9fI3P7/QrtJMhgu6hnDpN2KoKbtrjyX
XJ7jPfMMz0bf8f2+++JzlCUAwOm2AC5d7UXP61KWVuoSK8iyiew1H4ATM5Nisx0h
dw9BfaeoyTaxNV/Qyao3qM62jUOj9hNb9uTJk5GD++Z9RHcJj60uX3K3r5chiCtT
/715PFBjp8kz/WC1/nKmaMZELbF6LTAVScmwciZQfmKWnpyMniObacXAwOK7YHyT
JbQC6cHa/BYtgLTxtCF2UUmINgmqh/UltO8MLNMgrzz5lB5XrEre2V3mta8hzBAM
sD/kNUaPMjFw6iqRHPFQoaSlAnotV8JiVlB95KXkGT0Fd4OtGVWsai21MUoLD++6
Q6g//OFSxolFg5WaOHs21zIi8ica1ETyO8ytB4K2pnNh6oCSlRAVwLzh/QAm0mgj
08UaFUKDS6g6LcctK47uvm4hsBlMMBd2fEYscyZl6bxKruVRYQbFfz7KGJAFWFm6
pv1xzwycjIAqg2GLxhGBXfrSxRKLZDV2TdKTuffJCcsJZEfp/qowXfnaI3j8nNzS
hV4Hf7JLXeQ/rvVjmBFITO+v8nqfUbHXtOwlybdpDfIe02atXpQhw2FSvmDriMZ0
W9K6l+AxdLHFHtD6fQl1eq0riHQbnhKZ9YFf6THDNwxzHJXiFsrILqEo2Jl/U1XF
TQzEUFi7Kk7DfCYMwV1GKu79z5dS1UdYWu+oGfKyGfJHQ3hiowVDdKJ9meslNM3F
C0bcL8T+/5LkEpQA6mcugcrs1we1Fje7GGNWBgpORjtcLR4f7mr997PxI4CrQtvz
+RJN1zk5EDazkmXwJIt8bVzY+R36D41zzz8OK/a3jAFBwmKcv4Q4axOXbNruMWtY
a4/RmUS2qdz9zwDw2JPloWFZcMFQUpI4clbhkbCHeOMPuW0/6gLcjQniW6K479RS
TuHkuDyGK6n+9QX+wK1D6fnBO+pFHTaU40a2hGRVVFHfrlDufzWiaYDsxmlFkTqQ
cjYfhEzwgc7khZZVyp6W4uOrbEsQVn57B5CwXp2/v8Himyxh5dJoGcny609uikvu
E+1vsz7SZDRSzjs5YJfjW89TP4LThQ3nNRCOg+rTZBH0rbBNdaqKO0RD/uTZ16+M
O7mCk4pr4KpjnUhJTtaoAU78w3yVKhPNNgngHjR3hVLRL3YuUWi068C7HFL5aEEr
un8a09MePeybGwhilDGiLJSgJ5OzHwBZRfZ194kGDyUP8tw4I2u6CkYwuirezaFB
gIZxPs2tl/FmEZ+ao8NFFPG16L4uRZ9AS3mhlctQDjNIZQ7ZCGdfbVs6UbD1llwg
asXOHZnNcVH5/P2HJXyWCzoW+0DOso/MDuen0xLLnvlFLmq6bpv8/RrU/bUb+S6d
3buJMsQ6MkyVLm01Z/Om6+IXMKiIV7BVIPXI18H8LcTO2B0fBRSAAnPZhJSoU/Im
LELt/Qn/1k3A8ioqHBVxZ+jipNstkltXY3ftvk+793O+LFZepht9Uk+8ONY1Fhw7
vUPV8du7gh+xtn9C5a+jJQbu3su+ekJ7xK6BNriCFnNwT7x7hv9xAUldjCvc3dgK
AMhDYWKkXhSS3lk4C8GEgKXRno4KlirMufVqukaDREVC1uhFuxBnoZ64CcK4CmmK
aUMfVocjNEISyQKgpO8rgHjuuvG/wBq0cklLVJUfOxcVSB1pzH+9G4MDGiDpnap2
oKQkmeYJDqoyZtfXJKaVU3UvVUO8ddE9yAAQfoJOyCw/DbVn5UqW8RlARu9Zi20L
Nv7xsUqZgqZ5tDne5yU/THXCUl84wElXUpLW67Sjd7q0JMaToincYqLPT73DZ9ch
+QH6G2gequJiwFN2xTt/45zzfWmGE+KE6ZUQLa2ZUwA3rIH1HGSt/mD/oe2HBArl
yREobozFxlOO3nf0IfqwqhQMsvGFkdB2/zKycGYKRkgSGB2Bg7SgC9oaB3q/Jkxy
Hd7GqxMTt6SSjXjjFEhkv5GxOvf0uoYJ3LN8arVcstDmC7zpq9qOjvpaT1EDNjSd
AoToSYuH9Uxr9AcwMTQ/dlYJlfkASNcacT8f2L3+Z2F4Tcu23vVTFfce7fAd9Lnj
4FOxD3gTf0aOZ7Agz01UDGwzSYhQ/C9Pj+vW352cpewHMi79axMjoEbYg6mTARWy
Keyw4HoQcPNE4wQ9xQrppxUB1GyBKnSG1tjAdA6l+GNeD6kXb417wUR5GhXNVQZf
ZaEAEEJQG/cdGu3Fa85TaNzmJbGO+rWObZb6OW3gx1ZufeQQ5EbHE4rudL6uj9Zb
34rLrWV9DDF+nh0GM2l6NNs0mmqM8WUSIJZgV1Fb6dX+HtHmbHpvJsTFzPc0B8/7
/tTPIA7gYs9/eTTf9OTVJPD4j9jhYLDzt6mPuC/rz6l1n3jJX1125WVmu2xIWguT
gvRYUc4a8IlTtsUw25y0uSVjcrXlXlxb2MKLfEGKlDQOJkTTYyVNlqvzo6XUIDN8
YQbdh5SioGHtvOWH0xCOfIfjoobBpk4rXSAKrkdUqmZfLITXcFrAhNxNNz6mMnz6
oArFGxPXrthgatlSNbSkATp8Q9n9FCgijGpQBLxxMk6LeaHhSjrVq9JCAFnG5XGl
wF+ttKyUGRICVoWM5GTk0XWsxk8GQkqLzYZClQjbneJg4vfw1bm+vWrja5qgtYa5
V00HhWOrmknjvccwjrcoOK90oU5VjyOBFa/f0UEtTf2JcvcCHbbDJ6FeA1sLEnsD
kSoxInjTLo2J20WvlsaUZL50gp3bGlqK4pXO1Zglr2F8bq2m/nXC3nqxUNFAT5+n
NSQ7vIJ85SusyNRlbQ4P0s2n8xb67nQDRauyJo+/wy0Gbv8wK0B702uiHzYRwKNC
bSfcp4EOMIog9sVEXFeVE/UVD4TjS8LWcVV8gHRrkXOCe1oPAMH21Gb9N85i6tZr
lf1SxkP5nxG0QZUDCA0vIoSFg5PXBc38wFHbEYBz/JGRXC1va9z1ZKMItHTSUmfG
sb0GLZ8PkK0daHB+4cqHyHRsfQQFiDTvbjJUwavzpIdRIkrAGW3Fs4dEUwrGkBLk
Z2yyc8JXuJa4tbCXSV8/y/ywlHM+iVpEQkgVtqXMHYtWaq/lLVYIbFRE4haDCy0h
WEvmjRmc88Tf1wNdeXAaPFm7T67qQZkeKQQR9nybJBmq0pCmk+TouaM3N1vK12iD
nLKIgZO8bckZfmqejIFregFIQUNoS9vo4GujNJDRMNNIC3fZpS61TytX95nM1ZYP
jIdJ+9GlZkyD/g23hJLhUu2LqoB8WagkDaW+V2tDyk+IEd8/ECTLgeYyyD9HhJD+
fxI3iRPE02FoQHIfB6M2gh4a3KpZ34nXwErwLBIonm6Kdr18VRpnVd9YDAum6kT8
wKiq583+PDvkBzmYra89GH69m8+H/tda7DJl0Fl8x4vYFpVUfTH+i1P9rlV8fGN6
B7pRN5C1GlbCOXBkitZJDVZuQvaulPRV5+0bkpxgWKLgAWDlOpQeJLfJy315xFZJ
DY8mw0KUDyw+XgNg/qU7oF39Pyu4f6yfXfZcoTvoggm/54RYMx7Pm6cIo65PVxRB
m7RBpZsFe754dtQOulLyrZ0sFqfMjy/3pDKk6kUjAsaoGXlPZPNbhgMITNKphmMD
eWBhUdmwYc2ceREwtkYPs23Q4IyrXAxUgoLbHXh6ZOSgsDzPoYpbLww1MLBAGzJO
mBsoVNuPYzJTkxJ/GDddOKR7AL1KhFxR/RordkhNMiaqp3ui89aMeaPyqrGMjA6Y
NzubcnVcwsHb8frma8c5C/Qlvgww76DvdiLeWooVeDwsKnJqIycfWAql0Q6hBFFZ
hLtqEQaun+5hKu/mG8/EVHVX44aA613/hHY9eVoCe1ldvpy+ZJCih91ISiGjK3AU
QE0y9sc8Gi0swqm4ZT4gLfH7ckFoa7ovibinw6Gl+idcico2CHzOM5XgnvcAUCyu
kbdoPBOBkMpKNxFyQ8UVY9QAqJgaHHG6tDbswyKOuXB3JQxwE1rck5guksPTfpxP
DlGVddN9D1LqqXcKQ/hzjMt1QgOzHiTELVZh3IeUZr7rRLiHc4PQ8dSj+ATxUbfc
eE5nZo2i/SEoVgf4Skl5jyRde55ReipL1A0cixS0D14Pzsr+k/vbE2OvufRIor7e
fBUwMgTQg/I68uykxiMIt34OdgUmxd0WBdLWSCtbH6sggHJR5UsRYDdpsw275cm3
vIKI8LPNvpyOGhi0nXmjeo9zGgZ80KK54ywLMJGpe0UR+Tm2S/i8u6YRdZOVCoxN
FfEHhw+c4gT8jhIEn3CpmAORLjRClOJUHLDSpRoXlnI22WAdiMux2ffbuc3R+yVc
z4Iwx2dAmIOWI3+IFr+ZrLGRjnKxysf0EauX+no7Er92ctK4LJg3vDUc1ap36Elt
0HkdZ5fDbjNGvapgojhzlU1z9+Xt8SH+nyFuRIj3uaP+c7MzYdUtTNe5WkAss4zT
JOGFzRCuiQwCsC8oKsJvjaed8xlS6B57a3/s2LUsras7hiWAqsBcxmbDnejlSCdw
hNTZUNHKE8qbYF+5ZRIT3FDvqTOTBzWAOMvEiLlPfP2TOmoEPjyXimmq1jFcohxa
Rla7FLbyBIoSSw7F4wDrBHKl6bWT6u2iPHG8e7iRGTx2fim2EYzRv5ft8VpnLOnW
2jPeevopFhuAvIwB7ZGDRai7L8Nh9SEjtM8Kt686R1LbVvl8B7jqnsIhQp3gSR+O
5HYbj+4n2Cz4TBzU7NwnGh8TRjN2mKzWtZOmQpSjJI/Jr10K7UxRIA9ejSMXS8Wi
VqrPxcGgfyPRVAm6Dou0zA==
`pragma protect end_protected

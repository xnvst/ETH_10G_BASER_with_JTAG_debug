// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:34 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AUsrfbs3hNt/WgkDM/kVY7jyRA8+QKMTIY73LcfeBe+ZvNXcw+Pa4iK7cmAwMPI1
IAwdGJJ2EqQtUrZktlGdNq6OSaTUpJpzHmdZigNzr7M5mLX2JbA2vU1jxfDns5dk
M06dx12G2pPSbvhPnMKGrRWOgvSD2YDkgZDwVafMrKc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8144)
S9w8slwDSxmLQOL9Ik2wXyppiTlu1OJS30XKJ1mo4t3APd3l9fUwgA2jKPnr2lTo
Lvr5F86nO+fHrKbC3at0rKBFOxsvJOWWdTiKozRl7nRicgLwWRjKh8QCchXMLBIm
JBxsBbPQ5TkDnzyz19snPGw1NGeSvzXuoevv+fH4ZsTzxvKyC+ObD4dHdsZZ5zM/
6mCKP+Q1e6lyLrvOEpqZeQzf1ve6BhCKUcKskgsD65rUffciLmtYN/kqmHmz/y8u
gGA7y106q1tk2doGRg2nuMZ38WgNWsnENQd1L4ZgsveJzoygiu8qXSZTZPI790lZ
YzcccMYuPFaBr7pbLvSwpmm2SvDAvw9Z0bOmVCsALjAtX805qDipy1nDEd0o4/bA
XH9i575lrTgKj7mQmJFv8fEs/LFU2AQJ43IkHVhK5C7C1Er/1q3Nda8PTI1dRmx3
YgQxcXxzj1XfN8Ztee3ElhUlIMw3r8rVEntJWWuSvfgYZ6ldeyVmWOt5YVcFzbZZ
DdhQZLqjffaf5o32WDLG+kFXEiIMneip+XCF64Q2Fbqh941V1YKnmLrqIWRXv90m
P0PFytj2QUH7ClNW3FL8wCWe9SItiFs0ih7f51QLfpESKhw+sNHQXGche4hvkjy8
OXXI7d3k6MEG3DubvW4TqlarOc13a4AT1Qo5cP6O8/30/2VIIDwEYBId/4Rguj4g
yEhMV5xNdMbOL71rCbTvv041NtiifSQ7EYvHkYbRHKqsmN+9WHwY7pqOrjqCwNS9
I3UUvByF1Oe49FjZC29J+fjKcHZ/t1bdNvXcBJS2TDurpujinmp5m7zmw7055Q71
yqIMdEs5koKfVyBYdIFkllps9CbCXRGWmuF6EII1/A1Ez+JUsb8L3c9uz58YeqKq
fTIeF5N1dzhpqqLn9iAJ+CjM35+6XKYm3wwn2geerEh2OoQb2jjM1IeFgBTXfRrT
6KFeXBtVHhUbaj8AKiE1ARz0TerfkTFVQiZm+8svVdfh2Pr+K4hOq8PWhnkqDHtC
tHWo9EYMkMs5DcLq5a2iTbDo33XYyVXUoUnwZKQXDMYMpYh3+iZQtQqtsm6hEeXA
CNqt+yiDrSW1TYn+kPTl8f8Gl9oVK4LKfOQFsGOabQKpiQ0RNy6CQ+Socs8I7NCX
FwbB+7RkKOSleiM7WjkGO29Dk8J/s3GLQimiGCERldKlfHMjr3CbHQAqKi0kCaI4
RJWOzAd7BoimkcvjzSlUFCLaanUkQ+cqEfJztXQGKLhl/cwA50oPUgj8rZf75IaZ
HBbv7XAg/GJo6dJNiNOGhwKOBiu/fyroGLqZb6Or2/yDTQj63WoHnVrYgGx7SvYv
v0DTnsgmy0imgkjmoOAaM1/6o70Yj+VU7Ny6vNNKz0ekb0WhsLH7LMMWFjmcuG64
fCPfbTB/tO0uahfH5vrCG4f5LYIPl/f+oz9OqpGs+MkwcspqurT13XuVRgRNgwT7
HzB2hoO2A1Qe+pthSj2skxluiR5UFVZ5+Hno15bGEL8PzBrHH+b2ky5h1WR74L/Z
uKCMX+WIWI2G8SJaYlujTk8ZvkNHGdYY7R79TcqKjJpjuPkl7NoCV5HshOsfu++L
rCCKzxwrtDIGA8zUP+9rdY9ktxhM8lCOWDDpUWj4sPMM6m6R4/2erKEmsF0LRp8f
WovNOfYYqUAOnrmCLtwGPTc5tTkqEcfI5eaGVEfNPrLs+2AKA+DmH9RJUPB12PyC
ua3QQrle4Ej6uU9hJMDti+iiUb/ZrogghL/NhzEQKy9dm6jWb7mn3uqtWXKIPEk8
6vr2IDQTb65TbrIalDpvQTtehv2OPFMQqqNkTzVe05bFu4F+IJ9tGMzftjJGL+PH
/52MCz6bqdSfkGCtuIQvslDlI6+2EY2FG+Bc7zQmq08zi8cqqftwEsSg8WgFNOoY
fx1rr8O1SZu5IPSBzL/IjRKE94Jw2pEvSV5HvCSTaIOwYNTrnbPEgcjasTk+T2i7
ZW8GIwqJX5JiTrJ7tAabxs9joeAHjBsX/CzAtrgYBjnsytHvWaVxmHCfHSKX4v5N
tXmI5DB4ZBglQ22kJyGZSH7woME3E2P7lgJGjqc9GaLrUuaAyvIp+NP97k9tNuYq
REAAY41ooE/O6wIVGfid6MkXg5jfit9WrNh2GKmniOu2PkMMuisGUGwRKo52xWCg
8xbFZLGXRQdLm3nKqAqE5fsrNnOCq44apSYpM7wGYqBvqYI5NU2D2gQOrEdd0FFv
oW5MwFUzl8n9zjzs9Z3TlhieQw9GeT4VLMXReIqbzbTGFTuK7s3xIoOtjGDywCQ4
SGdFnsFK7JF1H8ZLvjJDxEbBtgMH/CoxWw6L40NxRhJ/B5ry1xy8lCNU4A2213c+
M6ZF2y52oArA7MidQaQ/FxCywcdrWT6hVXNpTgA8NuckHxhB2TY0j9zW7qZG67Db
4V0mOKdA4AqP7Orv/KJEwxtpDTImNKlTQUFPzL2fdmmVOjOEQgdnFYpvIHPSY3qB
tmyEvrlv59/+aqvZbyJk9dnUa/i+/+kWg8W4ntbWLTzsTynCSjkMbXIKJoRPBsl8
Vzp/fJX88LRN2MequznE4N8AvjJ84cTUJBNMH7x76Ax1LTc/2bXaRau0lXrLLijB
HU1q8mQfIcuJG2Z28z05mSfJ88oBcr5SFY/OMftbb2/raGCFZqhTIJso+0Hmdgby
p1+CIy/UE0nKXqOZJzTe/5thtw/jnI68QVaCt8onC46fwSwSAdKlrs4bSfNG8soc
GLmu1RNos57xDMO/sdg0rG0C/4KZKcD/IU8QlcnymIZtoEyz60cp8RtJ3YWXlAOc
5qrEpiFOv1h5jsmwPKusr62IpnC847WkJSOh2TxbHWJGbj/CCBEo3j/wHZIIjMd7
z8j7xwEi3kvtGbECoZBCHtuKewXEGU80JvaOujvTrNxj4PZiH22c3Ti0bnryKYT5
Ttqx3EaX1Es8kJpGsGvrZnoGqrm5ps7uUisxRlw5N1sr552EOUPROboMbQI4HlF/
r+kjjhHnhexTc5b8EJ5J7uHWq4CVmDbRBUeIQn0/wDmj+f6C4EH3EhoYgM6ZtPYO
VTA36t6ttRrHx+eYyo27Suz8pebOCWWr1XnEC1Jyzt/cDT5SzzONZaBAo7L55w4Z
WziJyjTqAy1WVbPVXDxSPYEJqsDJjKYBWEe6DQyzFDuLJdBN7GMES3bG2qvLoY4U
WI9FFcA3Es0EveHqStvmFjcm/VpB4kzXuYYxVpIpD8UhCmT/0ZWhYz8k6c6iBcJG
V82CGFsLogIIjelLBRSoCm/tpymNfQjFhu1gFUmPlSro1hsfR5vA8Mezz6HcoFgR
vBFLjnC8vcknFWyyAZ/GthtZLsQiq22Ybxzho/J4kFuUR8qJPJ46DPoPxB0/ZDnj
/Rg/Ei1otY5kJR34GSxdVCBTVpuzq6NVa8vYC2dl28Ri8IACI5W/DgdAG7Xvh4h2
Vh74LuCEhs1cSKCLsMIqYS6KuI00V/+FoRWIslKarkncTxk2jIhRHg78gGAPaPQi
H7UJ70C8mWWvwW+oJbMhVsTg5y2gFyN9ZylDgAARtUrjU0LSRSAJEbStMaJ1ULy2
drPuWp5Kedg5a9PNc7ofsB5nl49Rz+g7DdeJJte2BhgRzBFHBv4cYQ8kztI8xRni
CE7i/hhPxczdxSqw/wdTSijDLptIHD6GjMI9l7H62p2O3O7ALJvYWyA+BmnjvJSD
A/iQz5kuxMpv/S+rTSUDqjqcGmKlD+ZQ6jvoWhbf9h/pNw109RoidltKSzF2Rzsr
Vs1FXfvV5jJdEtVDvM0GhjYuRJOZ7NxCOTfI1SkLhqsSiy8cJHYlfNxEFlFzlGZa
m4cPH2PLj/mqA2289DKUTdJU16s8KgHXKi4vyVGz6DsPf41ysoE6UK+2RC5V/yMV
n1A/R/iCT3jqno+LBmzuFA8X8JZWBYGM8ZZEVbWPSRMISyiAnBQ7GeGSyFHIp2gt
MNewiS1CTOm6QaF+sSZBqNr0hefS6VgWHY99QCUk+w1UPVHLSwcjuT0+aykHXrS6
PmJPUtbm2rAgos5R6nA/iKhjtIOpJZIbn4frwLPPZgL4p+DO2JXgroKFIU/rxew/
CIMoePAKByJJd9srZSPl3XChE7eaSe+c/dTbblF2YPjxQYHTpsmYw8KTbAqDxGDX
VtNQyJWu18ebyw0FAwO7f7Buzgp75cCuDQh8KwEd37zBDI/aTbZT/nYWll2Wa1js
Esn12N0TfLu6Iitif1aKK/PYpG6V24WQoYW69SVrMdkq0eb/c2dVdJkcer1wiCbT
jut1Veb0tmqVb+nBjk41Gs6FfpeEFsfJOKxHoUhOHJJRyihpsW3b8AzBMyPB2823
w9m67+0aNOIAwky6uVN5ffCyXC227Kipva00e7ttRe5LVLb50zXoI+WuQOPAn78H
frA/gxoo+VhPqeedkrvw80jc7eLMoitu8xWHBLSQHrKE5s5oRkVNTuHsx77McATD
9ZCUfxOcooNmwlP5PaBPRtOxeitmg9eZKIpYzwNHqN8Ws7TAsH2jHYfmp23FGSea
ylYuLqryrBM+g8QDxbcTvjAj6ijcGfyM1dO8vBHDWViDgLd7Apn3vGRPdxy4brpZ
MdVURKOTcycIPQNhZzLxz+URMsXTggTNTySbh5a4euyfx3xKtbIeHUT/iU87D3h1
LIPhlHqkWR7V4G9sVceapK+YHlnSEiRV6DTdDO/IieEJWsxcXKpb5VqCqmyhFqGT
p1PDhPyj/ETv7qMpM/KyHUbQmTf62qH+Nixe/nZCYEWHLanY9I37+2ljtJaGWjlF
+sBGnngJH6lz9K+ihoqtMVFV/9LxtiiKOkMENT5kT/8ekp+WPIMz9JLdjjC//H15
ovP+htMo56SgQTzAmiklnSW+Qs3oDt+JPyRGKEhjE1wrntNk3pWh4D8NINtGYDmw
EgbSE0PeSNf9tdtkIFVLVfvX822vao+78Uzl5E8Y5wrMDUpUvasL0fmM5fTv5rq+
YJzVMbJNuXq45r3VTgjnxOsLcJSEHsrmmWAaFS0fFS8CHldMbbPj9t6AeKRMEVI+
rivp/1SiHqqcgjo/ObPDGb4HTSSqG/G3nr3f/CTG2Rfxv5exUOCir7mIkxg5X3Ty
V1qH7s3JvgTV9mM1cPQMloQyFwum3u71o7DSorFsv+F7vlJN/DZZPLNSb9uHlTqQ
3oLSCnuRybO2OHudL90ceCbQvvZ3QlUUSVg9YbHEdxsSiBW+TWmrFVU5cCCqVHYH
BK0542krTmuW/vNiIdNaIwhyd1DFicLDd+Li6JJJEWYIOmbr3Ee3uGn2Ai4zJ5pF
4hva1Q/6Q+Mx2HipR+YB/wC6xZ0in+af6LpO8bhw4QcEp2J1AxwWQshwGcIc/5ta
lN2xvCXhpAJ7jnKjP8nONaqsM4CgI95MiZBBI1J3O9T/0x899chxMiS9Ey07Y7tO
/2SKT9lStmuKWgrZ6gVhGebl5Af3M0s6vhq+pTJPjAzbwZrhUX/6W1Y9nnS3EB/L
MGg0NX/LA0SWi6Ys/nnnrPE5YvlOPD78P4/xX7kPJ89P2SbA4uXaTIEPFSsqyQ/F
RNzwt44zOmBLRlcwxZLY4uM4gynaRINe2uAxMfJlSz0qPusvJUp4QbMs57wsYxVc
z0MYFp5T8PneBse84eQulqf868rKZOqPq5PIDFpew/l2Jc+/pzCYQxmrv8Ddai5f
3nsZng0lVhRULudTs1UneDsFaow6b3XLp+0sovyf4RNNn3BIgD0/4PTEYQKwbg2P
e/roYaHxY/bZQK8EzR2W17Qj5Dd/Zj0r1FdU7zxeF9QNWYeFZNrzpiSzOiGUsMUG
ySyL3PV+zTTWSjFPyKt/7RM9duC0W6n4CuSP/uHFgif3kNCCOvPRSN5fBKcqj+kF
NsTRRs4ty30OW5BcqTPfFVKDor1XTwl4kE6vZGkpOPW+WRW1hF/UioRsRU5XeD+s
Vc0DU3WaqHje8j4aP4A88uMFtvL/mGLmEoFbdi1P0fVzH0iaSRxpi+KQzZC2tJus
wDcqPmkd+2yw/9g5lGyzeaZ97TuJoTxq5ZrkyxnoEQBB/ocVdO/kP30dAUbdg5PX
LR8zBqBaB0rYo5fzJBsavMoEIi5LkrCOKT3k4Xra2FMPQlA7nq79083fUwpjo0/y
zSUKn/SW++8wFeYo4DtsYL/a9GG/IaRKBmecDJXkiO1xUcNel/0cb2okKcnBeVlP
Ch9KVhUMvmbzHz7qHTnB92LA2eYZaCuMur7Zgd5jszUdTqON+tHaNXGfiLwUIYVi
vyF+L004e3coVxtXo1OZ8bgZ0JVBwY73bfymthPwIjDcwfzjXBht56r2aWbZTiBG
vaVPusOTgxDRgL6xTKHjL1bue+xTCTvDKtFC9K8A6/EMNxW02OrErfpSpdDclE4+
N61faVgFVwdWFec/y51a0mSAT+XTzuLhwFzRHa27O3qFqx5Ejy6EldmRe+BjnXK8
kqPikdZoZDviqt2hb/+69/MbQ5h0dFHFPs+v8tCMHtT2ypyXZ5T2UPybhmNx4b0c
kEoEI6j3+SFZPrrVuNTiUlpbPYdp5QqHheXu1NQnG7FKB54AYKAP76YmEQuALI/L
fBk9jZV7Iu7qmkARmdCzwTEOBxrvqBThN10nFTsbFg6PeU4kbZarIL0V4EBmeFI4
KkoeaujLHOxlyeIQmX1IuV9/NR2oGfRITO22Ni+HAYFygNxWvzwBIKOTLUrq8EdD
tzeUcwJxpzk3HdoB+AbYQfGJLn0s+QUzZLGsIBwj/wJ80WECt+fOAuNuI/FOZ8Ng
gncaMKlmF6NX+IrGxIZ644qDXRakOcf5//Syyg81mvUhf/E/I/l3SvK/jRITsRPX
Khww5ic72tuCZWGHqkIAEdFOXif+Qeqb8ftZX7527z4wnAOrlVGE5yUyTYBKz6bP
pTmEoRyXbvXvauIgajXRvsUSAP+PQydQB3vqHApLGZWXOLsoC61NmEl9/mZ6O5I+
yGXYc8YG2CG/dmof4bBqFUL1VfypruIq165ByV9aaIYNSOSN7s8QjiOIos2bySZq
x4ybaObHU7YBzjrHrT5azvgT907F0WA8b0PpuhknadC/UjvAc+15o9Or2IK678Ng
7IgXN0Jz6ZJXE+h1lVDvzueSUfRx20vL2mvNoEgS4Q5lSb/eVmfIrLgpswhdoHaX
ZU9OZaLG7xPZfumV/htfJzwG1yzPv0lKtcArIXcSKhyyz8HPfZzZaa3Kv78LahGz
gH6ug0iWXslBVyaFxEZWBmAEKtWXM/caYA6fB2i1C2WJTVBfFmJx8kVGqBHQrvfu
tCIFVrMHEkJWM8SmOjUdlsHsBuZcVFASwacKMn/r68bAr00zfkzQvTIDg5m3UgiW
anwcHMkt4grDjFny2ZhVuPqYPvrF4xw8CviLPCWx8mVC3j4iRVCwmKPxXBgNvR+t
YrmGIPNm8VDpHOMTl1Dm8xALm9GE1e5UZEXIL3gDWu/3yI0dzlzt3G4LIWYwVBES
yivireFl41bp326OYL3FZhfxpz64m02gpT5lmN8FFIRitzOTaUJ4QmjCIMBHu+Rk
d3WZLRsKmdhSWaRsviL86KEwaZIS3Js/62EvIQMsNyXFr2jXziBT2X6Vf8+DPKAH
lZyQUWsIIbjojUHC/78w/oR05sGIuOaUUShVIwsou2uFOB4vALfvpIwbO91coJvT
sBRGWVFuQpGqoJQ75Cfi8NXh0iLSU9Ux8XC87xrUULYJWD+QKNBUIC189K64bHxv
E4tB996ESdu825EajG8xdzyzJdxDy4/vFlXh2AkyDM7ThAqTPU3Xx4ZZBp/c7kpA
aJkhahlzPo5bK6RYFQtkaPflZXOzIXiaN1YR0R0Yha2en3Od9O3JWIVbGFYb/el2
gCDZVRu+f1MtrVYBaDkRfNPoRIdY1buLDC8wrTw7/a14kmGGYjq3rFMRsD7QxOrQ
zTGbD53NIzzum3WDCs/0b7wkWR4WYJvi8f/6ZB0C6JUfc69pr1o9IAfaInPVJZGI
Q4LuYY30dJSN5Yyuk/J9pdNgWrL+u+plTtYqvEt9ugA1Qlk4rIT79lLXEzDJ1R8E
YwpM9DevB0c08opcmB3FrG4mz1b7yfJ9n9KJTD9pDEWPZISWHNIaqkAI62CxFrsy
F7+2gooXXaCfpsEuoiILfXAQAvuUvdHCsyntXHjOLCOOQSW2SXPJlcUJQrN4ClnJ
/x1WnmuHug9dIKYW0sxAYeRDOnz1c8bXeGUhmmY/2SZ/QHWqZWkDqnCOvuYzt6sm
6dpc29mwURTYF7zjwmRTVrSoP3LsPFGJE+5ijDastpVLPNJ1dFZ7vAX1Z4w6bXeB
DOJonybjUYVE8G0P+MtNIIdzHbHe3Dojlu3klv+NfSxuBDaFiyclHoErVxG/nO39
yqfVAQ2dUOcnZYyUfS2a43yos2FGh4+t3G+riJegyW52Zy2rrptBgPjguyE7tQK6
R+07ZhrtLwKFpFanoTKAwggQVK0GNeoaaPCS11KIkH9/r+Ynvlg4R01DnElh0hIT
kOa9USdFAZd+N6TrPQcTdZx2+P2bxpMMd9nKZbMVWv3Qi7yA041TdXCm5HBAYf4v
uTLmS4nb4HwHwxRAA1c0q8EQLMqGGYLALn67vA5xY13kg98YXNYSNHYNS3A33Vue
BPW/I0sWEt/C8gTJpZqPpHp88iyoIwEGoLOyY9QC816DwPQcoqsEDFaaU7W6d+qb
fgcNaWOEQQqOrX+m9ufTN2KpdXY42dVK0G6NkRUkpXciclCTciLVimeOEK26kEgh
x6wUGgJgp1n6tz2HAIrrNe7tfv2/DDohTujJjyjn3dlhntmiwDygDRsvN4jVXuDH
+akmYn/T8+Zphs3LEDyHPqM+ccDsWgFqUaRCz9Gd6E/Gr94JldTE1RxjMi93vjUf
6P1+g1zR01EtBrTLQfZ0eUbPiJUhnwZ2sDpI2E5WCDz41zO0IklqNCkGudqH1ZqH
rnUKPYJHRfhIaIwHYgs02wBNVs7zUVvOfnIZ2ZbDIGU23/jbeKKvaswp9nvkv44L
y0SVcIgV/EmEiEOOOUIOMl8ayGVkJ9h2gZMWtGZ6y14Rb/xkAsn5dp+8Y2keW3ir
qbJ6k1lfYfdVlMLzluwgrk/ou6owEFzz5ZN5++Rt+yJyh0AbfREanmxZ/g+lJXr3
tsTFhAZBtRhTRusQfMfCOmBx04FTjEbInv+odgxlKykP+/XjmaGsigx9e3wsoS3F
rY173VkRVWu9mkQeBjovDpda+AmuI9U3mYxRKq9aI05Aq5i5gphczzhatJU2CuM5
u0rvN8B0AjZ2u+djocCcaSgb16fWy6m0XKzoje/EFG1Nk/GdyhhYHyEK1xa7wamu
8YZLRePk4BSWafJFXOasyQDyXDoXr4wyYq/IDjxPGMFtBb2q1hJMHrCZYYQ9sUxR
og4qV+66LOn66lRpacgO5R0Pj7zx9HNPVwg4DkaN0FiJvQ83Hd8ArKewkmwlg4wa
RUCe7M5fYvAEGEfQC9erIhofhPzfuFOQFFdNKEXIK4fU/I2EkcqZdPl9wzKDfB4a
o1q3a7hk0dR2Td0kSb9Dp6F7VVqQG+kr4MZxkc4TCjGrx7e9D6Nw30fIVOF95xQk
995uXcjSDf29Ae2U8vNnYEYgZ/IyPTP75sdseGDaChJF9SL1axpDj7j/1WFnBnVA
mrJdhgV4GvNlZEBQ5s2SaG7J61eM4OfaytPMA6Worp0zM/S0v/wkrTQflsRLxgmQ
gXTesKTAsbZ7hwQ1gBXqZv3hs22op18ccHDwstABNVjN6Q6EOob3qd7KZhKWP0mr
CrH+2n/aLrawSGG9qXykzNlYBrzT+pjuZS/8dh5lE06yylDI8X9i2MMt9vzyfdcE
Eld67GRJc+tZ0W/ZtiAzAB8yfCsVVXzbTi09Ati9MrbraaBdWl1DTGoQ4nlJzeh0
lyC9OGhFcpxx561+ctXH2092nEZ5E0QLuVvhn9GnY/PULOrYcbIxjyE6OXSD+Zod
YerZDFce3y6Ss3ZGJ4q4t3vMDUENVrFQNsKw9gneQ67U5A4La563Uwu9hICWtsJJ
BF3tZK7PEA25kLZCiwEB2jhNQR4jsHSOypKbyEtw+VmyL0MzshicpdjwuuWLXLwZ
NW6XajfIiijUuu2iRxUQi18ndkVVZPq3CzCGBJW3VeN3aRDBBP+bQXkpKjSqurPX
Vz0v3TLBkG+8VpTM00+4qcYu1OV2C/E723fepRiMyfeZ9BC9lPnrFsBH2eF+FpVK
8ngE6g1qf3wV4VypF0NRIt8DD889egfxg/l7FP8aPk86LNJLWLed+6QpY00LCbcv
IUUNbOtdWSM+ZVdr9t/6tdw1BM4eP+C4AewYiF42sb6e+cy52/rdux6kVtbV7I3u
QrY7poTQ28uInfaJu/IXNBzqusfg5Q1142ctVO+Jl0aPzC60iWS7qqhFD2N+098Y
NMMeJ3skzbRfJnW9/bdZwYR38kuUS99kEA41nZr1/basTiAnE5S2Q7XIGK1B6Kb8
FVpTvKSEmg2ZrF4Mf9m0uaRRzr+fA6G3GoylWgACIuxt5/Kxq3ZagSQeDynGWrfW
JXitpzMxT+RKlHTVsD6jqWDM7OAGehKrdt6FfnR6/DJwngB3E7xNWhsdXltaX0dt
T4mTJew0IOojlG8GQv4RX9MO9Iu3lkbffsSnK4Up/Tj1xnkFLWJFErkR0TUbMQL9
1goG27USRTaRkPl6xLvIUHv6FAiKCS/7RWft/0n5MupL3ro+cVflnzYgQSk8StHw
NNsgoujuRjTk9jpz3Hgzq/h09KlkEdxK/R6e3LywHWP4YNg9BaMjwoo0V5IVcEUg
dQGBwfkgaxygEin8qqeLL2lM/gvsrTftlCzjho0c/y8=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:26 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bzRLfcbeWYkMQmhVwD7Iz+bwFYwDjq7q7GKyLL1X57qBk83Tag4xXFtJO0P9MMOp
/QRrAhNmvy/LqwjutZviKq9PzV/OpGAzxTtpKpMxlVIn/WKETZnAcFktSVpi4/C9
qZwH7Z9nhj/cF4vS7MNbsfj4O0VrgkwtyOzAR1fkB44=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18512)
n4y9+1D/SaVRaGUReWLg8vjOil+dEqXp1iKCxCJLubgbA8v+p7G5dGh56qhyHpdI
tVgMVheoyv9zM50jFnveVbulNeaP1/UvoOsmeMMwruTAmkE9GZ0G9GK7nP6UJ9II
EwLDH5Cleg+NVeL9DZiInQKFUmUJUUEutxWF9Ep1yGr2eFbJfnpCYraY92KhFc/f
ODvCFIVyvbOKxq/+15NOK86X0l6j0NmFIJjjLS3W3Qo3KsXjqSubaEKXEzP4xnWW
WZbLszNxl52P1Dyb31viynnWsWHmZkMCXcwuxYk2rNJsN/72zwhxJe7diuieeo1t
Qk9PrArfmQWtWZmw3ui78fb24ak1S/d0vbkk7Tt5eeuuxgLdVJELs+riJl4Tu4xY
8O8bwQnBx1AshvdS+FWWr5zCNx6QlU41ZSgZ0wzyuFQG3XF7XHLmjSfKLmxNmynx
d1ACZdQdfHBE5et4jpnmjA+kkZdB+2I55t1NvsfhGPEx/kjSGQyZhqwYrZzqp2+K
oUL1JBqcpBgt4YRYISD/0r1BFSvbmE8eGoozplfumRZusGrx75CZ7SQUsgcm9pK0
bN3L5hEqDuK41JUx1jhJanKvexKnkERjvajwnESQ7SYm3I5RXWyR78D6XfE1ugRj
lIT61opi/V3EkSQQymYc3XONRSbRtFZ2dm0Au4bQb3igIvK6yWJJTImbjc5zcRbL
T17eWqMTHc1BjROC7rHADiwkywi6ACXVlR9qIyAJxKwXVtcG4/j/5KNOYBEGYpVN
7Ec3mtABAEVUflLp4m5aCXhk12nVSs4wTufPRyFn0Noy/EqVer4GYBORhM25N9tN
N+9dI/3uu57CW7LsXHtvAXqDsBBQPNJjCnsLUueYCOJVSgIeS+G+xiIlWoMsZ0FG
BlySCqEKGz+QLgR1Gx1icf4aovHv0ujePu1uhhMXW/RpQowAW4AH7XVn20uHwpz6
tZmzK+DvZb6Jpja0kyoaBNcqdGRktkHAhKVwUMSA4nZFg7s5goSbLtqR/F6tmlfh
jKX64LCxo0VFMBjTOBbTe+eKDJdqUR55f0FZck2DTlc/4UJbZ8ZinTwd66wsQe/o
dtiUTR05L11FrUGPsxSosSd7WGwpG4wLE4kf9KBb7DLYYu+euk5jhUUjYThEgMXp
2I5Z9tgheWx6pC8KZ/oamjHUMvujNrHBU3l3gYXw+CZeqaX/dsFtmaLBzYk+PA/H
8/MVaZaCbEQyKYYBhRglpNzqrW57LjJhVa/sYcLCyKYkR1YUFDQyK0pqoA3UImHk
4y2geLoXnd+UKZzhtjueGCflomKg+uNckUlBP7uv3RzDTY63n2y68JGka7o1ag8e
PyfnJE7FtiKDwwku+daeGj4G3IWR+eIv4Q2CXDlhuw+XsZtQJnfwQyugSdz5f+6u
WebZbKc1akAVlNdMGV04j4jYJO5FxdQ+W0pnlClFrM0lalXPx/5/Niqf6POAGw/t
UfTwj5vw1p95rsFKgltQsXKiieQ7Fl4yY7D9zRogIbXPXWv5i0YGsn2iKZhGlVpc
L8GiLxKS1rtmRDj9aYsY7az/aLEoHTqSu83RfixPI8TLgrWcKMvsl/iyAmfuoA47
uBfev09kYMuTCC9U/NqaHmIinme2zKC1W2CGT2Kru1Y4eyWiSLsNMgmJE19ERRn+
QP4QQdLPn7DNvz13ZIwEj3jTJ8Zi9rbhqfj7OfM1+r497v9saIJZ4X669hlM0LGL
fmytz4C0Ame63CtggquQcZrga8QIfAwzyJUIXVBVenrmAvSFcJk8AT7V7iLTvnUF
JFWpcijo8gPQj3kl66f7CMcf/5HSH6YQHy5rQZ/0knqj+i0JClNjQdpjTk1FxjLv
Z43X4G680CGbVNH7BU9JzeiWz3VXPQ3Eovdv+8vnz6AUF1Sb5lHV3daDN51TPrvx
B/p4Nz9S8l1RMMMFBW/GX8gYGe4CewqC5YtTN/yCgqOTMKTDbqzG5EEeRmwG6gqH
eIIhqEkUzun2WaYsJDL1MvP9PrXVHyVGY+C3ythn21uvRkiZFnqvadzP177RLN0W
trN6P5UzRJfKObCS0V83tgpZpO15b943oO1SZ2ZgQXD2Gscx4uebO+G5+JYH1FmM
ZxfEGCFnglKL7B2jJWmWdOif+a96i0C+tHwIPUJMogz7tpe/UUfgx997W75XHYM9
RjUtC3FFxFILELfSXtgYnoyrRCiXcM8e8L7hJt2a8+jxyovRURpbFzL4vzPinM4q
gASIBHEkagDPRd5wMLaWU5upEH2eSV5Qb/egKHGUs9Vu97kObWeFLQL5YWbkvIvn
kopfRyra4taC8rJ2eTWyxCM0rXU1SdAl6lhqUSt1EQGfGcIG5UfZYuecb+Qi1yPp
qb7C+sd7CGrbAU33n5g+Yf5Y2xXLal4OPyXmfSo5rVPdxe2mwIlOdwptsbAp6wAT
76krnM6Rcew22dF0fp+RJjLYggJHzqkciC4Z7dtbdWpYkyuO2zD8EPP5DArWNQXq
+4V/nqnIj+qdB8zYc6G94zqJ1UFKPsVBD8ZO85NCFEDZ89D32AkJerID54gACUpV
5kIqwuGtd9Xuyge7kHPX3DLoPLdP/sRNFUVSG6PPHB7CEdDYeNesciOwgY9o/ovr
zcNk0k8UUfadPU1DEitvpPfrXcNNJZ7He9EaZzIzSw9kUlSp3zkc4wYs4sfoK2he
vzQrsFDffJksTdzzCgxiuO9oQBiMZYfu9NQ55yBIFe/Xo+CS2J+WixBMnP7elJoA
WouW7gKV6QTNBJeb4vhNdD99kCMse8e8xLkYMDU5gOf1YFbhw3emyAsI73l577Y8
bhZEjkFPWnzH/YPs2d4CHmKWLE2zEP0Z4XsAAVU4oWdzrhszH9xHomWll/tsYLya
crxkJDo0eoRakc7ix6tRFdXJrzppTy18+5qepI800LenfrdjdljXWNyRqBovGYtF
6MMeEM58SKQvy4sbqWiy8G/rcOdjy7Vtc1UksQcvS0/ZzafR1a3V6WZtDWtUTpPw
Oh+XZgMMT3hcU7ODFB8cb4loRqqB47t37pqTI7tPSqaaukzNwnP22NZBoDXN9GOC
Vupmw6h1Rl6IUDcjmxmyXn8yTbG2fWrMQG6u+DKWvz1gBMJpkam+EK5W0UlQotzd
fhzDpE8gHTCySKJx/1uIlRTyy3S6NRamRSPvASNUNw5HGkxcJ+cF5aCqsqyJ8IjH
ULq0Lg6cS6iZk3kYD1fJ8NfdswLUKLuMXCVv+jhWgLawNbKHmGGoOzNBypKvkuOD
AOMJWojd+rpD9TAvisvPzEPZHYsTlxSRbwgiDwOieTPsP18SdQuv7T0ozC8yhmt3
F+MfmQgSEkHXfahH8n1PohUzq9gAs9euCVJbkVaqTBrdmwjDsqatfXUFK36w2RvG
PPA/mjbCcuS4G0666h7WuAShdANzUKLh3FZP/0qQhgvS4fckY4jibKGDTTs0htAR
/yHvQf/NACyz8P84qXR7Z7UcpPXBKQ36oGvAYMzFnPquZ0H5oL+7QMIxD4l+60Lr
Hn/1MskMmq0NnGqB16fVr/XPB9n0kEcf2+m/MR8Zi9TkvQ5c62Lc+QdQoPLKU4YV
EPNIX7a/rFRRRRklCGGoSKIcsw/JgSOyu2TiupxDVM91pyYSqhycM0dZo9BrRV4G
RpzyeIs6tkn0+Ipi1qimG2atkm679nrdYVt5Sa1+glqG7byyH3nt3yK04l6pOSTu
92NyxuzaS2xxaGR7Sj20NUuE9IN9qW+OzSZGCQbC3w2iRD8I4Zt/EWKOCvc8F0WX
mgCN5ci2yYolMh7Um+hzzM1ykBhwWkaHLlViwYNexlE9h8mV2OWOwJX19gM5An20
i7EdY1Chyepkxo+bBa1xdrcb+1bIRqZyBdKWs2Zk4kH2MgXZJad2OhOV1zk1XR84
kkWbyXy9hrQIXRCFMUrfwXvj4lGk8+JW+4clLTTQtYgOjodNkLTafo92oeG19khv
12Cmjz+dnMq1QXmhYD8i/C5c9UQ17K0CeY3au1lscrK9HYAIP4giJs+RdXYjohYo
e/+4De6v/OK2NQHBHEtV3YzyGjRvb008rvJYQVTl5krUBEJQRMb2D9XOJAwbDSh0
80DhSGBbSu6g6ZSo9nTsURGOnD9jRvZK7au7Y0XidcEGaLPixzXoP1v1ITnvblvi
u3dSY659kRaOJSsxlMNkUIOhpjI2rcyzoG0RV2eYV27pSBqXnA5iT4UY4bdj6IRt
DWCjjbjWNDHmiZht18kw77IRQY0nmtZGh7cMLm6Uwe2yG1v1tYxE41mH9hxshJr0
gyepKJfMxV7ONIwLMhrlZQY+ufBcazsCdgy0SHZ8k2RF2iM0dcguE2tryYQauX0F
1YveDHqHy7U3kGWc/s4+Rf+W8fwGKoUWRutnFA0l7ELQ6MfwxuDZiB/zt+M7AY6c
sVuZhdyUn2fBWO/Aso/05w4Ww0MxXGQazuv7DuoU35zhumrWU3Ks5mr5BGJrSB1A
D2yWCa6U1USL/ifJJ7n8MIClsYVM02QVI/I/J6fOUDxeq5U+sHmwT5zOvmTV/qAF
ftkoiyHoAUcoQM/1aNmRnloFr8Dt+Zl3DjMwmIBZrlN6UFVwkdepO4vTj4n+4ZPu
z//5MN/qiPFgF5A2zvwqsvQRVFwhcYF5fPEn1OEpAlKPZWh7n2zIeKZHeEdS083H
J5m0TsvPR1CaZeVwJvrv2G8XXgf7MhN1b9ZXF1KFUv7MqWTFXTYGmHSXKsM6zt2i
sQLkq8OsH+cr1U3Oyxq2ZKsFiCFEbEDPblBCaqVec0BbzfS/LBHUY4PmAooGDilJ
FZOxqbgfjHbycE5JsKsisxlbh2/rPgJVeegYI7sPKOzohjCwW5/Uq/0Y5YNK288i
r1iG3tRk0ONwS7kg6XJR+G7h03ElgVCJ+W8PtZw/CMWDAZl9051QKCKBtaYIuIBL
qQNf/JMC6ghLd4OCqYmZj7RZ5wzKB5KcQ7qmt28tlgF1CunobrdVz2WN8XWztlMo
IDl18VbnafONbGFYlHJzPG3i2IQOf/GkStmqPMDvvPjLp2RjYxHOvzF0aKcX6diD
qqafQgPCeeeAoo5lyzCCYy2V90eTIO3aaZw5NG3m7lTYuU0D2IDF5EXSF7gzOqDx
JxvhnR2DVAmKXXoz0gXSeykDnQUJLsZGTEQPMJq7Zj6SohQb7IbCRQ+20cqZp45E
y9SjOCNXrjhew/OAbnmkfspUHOdgvb8wTxuNLt+PICM2Z3lZO5LkEvIiik2KuTQ5
S7eRuhyXJOd/jAvu3PRZTQ1zSScb6nvuNSBDK8MT2FTBxnS0f3Fddvv94DoJM2nw
Eat+3T4AeYOm0o5VNquoiQVdPoyRevA7D5WbcCoOJDIq3FtRlBjQDydz7Vf6q4Uf
GLiO0poUglvVvvcUzD6aDavirdJulVGy0xGi5//HuXDi1iNLTyY5+GUKZwi8zhn1
nZeQkHlNcEcT0zj186uUM4G7sU2/MgSFJsAGIhiJ2f1T5SOFlfHTiju1Hr5X3scA
TjBiCSuXrWMOAj/QeALMFwikcSiiyx8EjO/suG74JeK8j0phajZxA0ZDQ4PWHYwl
hV3OR8GpxGp1qrwCe5dVkhQtHzr6jIz7OzscDoO3CyXe5Dz22G/soIYhlezTvYj+
wp/XC2vL89PbN483zkSeYKJuATATSi9yEh4AuGogr3g1b4ErQyHl4mWrCvnSHlFl
A1ZwEg+zlY5NMvBLr9OLcsuBEziyAlpjOJuSHWYBIU6YQpofB0NehkGG1kgOZDh/
lNU0NiK8mkVbqK9LNsJZSQFGOOq1XJ9fVY87VoA6ViwSN+7GLHc6grjB/36nRJpd
VD8+yLREzpUUKL8AM3TAm+bSGdKTmkXxZDWBs1aEv4Z7QHkM9vI8+B8rjqy1mOjG
pVBSgrqy4FXuTPnc7N5LQRpaUI4ms16VN/cebmKvJZdWjqX6EMAeRsVob/d3B1pg
XzYVBQqPGIucHYN5yNYMT6wAL5NT/kAysebidJ3M4zmiTixpxx/g7UiDcFicNY8u
5CmV182BnkxgFqUpEoSVnwwEW4J6246iCae2LqtsFTiaGItuhHD/t9IQw6zLxCaj
myFPVrjlaXoSaSo5JpQ2m3DzO3RG3WkT1q7L6ciNJZClKZOblZ7sOoCs+kjKx0On
CrEfwygUfE5nxCz8jS4/ruKb/ouE6RXO8yQpGdbK0lAjl8eHQRTqI8t1WI9FGDNE
OwF5xtWVI0xEW+rkGnAiLc5kEE2MXGYVyRbUipJ2OfimPKb9X7909KKj3ZqpVOSm
I0xX5HAHw/8+DiLBtY0NqBD2e6UwvxV0p0Ujj64XLnRlj72qOPC+YSBiwKm2Wzu4
F2UMLyNiicZU2Lf07gOBWlifelDwNNOvA0y2w04CrEVwXoufv9HMw/bIXAlGSKfH
FjMgz1vvLNWoUj3ZC30XTm5il9PiSS/MbjxldzxHtCBtt37kEV8q00ozV8/U07f5
t45isD1OdSzkaS9pH6XdMUNIvG81WtckV7GK2hW9iZgPSqYPO3wKXj7tnmSAoo6+
SsSmyDOnr+Z/aVpeu0gBcGD0tdcYrAlrWb8EQI67eAfueGTJeMDNCdWJGJUkiHx+
xfMZHvcuM6i8n92VyNPMaUmGedq5BBpS43pXXxZqnHFO5fm3otz5bo/1Cdi24AIy
hJoNyUaaL0pfg/jKW6PbmtR0sgYD4fntu2O0pR5za3D2rQLDUwn9uSCCG9BDvsDe
nMG4Do9NshoBPXc98XleuctbBrWx8NIbzr9zUZU5epirzSd6DOpBNIfrkjP7djIB
jRcZRcz/BTuEcGGaz/+iQzBz9bhYsbJoqAHQl+7tq4okiwU4TeES07zOPxXBpBSV
8FUtXl3SxMDFpZh3QjRj6yB2x46tBZS3oUYPaTVN814E8a1bntMxa456n49Pn7G3
CU7Vv3ppVKCUOXXU57j3Rxg4kkLp2FdpVeRnz79gWdLF+QZ3jnjBlSR8bX7YrImN
NfgHQPjK9P8s7dbFzl/XhMRiOCBUuaRWlGP8qXa8XrJ1uT9DrqUcS0ttXcwwujqb
8pmduxmfm4epy4uThBTh8+UsAyKK/Fv2eiy/VefJQgcMh44C73Dwwpy5DhF9eEFq
9/Q0p05U1nULReh1g7g2s2umhHljrAeHIzdC/fCGMiwpal95kGMKB/27DyWhukDu
TAA+XBSvC+GNZshgQQccNaJetX2mPs74yq4MxOaSmU3fu8vkBM2fhRBC22VAB9P0
KbDrw4VsvBwKJFf6/eMIeYB9EDoZJ2p7wJtBsz0L0wqxXHbQ6SLdgLyQW5tC+B4i
lp2CkJoVxD8X5KAalfKEcmf8E8uBThFZBumF821VO3h39zvFcho+fEBKcCmyAR/L
1MZe1THKHwxoczZSNffCAldKccDMClDuUHRqB2j83HngBsbprofpToGaony5EPQp
1cnggx7PTwzJ9Qg8j60JsXtJil2T+9tltKsU/f5wnEYTdZTBigWEeXx1bpAfBMaW
l0blCryVpNyGot0X+70VW2tYxhoIJ7q4TJSudUHIiIG67j3O3WELbQ4Hi4qtvcWK
1MQ4v8/tozmTiaABT+adQcuc+ohRFZqvH1XPmolh8E1Y/7aAPHyr6GqX9Z2TDYlf
zBRAoLbaGUO6SFWgY9JNSNs6kxZD/rmhiYz0rfU+kvlZVi0wuWH/g8Ru0U8FSpjE
A30lEGZtNT9LTkFgvj81DdqBjFxAzXw58FZZ/3F2fbkEGrCkfn4TyjYrG75nhxNL
STQ2CZDL7EPk0BOGyQMcCd8+2DYzNbHWcN5XVEhpc4tKFsRh66b3UTaeGpI7UFf0
vWy+DB7+w8mD3Jz5mcI71PF4YhgSuDAFsn6UeHx/IZ4XEr4r+48W7KKuIUvtLZfg
o7kWomwFQXEsoGOIpXUvyhNVhqPuNnHl5SauKmDDo9/dG63Ia4xnxBsSH9XFEPwP
Gd8M9mIMyYOHfVgo0DBq4Jyq6ru8TRAE0ff2fLp2biZFg5yJbJvIPMzc5dN7DAzh
mdVSGAaqBL1PHFKJq4Ne3J8R5oMUGG/4cN1AXDdgOKIeVoKp9BwsQLKPE872n5P1
Rh5SMM7cv+QEjna87RZovtf6qTo40x5vilvSAipCY7Yq5vo9l1yJml9/ZvTer8x9
l7KIZEPRGLtT9lgHuducQEEsVoKXaKjIPPQTGLSeS50IQ1CThTiQS5bjobaaZvz5
SF5YESSl6rAdu9H927Ihu6+8L1dYI0Np/E241cGV31TlSfGcuC/WhzsIVVs5e/CX
6uXFRccEsvFOzN5UMnjrRfWyhs+noYFCrDTgz9aSRjB+3dxTAuHcZ577WIlSZ5KG
T0bL8E+7W9AwH1vC8JdzzasJga3MXyzuxeLJzl+f+H5pRCr9HfqzZmOs+nvgrSVc
jue/0a0I8TpzOe7Pa0AkcY9/VS3WKGusRO4DRMt/x/oetPzllBERezbrHeNr1iT6
2CwzYwf/xwS/5Sz13ikWopAR8mEF6dMwJQvSaEDauI5zRuwr6S4GWr+MFhFEpTy/
2+Qj75d2AQNPqn4oPko3yd66EX6owUr25n2jUi/HPQKxoN8ZFaB81al/8gIpN7hE
ffIz3A+2cbKE2CLU/XzOHjc1+XWBOD2xgJDvyR8xxBXNg6aIRIfp+U7o49zTvSjL
bC3DXU5WN7BYg3u5GZJ9FOr6C3e7/yYCWV7J/IKfjxeiHnyxZ8v25UQLivpGsqhm
IDDuXCrH1wKIIWCXj5h6IrKHc2tfxB0e4sjfkueX5TLqVgErKoDyzRp39i1DtKyQ
zHHsp2vDCChff/xWgSaJOVsPNSw8VAeWtj+ww6O42xe8GRrtWatq++D35yW6zTmE
NIXXv9/PQ7Il7ayCnU5NFpJKuZp4LtRDz9kZA8I/sNXvADa0UQ44PcY0bPo27ehy
qmkhwD030AteYGB4X3Qa5tzvgheYFwFHA2WAmHqnD0hnANMrD1gEM66hnK9p+gCT
MpDFYVy9/Zd2gaUdtcfAagaSLrk7/GYKAH1Mkk7OL9VFCfgLX8S5mupwbaUQSOmC
Zq8BJnb29wEPEznNAadoZp1juwcj+9n7TnWRLgZ3CQELG6dLYEGTVYR1/cuMO/jD
5jZGh2sNftWHJDnXiUSEjAduMMRwlNATRIDAx1nlxeJmuqf0i6apeBjWRDEfK04M
fbvNYJHpN+s+4Tp4OfqFniqqv2Wt8v2VJygT6QmcEwFWJ0QOvp87MHYjtehILnhX
4U7t5hdWdajQBaFcdlaLKI67NmPQgaVnOUQke6dc7x+sSVeFOnTmGX4sCHqbVqbj
4vEHP/agYhWyi7jktyWtfRCzVZ9mpkM77VBrTDeM2CrvBjhh8692DYTD65qvwhBL
HOMFXTf8J/8otygkdah2BdYEVITjWp41XybKA+/qrJwZOSgsLkGy0mN4ZWO+cLMB
HDjBd0+OH+idR0AN9szDTvQjgGFklhM9fa40sJ9aN+pfTqytd7gpuWo7C3ypBGyw
wpvGwKHXvI5dty9rDJZUiW76pNbEJ9CFoYIdFr19wCjDuzqw19dCHEx7Dc/f7PLL
d1TP9Q6HzOSO34brhkYr8scQhIHfuWdARDGyuTNVnibOmvAhr8O1drHk2AGCRvhY
kt7Gi+4oZA0Hyr4KZ4U9YIrDyOimFmzgnkYQtMSYXslE88ciTMjbRla/xe/Eu7cr
zRewVvm6OvGJMkYjIN8oEJwcJ4LEhRLcKe8hQ518m1VG+QZHh7USnAYaJ0g0k8tR
B1ZIPrQHUsQ2COkOb5gEkLREnzdogsrgZI22t5k89Gp7gJIu8W2TcD1xB7iVX6Mu
RU6x21GKpn7t01gs8RL/llZq58abapipejSEoeg3UXVzv5wRGQz26tFlMElgo5N9
iUX2q2x3r/sKl53/Ec6mH2hNMOUkdWHrcoYDWcNTzyGgcI3v9aL8ws3QoxGtWxHj
V+jsKQtO1B9TW0jyICYw+cpYoOZDHxX/i0whv0i6ve8/Paw7eS0YZ4iLyr/vA/lz
g6OZe8uOOupoDxYNOyS2dbEOzVJmI01u+yO57itobXbhWkVKUVSIs6yxN0VC6IGR
Lvq9jVXMXqbawwc+0lNMsgYYh0gi8rZ3yZQqjv0dwg8+6HzezLinpa20jAZCBwM2
GbsL26CEG0ajOyylZyAlq2YIlP2JgDKKLlH52XfZs8STAWASgE/TsW//OnUCm+V8
MbRuE/6VJ+V5PzyeOh81Qz3ZQpnJ1Z+XK2Va4gYEQacBpL8PWQ1GDpF28cC+rPxH
V0ovx44heysVCzZVyXTVHDIDa84GdpffDTO0Wec8gIVS0X+2qY/L24s8XeyjGDid
KyHNsqqC3zT4Z8haEmwZ6ZVvpVkL8BKd+l+DTsy0l/GCEmS8gGE9Q3MlIvUZWeT/
9DrIlorQ4iBAGiuGzqwixsH3MWwyPJS3vNETwetN5yashh1C/P5QE1ubwHIeFN7W
0v7AsooauxM96UmMyx1dAXmh+SYp7PMTMQPS2sv13Mkb+It7hhMA3qI6XYf34eF1
OnFkNmcmdFM/ojBLItjbNPlQlpoROarxZGSjuY0DrjrMiXEkIuIAK3b97OYA8CE2
6ZD4qftmwavEvklCaSTT8EXzijl9FrR4A4kVa2sumtzfduNhz+kj7D1EYxOxgaCx
DNHrYc8fCX1fR7l3N2PZEhLIwP4Yrk3COTH4OJRC1wuPH4eLjWV3Kn0gd31Etvf8
45+dzUv5utJ2P67u3DIqe1396UtgesI3rdR61OT0ZQKSvcGhfYOjv0G52oFw5w2K
BP5DmwG61MRHTnwPS3ExHhU4QENJm7AbDSJhw0CQHTFecmlWOZZm+51M0Hu0J99K
kaipzgMbD+am6e7lwb/oZ7BMv1mzJ/QGcvVJgCwGUlJL2EJGRIw3thEUlzb6mX3G
v0cClaVV7VuLVPgCdvETX6PEolCzHlAT5YlUmBTiKK5EJcCFsJITobo0v7lPIRlL
0hvm4o0ohhbgnHlxzapDhOK6rTgzwFfv96K1A9TSIcyvBA6t69mV6qx2v3nKIok5
MHAjjhwoHOfMJ0mlxEyo78H7xd13LNoVUfszH0B6o3goz/0MXoeB181lmi8VYLsA
jgU/DVJcwNMTjH+GHyKZLCrqd2yiLbKI4yN8s9lIHGxv75HBgAOJzFZgH0lVVo58
S7amHSqYc/sh5NpWui346FM55BirG9dlndjAvauzwIQSHvhkYfn2gWFh2xpc5IFk
++qvHcszHYitC55dL51lGTG8g/iXbVxJ+QEQlEglSWXC+e7LXfLWGih4e8SFa4Mt
oecR84pzTj6iTyhuHVsudIYmSvRAElMXFTHxSTrGc8EzXiaYjbG9SxSCI7fukXeI
oLnG/sA5MVKIMjsms19pd7zHkS1del9DCW2hVQfUAggSAlH/AC8ljQsjoLTRQNRt
FN5paS9rCGF0vKFpPSYBZ55qLQhLfI6TK3VqI3f6W3Zn2y+WRhSyhZYk2+Jm8VsB
Ca0qdf2fpjAPKmErPQ4vm4jydO0sviskAytLRtZRXo8/Xd34wvaJwcpWdszinBzG
6t5rrOkCiZns/sQEc9LJWblA15qtpD4UTtp3PB0q3lZqTObAuBzCJOLRyiOFbZBC
wPolcij82gGyUNcsPPQJ+b8IaK6q1VBC9Y7Km/oxdrjCrW5EawdgCXbtUBbpuYQk
1sUpbDm7t5jjGKdZTx/T0J1GWPvEdeMviahDiFm+GBFIGSZWctJ8ZpDtC6RPAdYE
c6ao44nxAxDyeFavY6LWhLKQvlU8ElRoeqIOGOQPNwUbUS/0hxc5qSeC3Fd1uYkI
O0kvajXKshVrhLE6BUfweb0liBRZUlAKCRVfTWXCSt0uxiM872qvMMeCfNIyhfea
AQl6ksDJfR9tcOFS0c/cTFNkzFTAniut2SHdC/KKz3bgJIaXhYfupMO36Ic03F60
eWcVIJnh0sAOlWk7qosqcwZ1X5Go2f6VEHdihpZPuglULjv9uip2aA3+KU0V5rNQ
VVlJyFlSbzg3nBGzBkLdkahY9CSZQaHFcVfqULBesMyc4nvsSnAJUBTKICF+uMUG
2OPTBI3qZnWG/A7+g74N80aKB9Qa5zw/ZBSToePd4j4V0o0ezcAtfh7FpIrs9REP
ShbldQJHxYjfjH6Kj+ZmJVBcy0BC5AlxVwFSl7dU90srL09HpilbWk64sUg5adza
6xTJruz87fp3IRPg3bMAXvdGu5FwOuIQIWOAV0jzOlJ/10P/KbaP7FI6A06jaSWp
tQFzPvyMohPb727Sjzt9H4/ksk9u4sLXlGfGYVPsltnUtlkM1zfFbUdvlR8fKwwA
OKvvsyo3zMiN7YBMqjoEAI1RARxzid/726gFkp564X/efECRXqlXxaCQLZjt0zSS
PnvG33diKkh03niO1Xsiu8cwCYTT7/G9lEkOXXwlk+phfizY/joMiPYnggS+W87Z
nW8llekO8su2YILpYF8FmUTJU4hwjiIQm7OYHf0Mq/LSqpPde1po97Bp29bNFyCd
cArq6vsvH7sXYcPxghbrWfIgkjkupm8WZanJ9tKP3dP8zqXohbpejsmteWnpZPN/
EkTBbwPkzeZLUknQqTp4FP17q+sNG3CEQguIpX/9smJ2OMw4mpmF5mYeRAJ8RcJe
UFcN8RhEwvgWftwTyXoEGXp4X0gnuAMGCOqPc3eWFs1uIzEic5K+Lfjn12MAYr1V
uJLohA/tfyiOcUMYtivS3lf0PpiYmGAbkFTMq8jDCl1ElqxuYbH93C+KAG/YG+n3
vjNwfT71tDX2YWPgzZqxMkV1SSyfNhtaWvuvgsVwZN1tSTmet/QJMv6QZl0XFHJi
T98g3/8c9CU7W7N0KLJvudSquC6sDRB/JMxIDeOKkzX5uiWPhzMF2n+VGp6r34Xu
JVA1k4on66apg5IzmYkZ+H4wTzrCT1/MyjZDKK0S47H9u4Eh05ObcV3hSFq7kYsm
wFavwFVKvn61MLhR8yR7CY0ZfaUm4H90beIPvi+hUAvqrv8WIlwVJwAIIjJ2Xc2R
2xDtTPV0BnX7Q9Mv7FS32442uHR+v4kdGVjDuEcUh2KBwop96SGY9DBLaWsy6TZI
nTTEUzKmJ43CZzB217WYZtoYXin8HB2w2vL2XPekI0TRG/XIXNGCe8lmcIf6YzLr
hgFf5FX3Pt3ZIhgF4BTMkVHtYkuS/z/7SjdDmpt/ukNf7bnDFokPVAITqEbFpYHe
LFE3NazZvWdGq/bvSY1ynEdOVeJn7dGY4kagytXOCzeXQvD6Ut4l6X4i4gxABJfW
WMhoWjkKyscetlo04KctTp0rqqac+uXBmT2c59IA5Hq6ffOb5Y3kvlOA9qSyfLRx
HUT9CMTqS/G8+7+ZOm90hZRfKzRQFH/PAKOHEYMSEY5+Ekoe3Y21ljJBQYoGn9xJ
UjBpZszcMKwZkkIxGCgqqbEIl27u4rZAB5r6w+C/j3w8N66oN1TxF5w//1I+whOa
QFiceKZA5j+MKDrgKe9gDrjdRg8teHfgKtbRvHpUp5yOo2MwpYVX6x6F4G4mnyzS
Wzdy4Ziw///r7CUcC4FtVS/UPMT5lwMDwhefQu1Ca2Yx05E2F086wDWU68RiOqKJ
Z5McG+jNZcMO6p581P5RMWa2BX6ZwGgq3+1hDAB21LD7G62Fny73Bikldr1KLD5e
JHZHFKO4NP4HH8fJVtTv8xvJh6ehh2MUaoA23J+opB27IS9agG4YGkKHP14wHQvI
gDxgqwji0sCUKEyNWr2JWVi2YyjnNTrci9ZT3tG2oklBqfUsIIPYANjNt0fKvIb1
X1+Ma5S5e4j/xcaHPuJeWB76bPmtr+9C4eATJeqQlzllz5yeTKbYSUPEYRYXp2XR
Dwkpp+QHJJa1YbhoZf0QULn56IiaVHDqUCXeHj5C13jVDbZMuOJQzqJ4+4c7f2/W
pCCEXeEPQxkI/z+oBDssUA0hf1DBJqXGLnLxpx3ROZVGdz6YsKH9oAOgfsDsw0iN
LSxQJUYeesEtecVbroF4tX2cbVSGNiniAp1U2FZD32UDtjkR7gsYuphNZP0GSxoo
dIqcdyBX1CkMgO7Ea3riY9wIZCdmaMCNf4/2tJBplrFWXd/eEDmxekpyhKB0gvtl
0F8PyvqKzAK0r7kaCHtJUzATqxaULK0fgJWVlqJTDawPxU72HcMECNCuEIhpwH6C
HoEoBll6WRwp8Ou0VPXG69vjuqrM1lH9/4GjIMDXDyjLIJPWaqNKQrDbyf3zE6nc
qpR5I0WrRy7Wy40+K/9blgGYU6LEcpku1FdCZC7kRWv6bDlPnjgMGgRj7s0m8tLB
Mb6nUrVrjiP9dZiQuYWSbhZJ26tqLfJQOpUaP7lvTrN0mLLnvJwypKqokkgaXdSt
okQ6bx+KpYMjlVWkGGaUZ2q2bpDl1mSovkBYONlsZRbpAODCvnUYEtSJQZ0fnojx
yIqzy0FPJeUVMgfiPNpeTUJlshV1FNJszwvNhc6zcA8+Gyj2GhkM4ITL/aPblvnb
IFotvzzUQVm6rmnbshIC8z7YGt8m/86U/lReZTLcZMbzWnh0p9zPzNcldrofya/p
KZquz5tTkQMxhihWatb63nbgPtiryJRDTVernP4jDXtdmSOUWlntXT/kPfS4TGUB
gkc1eokNcuJOaHVZApes0VzhG5k1q6EnJPdz4pvehWnBvYoZ9HrfVCNH+EVuCcVV
Da7ube3TTeHZenE5O7OK5+/jM0DmxtKcdzk1B15WL6tOMIpY85WEKw9Fdxp9RNkg
/pTGnVY4y0kLrOXZZChuz1Q6fCnan6xJsTySwE3txQFMYIDGvYimK5dTG7KahIGK
3MBXm8xkypvaUih9N+x4c60sfhyLZrrn1MiDhshxZmo+iXbmSpuJQteSM2VuA1yo
2X73+1WcZ8R6EKGQ9w+zxgLOLpxN9GBC+eVS+2EbvHwANeWK85Bp6if6668OWH/n
MYg82PcT3Vv5KseqDs6jWguRKDPqBejQXKx42dqSvPQIdhQxuVhYFvtoL6xyHN/6
nqrnawpdqcZ5DXh/D+Dz0nudSnF1mT+g81h2QvoYw8gHdVy1bn/dXXK+e2j0MeE7
UBd5grMxhjZRNM+Fn3CNQA83qSnxZgjpgVESOJv9q8Lh8IFjKknx+ylfbiRJKbwx
P2fIx/sqftyzUj26uPlDfOu+973Zz+8+gnkKHxZfth/tmed3N0EGy/YsXAsZESvF
EuBjJdYsH49zCQw5HNATh/3N2n9Bqm8fXtHdoNKhvAKmKC2cD7uBKrHtUucz/xrd
CU2g3NykGTXpGAqSVfeZzfqa7nkVElUCoYJUV/1qnU6pFnhR5purOW/U1x2MzBtm
I7IVCkUgVvK8QLh3CrOtfjjY+pxTy1ckMSapQMcSZLEGojJ40G6Le7pG285zDriW
ZQNyYDdROTWk32LAJgMu1XIty7WWZAtpWmQ/oNH+eGo9xdpl53d92Mvq4Mcw5OY6
Fby2xENYBm+DkNPfW5eZ46Tiy6ws+h7tDJZqvc23EXe8YAm24rByqgD6E+UEzr3p
kLnQ98p7HHewrTtOMpm+7bX5jbqfbFZ6IKLv3+7EiDuROJvUDDkD1fSdNflv0cF2
KBC5/I7is9FiSwRM6q4TJtnuTaAzrE0irI/HYiXqNLgd6zu/w7bAgHFN8nY5Yn16
ENUXG7dGByai29ArZ8iN6WGagftFCNAacWOlN/VghmFmpaT7p+4FbWDoyyIi9GmK
pTua/nTehpn1G2TDEfA48nX4QjgVqr38oVpZFMRuYs4+a9WgIcrliG5cHl1nkT14
TebCA6OROuYzaKxP6yD3omvwf7/lBQNeb2vnIXjjUIRQIlVGbf+XaBBOX4UUar/y
yXL7qqKGuyEfZTpNSk+fhEcg15WuUO8ekH1eAkYytyj61usGi0JlHC0cE4THZAvY
pmeRv/Qh6/QPTHRNjGqWHxS18kxBvTSwiJMiPkCloUOrpwtcZASb/Jedw6bXxVZJ
LK8l+Y6u1UuescgdTN92jbjCLIH2NB5nowbLOix+Ef1hpXk2YyFX3h3VGjfBkFyx
513mK0mew3XQeCqHf+c3hRtQKqDHtSnx5tOJYpPPGuRW0X6n5tCiDor8/5k57lHB
f6Tb4aqsH+4CechYf9wCgDd4h3djLygjWSoBZtJiQoXLWCVLgv2Y2XW6qJXjfDaz
E3jxu0/+qbrKeqZjm1lLdiqrBY5vKiB+aHLCxOql6ofCCHKBI0je3cIB9BNKosw0
uPNwm34Qun71uyVVi3G5RsVNjOHvEWZUlgzdlooOFo4HDwG2OeXuKeeWKJklbrd4
R4azN3EoDoyS0qBrq4jbSyY6EPOvhvRBPDNgOff+aPcHxH7hLlLfcbHbDc8m1+Ra
IT56g2jUnZlu5FfPTY/r1V28HHSAl8OlQa0NuW6tyBu+94Hps/I+zdPgHtuzv10Q
63a3E9vnVJ2ukzjeAimIaTKePNWYJsiksBnEdeAfIjcmbxrPvcppxxG5VyiNdNGj
ubZXbW3kQq9XKCpFDDViFr3suH/VAjgtsnY324e8eTjje8JmoP5076DhUtDNl9Ig
mo7+bOicvv2IqLaYFX2dBbhyiv3PIB+6cVfIC0dMODCCuQ7mvco9i+CGqhvnMg5P
WchNGc9XRmPRAIiswYgw8Qku+B99eH/m6vdcAa9aQJ4ZC5SJShSlN6b98NFieT6O
c36A8vti0/kTn0Ad8WSo6yaPef4R7nyYFAH/ai7sI/6kxGfplr2lROhpeugFjxSK
f6lVE636y9Q2fGdeObE3TXz9YLgx6aoNhOLX8lsZay3lN9EVTzmY8Dr/5a/rEU3r
P5p5RCSDZVsZc+L50B2PRnuOOklwdrH0EEf2/S7u3sGfV5jM5Amn34yAbgGh0NrQ
kQhLoj656fg4fgRmKyb42gsR/6JLxt266C0xjb8wCQECi/jPRxm+mJWytN1QWAYa
rGEPmO+YfiWvBSiiU6lbSbMt9Ob/1KAOFdJR/7aVEJawpQzuk0oMkStvjkA9Pwml
f5LEOhQZqTM4hSaFfann+yUOrFn4x7UM75sbs03yPINRaB2Hrn63dmTKlqC2o4pX
sUmTi1WFVLIsJ8ocZgYbEtD/gf1lA2HY7ArcoKPxestm6Eu+VUBFfSGXge1cT3X9
PLPdfUoSdv5KZ2xfpg/6H3oC9kx8EmWVAMVd6yyIzTAfMe9e3WG7nF8PnxbtLe6t
G0fVG9yPjOe2Ul1t7CBF7u1cervJFuXjT9RuTUnGmnzHUFVRcmXjeiNVkeIhSmP5
SxfoQL+Kso1Ur3EbMIJcH8MXTkkmbloGVuGpI/rmJsMdin4/NkEE+sG02p00cMoA
uEPIlYz8itbKL3R4gSFejw7nNVxEDfp/mB62dLXpp3YbovPzfo7XLmIh5ktI17qj
7S13tHdRU3i4Vx6zKIx30RwLSOfyPJuQM3KBX0TYrNMH90W68rd0gEVtXZXtkJ3+
CLYEsjkZtnsQRnFgsV4+lX0PtDWNuyDyMkGoNR0RG27UVhG0kKVinK9ErbCOhldX
FkhDHnpirkkNKPJ9cGSXMLMEcPRaQTRW4xZDRU6SgdM77vFPaDF5Yw6yO8aVwEdt
w6/h3EuOAFO91moFbLJfG6hOAMZ70Xr+oxJnOuXJ+iU8PflBczW3Ibc92AibjtEq
kxjflWfG6pm1HRux3/u9zgK4UcSFKo3GLeTCvP72HjCTlWXvQH+QSuz0gXzSWpsQ
o3y+HNcHsSXzCSI2KtTMopmYkrtugB0G8RLMFstfsFmZ3X0tWkq0P9yQi6at/T55
7s+88ED4IffH8BiyY8Z/dW5p/XDO27OGqdynxg6DubGBgByhn1TLcV9+ehX+NlyH
Va95uxcM7LT0oOPYZJHVhupC7YpJ4BSbchRN/Tn2YgLgEycr0BxmznxfX1UdawFQ
sPHMLZryTbFwBlpGBWdaEth1boFgdywlP++LrBBDWsy3+whXIBQuG/G6ZsP+EGiV
pD8HxcT6kiBIW5W3nHaxmqtlEZ0Qev5Q0iS9/sX/5TnGlSsXdgAayV4rKdND59u4
/PaGXqIABQAbklE5IkqWFZMErZkMKYAWv27fMkmOsEW0DCIQzbcR7vXA0jw4ogJC
HqwGjHC1vZaCmXGTL6Q//qjhz0q5xEHWBpWGvNIQDnoqxkDsb89D2nrSGaAsOcko
jZL3t94K/yHU3+bFz9s+qSqxCKbVIekVHM3EdwZaaZrVKmcqXaKVnWr9RqOs5egN
z6OcThtpqXY+KQ7kQVkSXVkPTL9UIfYp3RrDfx0FlxdC2Joik0AhlX/uK4bbYSMF
KeYOlBxgPaqnxsKiJU7Y6sZV2ikr7/8qhtRXAqkJXYKXmyksBbq8KZSpFtX5D97r
jPBPRvxyBKXoGRn6V8kKZk6sm0EFCJX24N30Wr2rDBgUL91w4z025M5P9aHvLMug
i2vymGx/2hDNzHXSwXfS8aK3j6A1tbPSZyMGyJRulrnhq4eE+sx396YFEirYl0Cs
CqSZF+m3GjvW3G3XTf53vzmKlWUPKzBHyokSKlg/UAvTP1gPmo96moAFKoeODdRG
EqeX0VFRFRJTjZW6gDuBYQPNX9N7RYd68WO/10/v4iQM2ElMzMDOqTJJ8UssGG+S
jLa6KvVggjAlMwMAK5cRsc6bg7aWjmJv/63jnZDlvVMR9hp7P4Dnlk3ZbnMc2q5O
wfNnB+I93lgWK55z8KL2u/4fA7rNxDb97SH6x5ac9vSaTNon2ewuzh7PFGwd62dr
FfUZ/Ca8AsORnVd020f4jJjKR8bnKGi1+MLAcErPs8flytjK8OqUi7AiVBQPZ6ZS
F/ZGg6LP5desj1csDYm9vM3y4Xu+1Z2X2h6uGKBXhC2Nps0B/zlAipB5QtPUOBu+
yhOmBBr4wFUF2n6BYfm70hTyfa6Q2VUwJpYyhH2B0jh9zJgGuZhgZVEUKkwQy6RH
1osZH32VrK82EeJVXSqgoXUI+g4IY9a0t5YE7s54SWJFQlrJ7zcA5VufZaQyC1iH
L9UbNryOowGN8fuEyt8ioYgYSMpeiD8ya5hefrHYL9NZ+1pAryk8/AuJLWZpHdtQ
v4RW7Q+0rLcMrdyzcvSsvVFJb4UugHEWB7YFkvsvMsSLNrfApRitn5XwZzWyguaQ
odH9YNtCSm58EKXtsoRXsGLEMKNnxV1wNzAEOwUA1Shei5GG0vAh4hwAvAZBBwVk
4r0fB1SgGJtxPK3AA86d2iI3GY8PxABcFbhcIeQikctvunudiWOjirNVDpj7Di4V
9x0HRbGx41tTscpSGFG1q8EiSZu3DrVw7l+7VXkaT3z0IQXaSS/yr4IBG/5LHHEm
VHyERRvuWsQ3F+CBEWofe2pODRWzqQkk1v4tIBhELx2VepMKQ85UIbNRrJFMCmrf
8fN3BRqqBlBgrbyGxkxFiqjDUOoSzrnjUNW+Dc8jtLkK4Gll8HjPn+WNalH/nTpv
MmIikf9JVdtdEJ+wpuwkHxJKAalnYjdhnHjRWt9z+/8g9/yzu/hvvTO1e/3hL3Qc
t5v1AdhlCaOA48jUnRd2QEW/9c4PVecII4mxcPJphrfPMxpkBdMWvencvVu9bbOa
hfaH6bDcTSgug5lKAltj55gKxLuRQ/vOOHrbAuOQWfTqXkAEvIp67PhAAZ1PoQfH
B5gpSb4HmsxB4Pg0XRN3BxqA10+8/0G7Sf1ttIqsB/hbsZDPIQs11qz+cIANboy6
I1Y/2yvfsM+0pfWB7ZKz11RK/NOe4dwPK3JGL/rQeA87iSBKkSJxn/QV+zhb2xOm
+TP7FrVNtRuk0pIBGY9jLdnJOcBXnC1YKT+vXbdMA7tWNRmDBhh1H5ScX9pGxdRr
uIdvWw0SS03C2mMZcV91H9yljMGnQTuztuK29Ac8Sun7rQ5NoorMLVFXRoogwJaI
LiU6VSbm7e1ol55ZD4tYB4Rm44YDAmzk/Q9Tl5Du1hNWh2xWlGLLRv+Me0TpbYHI
o5MoKv5vOIBCDqlkOTxP8ZRs5ZdgIyDBvLb5Q8DWRVbBiMBDCmVof4R/Rcaws2yj
R7PyrkdBJwmep0wlYLZYKMt/flSXQS6jXPB8K9k+L97Zdo3RKzRBm25cpQGmlinm
320lAvUyh65oNlSSAI+DyuLYHVrzpK2kPpHAZjiRGJq30xHJbhSvSaWfHmxM+IQg
l8BhTu1W4mcLNMST4Bs1NSFZkvo93DP1xlAzd/iQEYH6BdZI5vsIBs0mJcKQNSvT
zoJNljwOrkU1gkfzNBHUyByOir8KYOdkxYr9k4T8HXQ7wIbPXFv1vjR6EcqY/5yz
8NcYKilM/tY9kn8Nq/2mjxI5MFJHQZ9Xr1fkx2Ym7Wd4Poy3Q6mBuOWO9FgvfMdg
/ikqrrz52OYGoMUSVaGmB9P6C+x5KExMagJnu9oYxcHOXZjpGtLVgR6aXRFVbgTI
lQIFRiqm38IwbANW7FyL/PvjEwf87MutUTscr4MP/WK3epr7NcYBrTOzyUL6Rffl
lQXR2O/2ojZWdFGcMwyAuymX9wwi0tndFJJfZiA1SMbjS/3ItqGlLCfEtFs5rUTo
ZFdU3dI669Le8v/yZKxhqgp6lglAXFQenXTrbvGnPkfBbKDbhVYpAaIl4KnRbKzm
ZPP1YwKcNUGNqEA1+NxBcvNYWuisasyBiuvigJEP4WH7czX5qMd5zYXvvHGqVTon
6azyIug1ITgT2mXtBAdj0XTia7yrV8LExYELRLbxhF8/fTfKnmlqbaGIUuZhtedB
lD8oCaf0RMrQbT+Evi7izjmMZwvFWggYp6xaRVjzuCFqd3iiY7IwisPY7U/EcSqo
nktKscyphJYD4DSXaEPuRjkQnLGL48yJokuj5NbCd4Px1O0WP7Sr+RW+KaqXf0/d
nXQ+45MwfUYACf4SPdLcDO1VlQrWwdoOMcg/eocO1GFd1m7IOyqH7h2yUdi3ShKK
qq63aM+jmGWvSDV03HekmLyIwu3xA96FfuSG/sB1wglZRGkI/SW+5dmNRrnXPMn9
gHnNZ3d8sorf1WppcPMfzI68NO4PYJTA248mNSSX27HD9kBiqTP5otMhguYu3VYf
3o6Q8xkDwVUdcPzdZRDijzgJV86gTv5R7TES1OyW+TH9QFFPvdv8TppV9NVuvAh9
/pi6KfLLNpTWL5u5JrJu0Owx/AIk6PPwSUD3I6wbtzVJcb7EIDJ1RCAewLGivy1N
IjwkoiPvBGV4OY+kLHG+SRhGlU6sbgYwB4vdhVVPS+P/x0YB42t8ooNgNFFy9e21
tl0IXxLQZ/5XUrz4E7Y4wA+6Dl0tiiLRwui01yhHIX08uyiaCXY/vVHdWwZRqsO8
aONILpgMgIVN1CmXekVTFIKBCmiRbYCfly9rURO69LKWkBDLSzdNyO8nqBGx+uz/
YdiIPtGYBrzGbxHMh+oxLi7SsbcT3nLfAt6D9CnoOnbQH3a6zb+Vp6ufzBd27d8i
a3h1eL2Xo//U8G4dFziElTkVCditeM/uTNW5ZYKtgDJHHykChChsalLgNLxHA5E2
fGZOp2fZp0tsemls9j0uKnPI5PV1Xn7iOrw5LOu8cQ7ejKrxNtJU2nVc2d73JFuO
73Yn9ipjpYVZZvZ6Vs7JC0frkaKogVW4/uuCT47eGMR+RPxE6BPWPTTBsODTHnug
/mtch3oCMWLlcoxwH/Y2RzK755KsQv7vvWy+aYr68YgFtbaSZa0zwSvF3JfVVL2R
JUnWTYu50YrWMCsPtgH6BL2sNZwxgGCyuxdcXRfzIa2nwCJU8Ml1VD6EB1h2iCWA
pNlIIFtaQWctLR01cGwXAKFXRwiWtBiihu1zNCmR0KZ1STJ8uosDfegW1g+8K+dK
/3zb3/zy986bs5h/YE+aXWdaiPvMzGF1+l+Jhr22M6Ub1/tG2LRfLUX4WI0JrYMa
p1XUd09OsSXBFt+ZrYqHj6nfDvlSW4im5p+mVo+q5ovCxW5m1k04+N+kooIKS4k6
79KJ3ndrai/yP4G4F6+/0VPHUNrJOCvFACveO2/vjWkkX7SirGM9Yp1YDJ7qgpDF
v5QPUxZ3ZmhAQxm0Ss10QBDAcEATncn1uxMwKQ7gInXq8/TWNT06YYGFyt0qRret
ddjhQlR/c6Z60Xm8dCkpfXZIiryZ5aKTQ4c+lk1P83Z9EHUKQLasX5OGsLvXEieN
Nhto/DtxGNn6+OJ01QQ5A/YkP468p0MJZA/1aJwsVZpvC32DIrNuU2LOKaSKcylk
wgwyCVlRsAbacr9GcuZcAVc/i8hdZ7aD8ltVUiQW5rgScncCL+FUnSusbP2p3QkZ
JTzVln9yiGdCqbWqzjVWqM/yvufSyfkPUENVMRUNUkDUYth6hNWUiBq4xln/Xmo/
Oq5YMD50TPCpP7iWG9KIbJ+vuzSOUBhzs1CcuEWesb7/3cfivvv+MWVa0sOD1Mj7
fygxD/+XECo7LomAC2fj7yXOF+pR15i/cI0FJm3s83AM5aFxYU9iN7BoCfsX2qVm
1RDySQdQZ3MVWr2FgDVHnYQCcTp0I5KBpB/wbjYtn8lqCbwYu0/iFgiUoa3DxPVq
UxO9tz8jO/16xeEX692xlolWzcNGbxzmT+AZrHEHViYcwPrfymYRc9LpWo5CC4XB
K2jhLMPUaKutLqUlHYuaG/cpyiBwPHVVqlxR1TccBhydyowal7frA7PjWh2jxX40
mVyfaxSxZA/vxu+MO3sVxpUfY+1eA9o6YHU5HBrjSB6viZoK9EoqDTAM8wjvDvqa
pO6zqgHdsnHL8c/neS1osWm4bNDO9hlURApcOkOv+3JsrOSfkwbejN//n3VNy699
PmB2unfC83bjuPaO8UdxjhXpmSzhzlaTSZ6JWf/9GTTCScFGrCVANuFXJw16fTe+
5Z9EdNqeJ16wXl9vw22/+Ydpl7YyBsK9szu+OEEkknnyHqxBMNqlWnZPxt4gRoyL
1sXrjBn5Z4BWs7UKq/OyGYLJ+IosQu8DBN954vd18GjkvtoYPoWhMopB2OCb6Hp4
7Yo81ZH8gAmvrHBIQpet3xjtf67zCWAP4WSCvexhmAQec+/UAJRudxq76jatDbVI
+73rn7RhumIf3he0MYstfI/RM+96MEGzSPVvgU8LyQsFE7VjpRK5HymjKk5umzsv
DlSTlwEUU3udBwMoTOlkS0ijRc58BJ2BBcJRqvcqXHfyRo/SaJeRTnmB5SAOpVjz
36tQQugEI7y3NPMKTsfoBx/jIo44ilDhTiwbbebu/92krgCWJhjG3FSVEh89BzFI
y4sd5ucpeUdyLHN/R4grxwTBdoTFRJy+nI3dGzmehvhBHv4JKlOKsifWzqlwh4kb
MpUkLM4rXR4SyA8k46gacE/DjwxhmkRU5JtrqICfFq5cwhXGcDiTfjUh/JqiQ7sY
X0rG4UB3m/7bNcQ/aV2d5cJOuEU9TNegk44M01z0GfqTakU4g1WjTug9GkN59NRx
ZfHKDfotG29r+dw8h4RDzP092FTN6AFB5dJH5RJtUbZLMO8UQXuF/rhcr3VfVnqo
9ym+x/HnzONumMSunRs81PuUMgsfe5MqUgY8ZXXlMpobLXvDrnRU54F8ydxzbQ5w
Phxe/V1DSaU2wxf+V9BiXsL0ZGbJGrgPp9eDdeAAIeUVBKW0qsU70sxHZ/nhUYra
ac4h8PbCZ5kRkR3H6rel8evguyrr7FVmE4Px9LHw2LYYUEZhjn8mA/7J4ob4VSx8
Ia5GNAcKeReB17Gm3qDufWItLAEM/nKmBI8AOswbViK44lmkKQG4e3ynAuDAHmOB
rRj0fXGzgEvxgHwQdWgjSettWp5N/Op9ZjdKEM4/e52OiFyGLCoyNQcs8cRJop+V
9Tm88knCnrGqn7RuDgadufFjmFUHmIVAKsRjT81ontKOuoG2h1A0pPbhj/BAzhE6
qp/c2Xvwc41sRLtBCljubXl3SHf6bChYAPJiuwYC45rEYxPSZorrTBXUcjU4wBpw
ucXXY5LOc4sNitrvveYsgl2ezYLQXC0EtyH6S+j4WZc0g7afYj4yyg6XGxQOtZjd
8ClbZ4600Un8ToY0DUNOX71K3N9oZ6tTECZTcfj49Ym5Ok/8fS4akz6ms3aj05Y8
LB5/F9bDXyacsnIatZeyfackcMCNfm1hCIt4k1vjRpKIKTN21bk+JEhHnYzalb5e
zmK3QHmFp523izHYnVsC5Z58A0KvddnJOsEvlHhun5SbwMtUauGJX3sK6osCu6kV
2IiolvYWbOJPb2MSfBaYq87VIKuuYklp8wVZwxc5UwjNoFT47P4iL4Xh6asoEQi3
c1+yumXx+AIatjJoGTwTJgqWPnZDbT+mHW/InG++i+ADHqAT/zqJeRLH8MRSEvDJ
f5toP8pFmsi0fIw2Zgj8geZMTKk5J52AklbnjocMsEOn9ebiCxCjgCx2Ik+cabj8
51yKuEPSyxPbc2+6rI2zOrWLguSq3UFApwJ7mH//hBy2Btmq4M7jXIBLyrRT7/gB
Am8e6M6oixGTQrdEv0CNP9uDxriBwtiLe1S7iVthZS/MFvf7ovwlWlHccAfTfplL
uY1PkCdpiXv9pfceBozrWpnQMUfpqIRxIl72AE2h96xj1k1RtfOJYdjzWIrTZmOZ
eU6pA0sAGXfKH/0XlFd65g++8FJmBkvHd7tjcWPvZ2jgTV4aYYJgr7zG/jkaPZZM
FroNoDF7eX5JKnGknMwPHEulRSz8j//Pbapfzyre0q1XjYA+a/r1TYCvcj0tnRHa
IDW4nFWJwblZ+hN7eUR24G9ggZEgLmZUqC38hzSil1c=
`pragma protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡j��-��l� �3Wʴ ��ȟs�/�\�Kڰ��n��T%�ږ�����#4����*��Sv�=~yQ�iy�$��w�2<���0���xoV�NFE�`mւ��פӈRqS�h4��yx��7AI"'�!��FP����:sK���8�1�9:L�Rv�7����M�[�3X$ʦQe%�GA{�DN��� C��G�L�U,XWNkA��h�x�Xq��f_[�H�Goܽ�",F�b�����c�	&�ΔG�t�E��;T��0�v�-��d'N-3T����k�Q�D���uh�2�GW6�F��F����mb�)#�ʭ<�+Sa�wY�e��Np >?��GϊFYC����ܑc�p�5R�D��(�e�8�4f��A^�\�������mv��g���`�E�j6%%;[#�)^ik%�*�>�Rw��������h��rm����K־��q*����."�Y2z����<�)u+�ꕀ��M�iw(.�7U����نS9�meS-���dSȟ01����YE���t$t7���
1�,�")*����`�.{��rz�86n'no`�~�6�d2��է������y�r��,� �}��W�C��� ~�µ[�U�8{o�i������H�&�/ZC����As2?�P�����xұ8NP��>����ݶZ�~�lґN}vT�Ԙ���e�jǗ����M����k��J��&.rɦFٯt�7&�l@U�\�Ʈ�`�di�FE1�=\�t3d�)ǳ�c�/�֡�Q�@�n@��]�_3���]WB���GV/�����TAm@���BV�q�Kk��ĨUB�Jᩊ#�ư��T ������r�6/_��̥~x���)�.�w�;Rl?��f��_�꽿���Q2.�`���d��z��4��fe���L�5$�E�u\-���&d�\d8E�1*q���z��":�t묶^�H�V{{l�π��Dd�6l�a�]�b;ь��犨g��Gr�lŽ���1R�2���A}�;?:vd��4M��٪� MH��ћ�,x��dm~xC5� �N�2�	����k�-A���a4�a�n�4�|��_7�ޛ�X7ˤr�+��T�մ�돎����3���sch��x���BP��vr~��Ny9���}}�щwF��fZ�tȂ���ҁ�ś�?kp���ɗ����:��Zb(�� ƭ�q�y���H��'hA�uC�Sx��3)���_K~�8�ze��y9�,jyjS�@�f���Art(b�����}�'�>�P�Z��`�*ЇU�Cj�� ;���r5Ju�Ϳ�)���uEʐ��5�>t�uw0^�ˮY�lל�c��Fw���Y�F�%E�<�`4c"�I�y����I?���;�8�#�����8m���`<��e��O`���
a��aK,��t�7$
֡B�|��� ���ܖ�
�(��c�s��Sz�*_m>���J�\S�sD
	�I����䜳 "e��]SZ���	��$`����7O�?�+�jZ���7�K0�Ϫ�I{�X�&�����V�`&Ǐ\�k#��.)F��p��/Kː3]z�<wlה����{H��C�ۃ��/,<V%f���9�<+��7/�'�%��p��!q���9YG�8�/;�s�cS����_Վ� #`(�G�+��Ǯ��[K@B���n���pZ[����HA�E�����8и�M��6�5 ��?z��F��E��U�]���H�ˌ{l�ʥ���|A����wWY	���E�r�?�'��·ם,!S����v����k	�@�I�m�t�tC��X����7�:�y^�`R�h�T���`!u��F1���"����qM��Kq�z%m@��G12�5?��[�������*����t�u�Pn���%1��8(�}<����+I<A�Ѕ���@�xU��Z����'��H��f͊�$-�<�O��� �a�@M"/ l�N��âJ%��)���������!�͛3vdRvt��;Pd�-f�0���:�Pqxqv���En�a.��z<u{�~���0V�F�C��� �.@�]���#:��M�--���J_>0i�qGR#B!9_AC��c�~�(���(9����lƖ�K٢隿8[F�����˩�?U�nx�c���Uj��IB�u���2�"�Z
t��I�N̉WG�kI��b��\'�%y�!�����	���Y���-�eo������_J�4��B''b�����3�Up�}�Z��J��x�l�Kc)9�47	�\�ힺ�&�cYo�&<Gd#�k^� jU #Φ�I���$CF6� ��x*.��=$m&�56�ZJgB8����i\I�ɹx0�ʆ�+�����PBM+�OO��z3{��6����f��d�c�ix����k�a�oF�e�I�ah��|ɤB�bѧ��.��.i�)Ω�C��?i6�� 3*~~f�\1rq!����� .߫%��E�������E�6��Y������rĈ��<��Q��#� �}�?�VX$��_�(�hp��u��v�:��Е�,(�r�b� ��a�=�k	c��kaۄn��!�@Y�%�>_��Bq��j��Z�� ��:�!�Z��G�v^�};�*UA��fw�z�=y9K#�ג]��U�ܙx�Al3|%�!=�!�'��d<�#�PN��Y0���$o���n����V�f�Z�����)���������r��k,��R�6p�H�1"yB�В�6��D25��/>Pr{>]1�F	i��!��Cuo��HBD*�)V��+a��R=�;dYD�b�><e{���S���lk#�t���u@ؙ𭥫W������=bt1�wX�􉪫4�d'��Ŭ���"Q��^�y{�︣����߼�a�ɾ(����=s���0d�4��� @�bm 6��x�q����a���Lp&W����(�1�#���:p|�������(z��ݛ��ȹ�O���I����Q�lR} Y��_�Q5L�躝߯.��W���R��xq���x�?)�oM��ښs��ԯw;���on7�V�h�SQ,�2[����l�&כ�w�����5��������渹up2�9"���j��̭��z1_�S�.ʉ��Zy:ǿ/�Ł$;7���kI6��=�1(�S�T��8�/��� w�=z�s�Ծ���:�|k���Z��Я[�5,�k�C�w�#XdcP�	��n�Ѣ/Ύ��z}�y�j�(������.B�3̼�x���2����v��l��c�4^�HS�\���2�M���V���6��HW|5Ù�od-���0yD<�RdR�,������ >�.F�f�G�U(���&S=�(�6~Q�mm�"�D�p6�Ѩ��
/3�ů����9-�o�]�o�|l9!���%f��4%����Mj'A�c9����m�mбF<�QL�*-+Q�+/�o����֮��!$�UiV�b���7�vAv����tX��ě\V
��7�{���=bq0������{�5�}2x���S��4�Dڹ�ɤT��&a�Q�G:KC�C3',�6� �������Ll+7�7����!��5�Ǥ����U�L�hQ���Lq������jm1Z�xԄ����)GN�J]ݖC�������n �"	jD�c5��)��>>`�@*�6��{��@Id=]
Ã�N_�Z�b��1�߾���g��z��z�=����D�������Q��^s�=�����^�2p�B²��\�A�w�xAkc�lA�����,�8X�u�M�ƆV�K��<rN�J�o�Q�MR�����˔qo�8d�����	���[W2���qHҕ�m��ōD�c��-��o�̲")?�˺�-p�D��Փ�߃T	%<����/��~/��K"�2�v��m���4�%�D�T)�w�*�z�Y�8_/��X�)�`����M��R�� Z����1nvjp8������$�jA$�R��w��UD��xx��fs�x8�S���>�|�:�ʻ;��[|�:VATa���Ky�6��u��`����3�b���%� j3~R�-��РϺ3ȿ��&���^y1D0�T��	`�'��3�A ���h������E�pEDm���GΘQ��^F�DD8�, �_H4�;DJþv��R'���v��m�� ���JL!Y�P9��������w�/vpԜp�Rp��ñWmU��n�ҡ$I��H*�����Sm1m�C�,�颫������ܶTBЅU̍X+��!Z�UA�{ܼ��p��_?V�F�lpN��:�|�\�3�͒���9)W�s�d�*�PI�����ֱu|�cSʸY��q/���쬡�z㽋�:���$��������?�v �d9�@���%w$�"�Q�[��QM��o�����$j-���`�*�RjBc�	Pvrm}#��:g��G:��)$>���2{��7�&�/|�.T�������#�c|�r��$3�6E���>q�6�\��u��&-�wul�`��(�+���->�����XJ�O���h����M��|�w��,0uy�aFB���R:��8޷ 3 oAe�.�����]����8Ľ��*-'��N���ܣ+��"f�~���c�'��k����]Lk�R��-�m�$���j��'�.M���D�;�㯝�{S�1�$�q̍.@�f�T�����^ ��"�و�n5�$����BtZ�������S�Īn�&@NA�f׵DR1�a�;�Czեbe�/��/y괂s���zW%�A����6g��SPu�68F?�b>�itO�F�#Ub���2of���2A��}�S��wToR�},א)��B-ิR�%M��Jұ���5�O�Y��=u���$y2���0�	2�Z��$zW�n!��F{��Q��ˏ��o��(��$��@��
���U�c�{���m���x�
hso�k��z}�\-�Հ;֍KJ�y"\�4��K���#?���n! �52�z�g�7լ����3=��R�9�'"����$����Ѯ
� #%���t��Z�;?W�WE��8^H+��H�%��"aU!�}S���iK�3kc(��m���*J�+�a���>L���oDG���[!oI��"���]T�s�V��Ț��6J�b�K�O!К>��z"+5��.2+i�[N7�Bg�Ggwa�\��Rf
]������4�M-8c��4^}�(2��1[ಟ�*9�\�<���8��/�ħ<Zl�)F�r+��d�-���zFOy%3?93{̅�V���9f��w�Z�'�/fl�)��E�K��!�2d��$��,*��H!p���;t��]߆�a�mCml*��m�я�B�\�-�S��=�@O����	�g�+�>ĕ�
�C�;�m���[q�J�pW�-~����J.��/�>��)�.&�!yU�&�v���̊�j����-�9�mg{*���+��;*��# 7�sz�Y��Jc��V]��ymdI�L�SN�ʃ�vYR �����!��6�q�Pg  ��( e�H�Z�a��-�N$LY �ϸ�z����'	h�NM:]���߸>�]�N�y�Z�s5��N�vDB�C��������Ic1P�zZ2����+D��G��L����Y6�&�0{��Q}C/E$�`���`dhȏ5
��S���AAwx���'JF3]�`���]�ኪ�#�c1'�t�S���*<��B�j�a��?B՘K��4������
����=�J�����A~���^n(b��\)�sA{(,���hj��5�;��9'l�ʶ�E��җyVgE�]��^�J2=�wq�@�R�M�̻���5�;ќ�53�G)��?Gn���p*�Et�����dy� H��S�XKL��%!8H��P�M:Jk�F�2Ә���d,�D���o�FJ�9���[_���n�Bu�k3�U�t��-��z�Q��ˏ�%c,�\kZ�_pi�FH��h�&��8��l
!���C*�J`J�јn�d]��z8{+�� R�Y����#5y�}�B� ��V�<��~m�UԞ:E.�ǢY�-e��x^*͑�qy�$ Yj����E ���ZD>��,�q��U�����=�����\�?ZO��=�x��Ru����Q���n�;2��ּ�pw$��a��Kl�"�1��&@
�6�?�o���ql� nԆP\�ޯQ8�g2M9�)�5���˪Af�GP<r�]u��AX^���u�:Qj�gu4��P���z��S�g]o��UV�q�i��*���CIR�_Cm�V �R���u\�����;���`g�+�/;]�PЎ�z�j�6�a��+$�=§����D9�N����L|L׊
^6��t��y)U��-�=�H����2Mj��|���@���3�CU��,;��������AL�tT
x��4��u�ս�/P)�w$�3D�\�9݂vgן4����a�ʴU�U�����������v�x�ֲ��3��K�>Й3N~�KZQ����pvJ1���z;
�1��'�}bG u��q.�U��6qZź�������L*+�F����es#S�eO�O�p~pmQ2� ��֘�-W��~Ҳ��Y��7Z���((v�%B}ڌ�Gv��i1v$��s�&��N��q�S�;��g@�#쨅������˾8�J��W��ȓ�i��*���zO���o���a>��Js�+��Kň !VJ�8"2f��8Hc7�X,�gJ̀H��Ļ�c3��k��\�: ����:嬦=��c-�6��>�Ep����d��/�L����%�G���S�@{w#��E�~�(өIi�=�$���g��h�3_2�u�/�&��KZ�rv�j��
��T��u�ou*�p��^�xz�ٌ^Jlz+
�s#c���RX1��Wg���H�1�]���̐|`$m��l6��vkB�0��ezطnSa����>1�-�d����On��@*L���]{���_"���bCw|$/�e���7O,z z���iv�uہ�����l�����c�ˊ�����ʱ�����������U�:���3������îjF�����1Y���L2ý�X\>-ŵ��(�<Z>_�(�6]n���6-n,��P�Ҙ���F']��\ ƾ��9�ب�ȼ�D^�`�?*kZ��Ivy=&k�nƅ1�d�-,/��ohk�>���l!�D�ο0r��-�$�޺��Ҏ�����A�{ia�U��
���o?�0X�;047�{ǎ�f�+�x(��VG=j�����{m���6$��M�����ѣ�l�H9�P;�Ρ \F���D�yl�˰�#�ΆdJ5�ؓ�����8X[ѐ����x8U\ކ7������m�F�V�|�v������<�hL��J ԛ-�%���bT����3#�����"]���O�{{�O 
q�Xҥʭ�O[�o�L�PP�'�{'��6Ŷ���6����=�I� 2(UC����!_����(�i�)CK�~n����8�����:���Ć�|0_3�S�GjdҊ�
��1�-NRv�]���"��ȵ������U�H��߁���q�{o�,{������1�\�\�BfCo]c�]��NK'	�qc���� D�c+��J�T.��D��'s*2�@1
`x����������l|*D�i�!�I�T]�$+��q�*�mp�
��8��U�d�{��S�<3���J+=O �O0�:G��mA��[Ƶ��K�uCE�pKB����"�]��)-�&Hw$g��0^�15O�L^k��[U�H��Bl��,J~���`����ɋtũ��ؗ9��#T+2sM�R�	���U�M�(�K�E}Y\�R
$��C]�~��.dK�G.���Pn`��o4�=}�G�~�T7��;�P����G�&�F ��EV���DF=���Tj��,C�)�\fՇn���e�"Ç���"�T
// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:25 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bAFCMmOcVNrTL6Oih9DOpPvPQbGwa4KT6DzJQQMUeVr79ctfqP9FKqdSzrv0jAyo
5iOLMMBjJTglIiyeDxlAGk7LQNrPX2QAWVEJR1zvFQprCYGVE7ZlkzPQMujMMlsO
izeHLxkjSCkQ5NYhXIGUD4iacgmEbCpO1DhCfFiQOVg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
1xeb4eVd4v43J9i/1yWwcPxTiqhcqFTuPYjGEfB8JYsPuabBhoRawlz061NFZ+CH
Iebl+QE3G/sIFsjSqRDqyh+Klvipuyru83iG5iwkCqPdhHCCcw/XAbux024wjoD+
ikkVzY2TjCx2wO4GBM/6KXgeN294IUhAGrbLVL8zrckWLNzvX3MK51d+CJYS5hgP
YbBZ+yOzS7RJL5ZUHvEqLYKHVXeVb5K2HSeQcFb7vbP0gECsHezZYQxhoYO4SQDT
d66Oi7SwV2Mi1NPdXf8YMRT1pzERdN5yHaPxC5zI3pLqUbbl3oiJAOwO+MhoW0nS
lzuivxGF+3BfxAsJfJdSPdEfGHLulcrXfqW9AHi3E9vpIpo0OBxI3C6emIB9w4/h
HH3fZ6CGE9gaqgeQxiTIiyF1ih9VWwDkmcMvKrZseWYRXhtWEnh2J7yEXpeF0aUg
ALoJm0V9G5frz+e4eHLSc25rHFXfmNrjTi+bmoNuzKfCmf4tsfEDWM8wwLUL4phm
G0nDTYGi8agHMdLk+2rH+D3wt3pFy+/rM0WImpXZON+NuBcQP9usbS/jCo+UqWXc
d1tflRbp1d74mOGrUPNTG/n+/5AvZ3gGBqcFufpHA+NfmWLWoTgnDqSz1mp4aoh9
Bg3h2Y6oDYELQ75SIRDKIIBlusZmn+wCBhViEqhyJUw6HFlrK+4IIKuGVCl/rA9z
IAOsrcAEYhWlZwIckH6T1b0HuYXkHQ25ZtuAcBTQiUklB5MtTdb8mfWRwNNYAlzB
cLmrE12SgDe4WVvivdv+m6fBkTUxMf/1uJ7XGjYudYrZN5EScsBi5MmcM/zIJp1Z
HNYL858wCgDuLpV7IGTZXuB4i1pTK5na1dwffDtMbh6p79WyFRxMk3gRxgek6Ahk
PIihIsUh1wyrErgELlS7ii3lYZo+vI9NnyjB3htdbNrOKUrZT8xbbg6rd8cNejlP
CF/eQFyyty5Yk0SX1lN08/BzcIG7e74dzIPZA6VaGUEunWxYVd3DRDjVnxwZYZsu
hEwCfuKAdS74Rmu+mh5/Ez2RgD+c0gt39QAHqZjsC0CSgPH3Z33DRFB3NBst6qek
izG7YygWs9oJHNaqkTwKt7QHWabdbQo3Mrr2LnL35ynw0oSbmHXztdF8hW2haM1d
Dc6Nn0GHitHi0LK0qvVs2odFOVz/NoLdBU1OVoVGBsChd4LVQ1p/5Ju0FeQNQoTA
rg5g6d7M1FJ0Gg2lsEZvW67ChgCpXlJcbJzfkhEnjDA9r5Z6J7nZ4HYqrK2wmzdh
CdrDmp1O0wtHQb85Nv+9QFlyObAA9Fe9V20uhHoOhOdW/X+w44t7tzwBSUeLWRux
/9qKfJ5sfMWO2rrhfRpRB6dSSiZUWVOMHN/McaaRL/Vain/sMTWqSZgP9Lzecqae
k1QJgltoT6IZ9GwYNZKqbHvnNoAAA8fI01ZB2ykdC/tiAUyIboPIHgrQiT0JaGhU
/oNzx1Z0I+PiiInQuk4eu1520/gvnq8cmP8dyYZHA5Rn2f79dKjs+9LJSttsSg8q
Ta1vcMTidiSQSxz8SpFRwv2ZLRE/ymTrROuvjWuvy1INrP1GMjwIaTTr8EhYIDh/
lvnIfwhi1PW7VxinS1lZF2pssEpZkwuvacx7XZ510RX9gU6werQk7+BFG5bg9BMH
jB5qfScsMFyrs93WRRXuZbGIiNzaKI1M9z8Fr5Mws579cD/VvFbsEPSu7QBO/m9F
g/dKHqTg/+GxirytvL5FwtFXbD45MP6NIR4qpX3+7vU0MFdAC+1PePQhZd/mupEW
Md2Xt2ZSg4LSkyULDps/s9fm+9JsCHE953/TQbqJ20r9h574SPwf3bHO3EO2EVSH
wj8OH/cgoHDSA2ahh6oj7f/bKejWU5io8/Ms2DjMlMW0dusYf6gg8k96sUfwFYPi
swe7xlv6U88o9bQ4X28AuzcURMf05SRETXvsQ8jUiUpakiZwmhhin5oKjhC2zWFN
w0cvoInRGDDzKZBnMmAVaMes7PQ+L4aGdpp2ZHvh21+xKzOnhC7quz9N3ser2iBw
Mvw99Q1r2Fa50nWBg1dv92284vmxhIzkogQXsSMKouQkE6OhYR+pkgwurWhzii0/
GiF0/bI1TyokZFZr/1X63Tnz23GOHLxpIPhpwyuaqd7uqNgsg3GKnTRS1ZsP9953
NVUusrrj3bjfJ6m6lSZTzQ+QJ0uKSa3FCcDjz92WGEf7ejBdIhltIXdWiH6dZzHe
HwJWQfAzIDDjzAlRXfIfrldi3xS+hoxgUGA7kem6DOmE7Kqejef127vdG4b1hagl
ETyPuZ903jGOVrPrmS/34UlNJwINptQ1z/PPe04R5ugkX7Opcik37QCkaSYCkN01
1idOvgRifMWpGc6BXhmpWnZHgniZbBFpm4FNjkYMHMr10/Df2j6kq2yl+uhCoT57
v90gXceUb6sNH8lSSDvM6RMuQW4OPPTSLfpTWUszaLoGWrgvufN28t+odjL/sqAo
N2ayC8xYziunsz3yBbsnHx8Cwf6eI+Npy6qsiWRNawWvBE/v85SXZr4tDy2fM7zK
PhaxVveSkm7eSKRk2zZXQ+OrQ/yzeYhgjoYEhJH89MoATgUhhs5mD2crK1PaCSKA
vXJoGKuOaaxCJ2a3KxIE4FGV3BZAOO2NY8uZDYvMJjO2Psje6yWKuBYhtSwd4Igs
+6fq9ekPuix5GcJPkDtMH4TR87wpE5bGCYIgSMXJhVyi5iKxhyi5GgO9NNMtD7mF
EmPAexueUIlxe4mSeta46VRO1vEbt+S+zhAG9qwKkyRUi7ybHXe48eet5w+rQGnN
TLhrBsPxhOVKM8SsCZIeOrnqZa52POfAtWix8ncg2h5e8FZXeRWcqlUnTdPM2wsd
k6J3XhgaeN6j1EWa2D/GT7IecJH4vjOG0QhySQOZEC/xrwt57MQCAoiRCRGZNZwv
BNIw4ZDE/zY/8VfkYN7IXAgBjFRML8MHBY0yJV/xjNnqeliCeJwMV2ZtlLxt5Gm6
1NyAW+IbhFHqw/V+8OnmCT0X9Prja9QyhmGMaAp06Pzjpy8h5fZK/lwEncTK8kzo
5ZkuCZEYWZx3Mv/JXtEsEWd4vtYfl4TWG2H0c5iwA+Vb0h6S5vyx/LbOxv2ltm1y
CVt6WhevR0bL/BipdGLAYiz9t+JoYAOBc6H26Trq9MT0F/AciF3/Zd/2/A/PiXS6
+SL1vYwqCPpH91ViULfGR1Vw4ibRwtNBQ4PjjWdUT/BM0QjQHX9Kg6XpBvWErMbf
W9FB60KSX/tu3IPYu9ywjsOi895xnIet7/RQfaOPGW4oJHmIS6iuKmmZ519eAQwE
xYSN73l/BOGh4ZTOGVx5HeCv0vE1SAZhRsRspwli+NeN4R7n1lqYKpYI5oX6qZU7
8yOK0WSMLy9rw3DKRwdXaFq2rQcR+7S1Rm0fiWIXFVv2hr3SLl6SpX4IlzZOEHhz
jQ/KI2pC5dDQmmWrG8IVCs7iNK8VAHoCyHNPf2sUa3/awyKNqK8UA1KS2xaciAek
etxpTHYNrtCDDMVLLxPV0TDtsMdcHOOW2eoAIU5LXiUGYkvCw9PjIl+G39YTyLij
rMMRXyMwIvMqYCar0ksfqPbt8AYW8nM/TkNxLgimgtyqrMvjn+LQiBLxhk32Mqkh
vZ71snhEtYnL73nulq8Yy02qu8ocnaO5bkkgAE5QCRFAQSKYWGbGkxSSGlM0olLz
tA2H7eDx2BrCqcFDP+tF+JaM1SkzlBgXn29zf1l7u4F8zIWGFUgXCOn2wo8XsJPH
bnaE3YtHRcr3KU+2qU8+XA7tJcjw/BTTKv1uxKQQ7hAuBpSnYm9q6ojKhR8AwT3y
3S3LDr+3lNH23UECS1tRUiDPKJ19oz+BTnPCOcoXv10BZZFbtHZhimG+g1LKTVIB
ze/t9+IM1UBtOZ97WVSQRXopbgVSI22nie3R60UU18S1ywY+wcEl1d1s2XUKuJIJ
FU4CkGQ9lnGAotdQL+JZ/tlca0lUoKXb5navXiRosRZ1HODM+SCZKXi4vGCy8Q/a
LK5Bjs4ZBPVFUo+rm4nZ6gFnI1zqtWcpP2EGsoZJkNJX0vPPCKTeXhQk91iPO8gC
5qijAkNYFz42XPr4Lvt4+79/QLjPWGdnNP3F+R7e+VIpW77L+qE8Ei/OEC3VuRFw
paixo9mQysX9Y59ipRINg/hPg2mx9J4nBLZTHvgdtXO72F40+NDzZo8azEtRyHUp
UcOftesxTZXxhdYriUGW/xNI2gLsB3DYD2Qya5GE3n1QBoSgqnknrfNTHtmf8QP5
xi0Vly27c86zgmMyNOV0oxJ1kgHUYR20nNzIFqDYLt/u2y1r+fpRZl5BswwM/253
DhNNlG+2r6vbubysSDcCIEn+YRXKEjiJnezQ+dDqU3yzY831Qb13mc02Pbvh7Fen
/jJEaiHaATMHhJDzuJU20WBvF+ElTt5b0v2Cv/Kh+YeIRcYRHrHFRed0YG5tr2d0
SYGe5K4TEG5aSqOvcoSAP+HVs/9Nsj2R9XiHmBIqj/DlXc4OQbkeCAfcvEJJnSKt
IdtG9o8fo3velcAZZWgYEiwssuARJQ7ciwzRZM/XSIRDRq0p8Eutgz5OZ1N9kB0A
s1dREepywZxcX4wygzHtZb1SbVE8cUTJYYtYKJJzZAGex+GJ8WgKX8pLzksrETIm
rhKKvUA1XTUdh11BjBfC3XFD3oDLIOOx4xx8msrSzLJnSr8YfvZaYrxmAndcN2C4
jD70HS46Q+Ext4C9cehdyIkagL0OT1XfMxmv+l/JxE9jqCOJwaeVf8Mf5ycAVBL6
7eXl5HR2ecNRKnnV761uPyKsI9FwsLW12FYhn6KXZYZ04Ms3OeyemFDPEBhgKRvS
EvPdU/jx56KUKNg4DTnveg3i3blRND562xpwyuNMNgE5tkg7bHROIWN51Qs6F3I9
ZQuywA6y56KjrydAICsukPpyz2ga7dMh0iW9Tuhk7+t4immFgd2kX72C4K5mfhkh
zV4latkbqOvNc97XYkKQrsZnPxIOjcXFLKAPoGfBCE63zTrhDHoeBFSjdWsJphjH
RmTLIlVyroK7F0uGPAes2IKtzBZhycEvcZVWrHqpeF6bkvu6UOkfSXMWF+NgXSEn
iroZKbvirm0UPGaeU4YXxagqpc7nq94I/dthE4N3KwtGX8v9itkOWwxzQbsGrTQ5
aX3vahJisaX7hMwZvYbNF8hBb6UpTYi8oKLo+yO9g3GsNCEroItga0BeA4jZ9icN
8LSX+2aE0D3q/HjJ2UypnqMEOv8f5Y413qKKYT7kjHTh4Hz9XxmQxBG9PRLi3r41
rOq683qAKyiJp/SHndeL9jSHOf9T0fMoz9VRpGT7RA3WugbRC3GlS/kIoqQM6k0N
/sops0GeP+LoL/yB4Ms7qHKH3mFtBLqXXYe7umRp6+VAOSbBzoUj0oZCe8EiH7Jv
LOlynZXQB6ymWN0d99XiRni1yuFGp2QVFVzDNusij1ssURPmCbw3f4SS5PrlWESe
V4Z+mBIts9xUMKmjYMOBaK7KQT8AgUCwAaZUt8db3GF98HtxZMcB4JB7ihZrNIbL
cLeiI7C7wEXdJQTSols6J2jxpexsSxNDGBM6Hv40W+cHqcqdd68SlbYmN3al5TGJ
qDYUBTAcuC/mLCjZyfmOy1p1G/G4raiTHaYWRzBVCl9RVruar8q83tDRAd/x4Ho+
H8pCfPLkT1WnvCW4RN9+uogqGEeOOrc1fuUfMXsFJSQ3zC1amQUB2SEo8E6hWOxw
z0i6neabfKPe7fO0I+80ba6PNC2G/x8Ezb9qj2MfN2ln8Dy8d7CB86Jffly/ltvE
L8itaUrlpm2ru0CB2OGNwepw07nsO9UkRkAQRK0VNQEZ0JQXtjr6xGCZiiNO9AtE
9emGq7kMUsutmKIvPX0vHIi7pTe5QBUOSTREvjh97WZA62rhVHA1rEPhVQuKkipZ
ks7spgp7vGxtlkshUjvsLAyqjqhPVEcJLKFuVuCgOQRzkpu1tR6Vx5GKIXeY+wHd
zYk8rfuNx07sTzx5pg7jX0xRTomQ3vh8ER5kHPCNcjdIRMGmEejIsVmFR+BcRgMV
F7ExX237FsLWQRbjmH+CUUsX4kIUkJGX96cQpMajntf+4n0ZxGsDHKKgYOlmL7BS
VQs7k9cOZXAnpKAZAfv3Ck/M9ZOqRk4q4fk4w7y/HQEtor19RFcPqReHNCeZGIq3
3JyUpc0bcdiVJ3vJy/POFQDTqI6HKo6JJz/dq4hEg2y+g6E99VUu0IZPa5zpTUgT
ZQsf2Ah9XQgRYvaFJpitUDOIeJRvBkgVXecVfUUan/9Ec8s7RHwOfjHzJppQBzf9
EM+YR5w3e3Ldb8KslaK8k/Kjn7ptF+VpXh8xgxFOge7nce2/W5PmjJhr6ncZNRF1
7nqGUiO15rUpQAEcIifLkWEmpS3w0NLOBqYTt5kJeCdMOtHYqfro41L9K7WF2QaC
DINZ/iontWp9uS4Tn0CXuExAIAqYnysYpf3nnpld5zom4FKzE1XomoGg9sZgILr+
AWXC0YIeBJvY2NI/s02yWRgQnOspGu65oOTjlW+r012D3un6DliCVBDGproLb6bO
dkPahBArKqwV7hv11GOlDrquZGYTM79+e2fB4xmC9faOw1G6Cy74/DDWLy/moJLS
DyIK2NazkX1bWbmTqWIyP4NPsoTeLaBO6+q7sYMzSpwHVh4jWwHkszTK078phX/r
hrSYgZF/CfhvipDzjwTDpJIXdU7HV3snUlZMCSXOcaS/NKQU6JAytEM/XjRH1Ssc
OulwrgevNx7iaw10CBeHN3MlGVZX1T7j6y+Wno/LyNpHh49kLfYdDMjZGjPQwzrC
Dwclpq8pQNqlVj65RweHTyNRVoNM1MKCrvK6dAQi2pgnmAj99tjE3YaMWfDcRtA4
SbMqfGCkv2QrE9Ubx6Bs/cCxUy4D42ts3a3jLWpHlBfsboYZ6SmxE9+fGaTSFaPl
qCNFLWqvVq1kJcd0pD7sDeDJgfTAiNN69yXzZ79QdMnMhHXVORESEizKHsxoNaAt
heayqqQInIx9JxGdDJnKi//k5us55Iy6XoGyIdCcbHXkyPHzBhFIDbL+uZVQBOhn
cVjohZDkNGu6QlC8xfcS61Cla7rVXQM+mlNsufjIsNGOW+nY5kF+szKIpXshpqvz
COxxSmj+lD9gMC3dfa+6ZKl/6nqaPk1jpYJ8i73MJQ+H1cEUkut4JBN9E2r4cBBU
D1PyzuvplAVthFYhGDbhYMYkr4LiHvG5dT589vs/EYwFWGVxbPUDUD5gornxF1xD
RhK0bzBeGT52ITm+gXCeTgkEUbBJ8TgxcI9qZU+LfrzZt3ZsCvRmSqSBRvnedwvZ
ijXkgcDumqIa3iWVtzF5Vyf5NqYHGSqRuATxDol/wUkxccBLyojtQqWjQaVe1Q2Y
yrcc/b6D3iAbhGr8ATJr8lq6cb1lPe96Na1K1xnfCKQi/WLRTPbND6VW0Wu7S//5
QUyXM6vMvTdtad2iUPtTccAAFQ1lk8pIaeCNcYqS+wEqJoDfdAiBsgIvJhtjkUwh
BNoqGbGO3H5G4mLjZqU8Ho/10QXgpkLbEmwil4b0cmw2C0VfYpY3p3Go8yKZRt5Y
wTLOIrxnmYVLC46vSeO7xg==
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:33 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N6Bj3ikNOXs1BfxeMvg/7mia+EqTYnalNJ5mwDouXwEZKcMFJjo2oeoOMIogp1SJ
+x3ibvohchRNPYZx5xuAGlSwDm08PPY6EAsuwwc4l4uf7ItEVfGG3ZWdH5Ul0GjE
yqgI+nwICdImKCM8AV78QdiHJQsjPQZ/cdckaXUss0Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
pqn7eeB2QwR4KpbD7uGsJUfYwOuO2UUoyddXp4/76wMFmufDE4aPAQ8xTYrQZ0ZD
Xz6OeceSfgBiEJZ4MPBc5mTk9uupX3QRwJ+RivRoGzDB4qT7R+Nd8slNw2kibt/d
fsXWCsonFQeLykbkIL8ig6uonSKR8FRTGkkdehYH8oxkrGeN+VN0QlfydR+QjxPQ
oJ3N7/PiadtC3A5WnvykSBbNMxpTaBiFVwsnbl2TLHQwbny28hfjY2JaryCAZIPU
ekdywFEjzzoFc3ShKM3YaZQnQi7oIrs6m2vJlTyJ3YLXM6CPi3gd371WW6b5nCBz
8z/SK3pkySETrH3PwI6sEY2Exo4SQn18eX46BG8GYX9OZEmepwOeBsjGkkpdhSXu
cQhfl6j96Byv/deBIbc34ghjEqwlcSWUQKbQICbTmzD5EDZOwJMX62WcAd/SYpj6
sMGKQNbPu5y+WVnRrn1pBFEHXvmav6Mn0aQ0XfauDYQgHb/ENLtAnrWBYey0YZiM
K3LtnXnocmTzHq/99F2daWqJSaHScaeb2Sg5ow4akfhYyusm3zA8xBME5Ltvxt7u
cZk9PDiGyQBvWRtHJYyUChKU3wF39pZl5WgCoKD7xKKVeZs3iMgIDXZN0x8dBZmQ
1Y0r/AzgnkxOAuKKBRNjfqaB0ebyxmq/PyGS6HeptLvZGkG6TNI+slw+bt+xvH1C
whRVTHYEeDTKBFFIJsux3pQbsq4QVBFDl3O/yO8x570MCFDM/nIRBIOBLoFZC+Jw
XECUMjYLYc0AkSNxb7SzvUVHGkONN4hKCvqTGvfDPZ1GZgC1hUkzoG1jdVNQpAIi
pY2Cq5Lvp8m2BxGVbu4SXCnClMoui0P8LhEZ2JZMNjFTnV8WtU5IjrsVhqT4ExCq
BmX0Lor67vAvGAUAKeG+DiO9BQNqwYyYVyvl9IFj2w6w6cN5YsfwZ/WgS9wywPuX
dc9cO5T0dRghb/Zylwhi22BfOdZeq+PqP5m3yA+R6JlNHJIPOFtWd+jHb3JpmpM3
O1GO5V+0GpK/X7GhoKxYIctGSEicUy68Nv5q8exmxSg8NT9iGd8YtE1PuxqMxTLh
AExFkf2vO6ktJ4uNYuaDaddO7sYryUDw/n2nEC4nd+tKUW958FFH9xXGazhzFF5p
3uhk3qo+dqt4nn3sM1kW2Lwnx2IrzoKeDsHygNPJc+jZQfMMS5xO0EsGKFRdSfET
ae9u46C23Iyl2hucuw4bdXzN1WXgw5Z/8uEBTZRtTcSxosA6qwI83lnwwlZAKqBn
JwDOZdcaBsw6qn/mevLZIQZPOCNoPYooUoV36YQv3tO/FxoLbjFLalOA9tqbeqEo
1rcsz/ylB9NYb2ArhpNIw0WL/VhUuImJAtN6eilg7Rf5Nnsa00PRTZ2D6wYd8llK
9uJblu4H/r7fyFD5hG4LLBfKuEHPkAoXfspZMRDzHyGpyn3vfBkdWzg0A4nCTDNB
FyMAl31UhlH+yowNvYAUFrgKH6dwwXrPgq+yYNy+lAgF8WOVAhmdiezL400MJQ0u
myQrEpxIi1jOkoqEJ8fxHLmwh+APxe2LtBmuq+d86fD1Fqo2FyXSNf89YGEXQjDP
vSxKdELvcN966kRJz1RvsinYvipP1XvZ3R9qQ+QD7l+lwJ3HgI+6VIDHKiI58JSu
gMoWZIWi0DlBBkr5I8++Eg3TD49clHKYI3JdLbou3v8iqhbmKa1VfC3DARxOV57P
QzvK0/NjzEeHHN73XMRPoQR+i9WjQo1zunWsvWFPYWqbuQ4WboYSQcpQuohpyTgF
PzGVpNMqdMrA1bDC/tFaYpTSgS+nEB8aMG7IgmhIlL10RTVLEzuVEOFzF+5iBtBU
zME6uS6c05ETygt7q/4twQ+RJOVXTaN/LNvQjWR1zG1v0FYPdAIpslxqO+MMuUs8
9ir9jz3F4Dq9lHvvqzMTECD5loZFo3v5eA6YsGXBt1hSmoNgBSmAb5HckRvNB2gT
KpCvsWlId7Ixu2Kf1Qc+9cUESWdpD510+XBPA8HXyRwE0T0BUjRl7Z0+imdhh7eD
B8H62pH9yH44InqvJDRo6aEwDAcWXnL8DV3Mgvvv3M/Ge0Drc3bavS2ABxyTyxRn
9o2sjrZ/Ig5hbRwss1nZZAY1pkmpHJ2YrRMpMLwBowkFTJRDl/7/T7oud3cc7u4g
NwOp56nsrWwEaAJV/zhXY8PLN1GxXIywLkR+spx4zUFuH2rrc9L3XxYfos+DDqxa
0BdqKwUcQknt7fuOpGiqqwaGYWr4DeP2ZIXI7mZsDXcp8JwIJYBojtOwIE/bftkO
l1SgMfHB4beMqbPChBvtkYA6yTQwVM92AY3EgnXGnrTR9QeoKR+PkLjohRvEZlc3
wwqZ1O2eW17n5TgQUw5nPa5LOZuzrIjbdAnwx+hra2hFd6UotFCHja1sEE2Bb5ZB
P/XJZSmz2vCEVpsGUza98fAjTBgprtPebmGE9qn3ToFzXdnjYBDjkqiJ9vWAyIMJ
3oJR1nAm/xnnU015cU1RBoRY+MUqgU4IvvwiPgL+kLbk3ppXmceT7z4UI46Ok8u4
ptaXXyipf/bNhfjArPBNM19AbaA9Aq7XkqaUwktLouUolz2usQpfYftGHn20cE4F
KA+Ebik89hC5GR7yK95Ts5uPJrT/OGsTiiUD6aXsbBkB7PC83315Ou9TBle/YCkR
rBpHbQ2JNHQd/+fiv3tUJwI/Lt3nffMztOLURWXdSB4jVx4wYqWqZ98PxvDIPhjS
opHEB1nMNiJfPFmrmgHC145Cm2Gm35CvLp7sfixaZdfXLhp7o96ekD7rJda38AOn
IM0ez//ADASqDV+/j0Bd74EjhAgKFWWwZrF+FWSr1c0Klm8VTtpYv6BhaM6mUptj
C3fwel/q/4WpzwT+GPJH5GThoDXsCi8sKA+Zk7MbC+xcxY9Bbe/bRThaN8XHe3b+
xxjsAnFiq6CJM0OIe2Kp5/iBN0iuoC9KICkPlELg+MahkXZBbo+6qqCAb951lH7u
6DdvTI2E0RGqNCecGlj+wSd+6ddyiqAKvROio3ng9ZErnAidCSAPAtJDXK08+lq6
pNmXQdxxoT0Nkj1puyDyyQ/mJLup3220oWxqemtDbEPSlsWxawIjSZdxY1EhLRs/
iVCOMlyQTKfGFleDf5H7Vk65FeS3i0qHcwmPS6Yw9fd6O9ViR93csZKcvBH5bc2i
FmYRU0txxIb9pVMcrmFVDQUH03SYhNJbl9ra1uZH0wVU79QswSy07DFcqhe+Ydhv
SVFkr3WhVCuMuyxETrTbt/EDOGStfd9qYhkVOJudAF8wHBT0ogB4Tf9EWChcKYVV
PUaPB0IGBpXN+PAYVk0MpMKMJR5WoPIa8Bca+3dpt3Re0XGkSHZCL/oRgMPLVPw0
P0MD2MyUsmT8wHgW7PS+FNgocr59afVE/6+TkffUbMO+FJLqhntSbNqfbtcBtZ2Y
Pb3B1Y0PHNeDDYcsHSDH3v97QjU7gKrg0zmzKCi28mBipXxTXHU80eIcpgFkNbO4
E7z0xvoi3HpnA111OaGMXRwdatmrsRSa/xMWTfzi1uMOHXULXjg/iwqVJsAPLzqf
FXVdZmLN1lLZNPe0JeV9GDhW/p8NcbqQzTY603FH1a1N6KD+fgH12ShtYrTJh3Nr
YDoqNcimM0ltdVK7YMYAkdAzzvUCanwT/Ei8KMavWcPXtIbdLfIrslhUAi7xn7FI
XKoTR+ROmtmpYDqNhuaIpbO157Qtjhqlr0i7mO0/8j7pil4aBXALFBJmgF987way
dvR989VtcZbJPPHGgZMWNGP4iFNJVmO5brEZ/pbXCSihiD12LczXYYljQw99elpw
h4QPUW/Ft8E46T0oDEfm4pLoV6pwSSVEAEyQOSNR4mESkrsiz0cT0UZcMDnWI8yU
LgopprxPB2996+7rkwzILcqa0RdHfFc9DEpeWnpkZXChjQGRmW/Jy8vG2WfwRdC3
WDzH0lum7qjOTuliwsoFw6fipWHuM8Qcf6t3kELsegbOz2GP9osTibyYD0Q+DK4j
8rVcKWB+7KIodCH9YRQNSOsLTdiYJ8o8xI0dzTE3txiQCtEqar1afl6VPoUyHaV+
zkevS5/s8njr7NztIsY64qxK4XItu/iMyoifcPdpHq7ez3ak1zRb1IWa+HLvPsSv
UwyV+ACs1wFplc5UJyvOshy3tVmpsM70mv+r+PJW7A4aqRxdOZJ8f0Md5+UOSw1E
KHQWdEL80DWBUSNrZRUHdj/q32Pt4NhCAQOaFGBHAwux5hUd2GVGPhMETZeMaocC
MPlAkADqvVU5409oiK1ildfQIOofdpeIXrXi2Cwx9zetTW4jFCXaANB41PU31SnO
/Vq3VFSBM+5xcgGChGhY57/JnyYsH2CdNDf9qAOrKtEu8TdEOh+a9Ip0TJrtRvOe
Ou/+22uIZock4xTP36rSQHQJKMVXfDZQDlIkqD87deiIA6iP02dfVzdA+1ZjudSB
T4fdpwcNznNXiZNtiy9kPgL4Dl7ALt7gOdh5Nkhy6i8b5oZzoI5l8zSENGWXZou3
ugwNKKjayREhDM2LjQyHcwHCPbLt9KROk0Dwm0cIvPIX8e8ozCC1mptvy8s5CULq
Dy4t5pqnjniJygYv++mcFNfaTfiVzekl8LgtM2kbNGMumFrcnxka/KHF9unmIO0L
88r1bs9r1+AebVYYFeMeOjfLKR5kkixuctLDs8L4XVLwZO0rp9bbGXQUlwzRzNgu
K3qe09I5Mgaw2lt96OENOz1vI/MnXMogaVoAuPjpB7oVMoHr56Lv5TzMFeUfyigT
LhPCIt7iSzPhpnSPQBCQJbY9YQskwHZviv+4jT365qfOu3iKwDJ+63VM3IC/ywec
o3fyxMzpjrTy9dXlVF5HVvYeR31aTQFicsVvM7hRoacEPcHm1DVom6zz9iJM0j+v
/GGroJZXweYECBuf4jrYPu2kM2JlSPUwX7hoOhg4dJ6fF3sp7SpPU4FskNuwTwe1
BPq1MxtvsxKtfoKp85gEFkgKPRbgbT2q3rPsyvcjK+D9IxVH9s9V9EHRul4V/uBq
dPeKF2iRZwSZQ5Gt8VB7o7vYPqTZlCbHMetfVzo9PdC8WwApX4Bjewk2093qiFXW
4bME8eaq6h8uoikaXKJ5lIPMTYVWOxhbv+S2IdV2w6hxKuo4JAOFR4tOcQBD+0tl
VtWVCtF2tk5ddTsllPiBskznB+vdc3vYV7R/a0/ROQQ2NL7p2OLk7S3+trDfnyhS
lF9Ppnk1PpRDPPT6WzXfSskwA1kKWs1oTQhfTl0i884oKCHwo66x+15Xq/Lhtb1D
fk+NhgmR3cDMgkNSiGa0+8zNMj/mEVYCgHzYeuzFR329phdE+Rpcxa6zqNQ2YiGS
5dubJI5jF1P39GIUkR8udhNMXB6hkZTGMjL3DrwxSksl06R14qIKl/raWF3K6cHs
G9MoqzAja4H+TDaF7JyR/pwrrddojt/cUV+CdJom+LzNEIdWswWugVzg+MoNXxHC
jT9ReeUtzIFbdgaMBltpBIw8aTo1c3t+wNW9mpP7LN1drzmhMwmhB0Z+rFY+PaRb
Pf/x0GmKYrdCOe+cCYgQTwgxmts6vt8NJQl60aZhYuqoHwadAVMb/I2+u9K4wqVI
oMaW6ErS2BIO7ySSiaj/NNO5uetVhzW5wPUiXrNq2UJAW0wRE9rTXsqM3ksEyU1h
usYd9A7Ps2Vh4MOJ913Om1ZsC72LBMSjNiWMk2j3zs5R37GAn08ePpj0VDI5eKhC
91ChrJSlGcaI7gZZTZA0cuXDKrQjsKx3MoZFc8uCvzy9QajRnQCpCWHY3+czuLXj
FIKjlCV3HEGjk/3viD4OAR4HMJGYQW4QxNPKEePxlcN+p6SUGZwlu3drC0PgUwS1
LSDypFhFAvfko82xSNKNuJL7czDj83HUPXgPYHw6R21t+tQbB/FrDuhUUM5j0Nq6
Ov1PWSQOiEFEVu7mLMO2SpMSSn0Rc2pFyhFUNmNhkmh9PT52CTjrykkj7l+NNUJ1
Yz6TNql+AEEKp6Azrr5TbRdcHX5pPmZpuUeNpbvC5UNnUEb552bWLV0r4QT4xcHr
Cy9Q1SAMQ+WW5GNGubNhNbfSf5qxbP3soixkzAxQm/YIcQvSw8XfDWPNyXeroYpD
81dHTAprkmpC1rxDAZ70tduekaUn/QM+9Nv4qRWiiX3aYzLPV1yIbZ1Jn034r1vn
PVzVPzUkqcxS0SELb4hyiWxX6+Cxux2xHTXwvqwhPxLSmzVWXeXCWfnIL6cNM9tA
bGpa1GNZbfzUNxc70rJpkwHkV4PTNjLBvAFnGW95r/5zA7WTAbM5TZFVBPifDRFk
cgV8osq6k5IWEQQgdW4mgXWfbUQyhPRHSYOCMPRIJUTfPDU/jIjRqdabdAtrVAGy
tCsFtle8rhJRlf2emZphdMjin43R9i034JIU3tIfKsKU0nh5os6+3utcgBVUMT7A
zNBeGApicLkt+xdRPVSOPYLYeZo9Ni9SbY/+Rfv7ZhT9yJ2yo0xh2WxacQ9L9HUy
7Xya2QEr2D6b1gsEmSytvlzVSiAcFu7L8a1IT8fFnkKCo012FRhIRglYevdoSCGU
4nFGk28DPytngMXA6FyAF1m9f35XU39l1Xp70B6XaWMZMg+m78T0NIP/cepykmJa
4rkQI8x/kBr51IiAUitULrMQGY+zHmkSL4MACc405zwNFRPBvVdkCN+WayJ6Jke0
ZSKdrL+G25XJVz9YcVfF2czfuWJzt1ns/5gJt7zLkNTvBZgXD0nZd9usZ/Ybjjil
jaQshDnlSXuGzhK76TD9vCSPDuzjF23ZpmVhorLk82taeZK2RiZwOsE9yWD/yc9+
kpR43htkWnU7JQRMvJ9U2c/gW6fq9wQbDdWSNXMx/tXI0jco1Re/tnNBkSSTpsiE
5tESbNUjbKArl2dr7K5nDEEq6gZLOmXSCYMHACspsh4AJ0nc8xjZr16+hIIEdb6D
QE/fwypSUazYy3kJwRsqf0isx9dye4Mf+hfy4q2V89fKo0LDb742RPuuvesdve/N
9nn4+I39aHI+0wivGR3vljDdeBlLTFXlzBhMiQl3cnhGoWjqet5RyGib/FXZ0c/Y
NW90InxSUIvF7ANcuXUTIkhlCjTXctV7IMJCKoBB2qXfU6Nb8qtxXSLMO+i7wCdR
DcvTiLC9fXvYvImtHmuq5Ik4Grcfm+wWS+6bVcfdydtNdFl465K6taR6LATPbX48
qJFMSu0N9J/FcK2LCxzOqVHXPQaL+4ZVTAtCCgBpL8kpnwyhgDRtmDAJ8ArMGNc7
FViTOO6J4TlJ1CgGJVwEaP/9JGdT+H5Jxc+Np7TiwBfS6fekNkvuWllD6BKk+Ooh
eeT4tAp5LzXWml8In6JOs3eLVEHrpMrX3+wHgkMx/ErDTJkTBL8BUw+i3lbx1goM
cEkR4xJRP1duOif3j1EHGSXBxHRsq75OEcA15LTT0q+wFIG9bQQ5kkXOoag+9Ylu
lEGLYjukiynCGCxRnn7leSNhhHe00X7wj+ETayL7HPgvWuc72+b+9AuhW5AAvdAM
`pragma protect end_protected

// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
nV6FNU4SK485GrzdRUA1xchswzVqAcDh84BSzdoPmPohy3vbHK37pxz/7GLCXpLlPXB1ifPQY+6F
Fq/tPwe9a8umf2oqz8ygbqreMlgeCXL3vraBCNADilIbr83BPE22lu3qLFJ+ClhJz6g8/smSkyVv
14HNI43In0P33//7o/z51BzxPY1M/cQn1zFZwwL/ydKN2sYhLio0NNykIjtI5dPUPfzc52zwCXjt
cbtK+3j9eAcpMkONh4l+ExxDCKtk7ZSEu1rWGGvCEymFJ2v5RQPjvQJgdrdzRWjCffWFXKSH4NQi
CX1chB0mHSVuBeRcG2qdxnp7vQUNS5TKHzyZ2w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
UaGl7vObFxyhdwWQt5X42wCwYYxvaNLEDRCq5Xp7MQjPJLoVsMHTKrykLEuZcaZeiQAQ1+4np1jZ
pFULIGOnPDnAuD5pOGLASKBZotZ6tzmHpZtQl3vQpsoAtdEcH1a/7C1AnupeLhZxTuBaxQmfvYLo
sen9Uj8IFD369VGZplI9MoDm8EuX6TNFItTtfAGCf9lE4MkK2UnD6VpptJqTiVOvjtfhvYoKB8Q9
lEakLg6Cjbs3NOpuNANmfk7zgmkCDxsfLVejMH+hN/3OJVohAMua+ACjjNQDP/vgY5bFoWb6654L
9jaEmKrJNYKFBaGx/UwpWSLbet+MI+FSiMg6uJ+iRGZeHE76h4egp0Qs7MnrwltZwGwfnHZ8Rg6q
04fub7S67GL00kKBgmECuD5VW0BcXrVD1/WA3+bt2KwSPm9o/lcm9cr2RJNE61qQFpqFBROTmDMe
8TMmEU82OJkdMeht6SLBInlVcjcC8S9HCNp7E5w6QjIwhCbCO3Z8A0+iBe9stqXWOCAIwYKq2TPy
tkxzoZsX9nIxIrjd3/OXJePKWvanTOdD7VhV7tfSc8ONA5rC+QEp6WFor+MkE7DdJc5lLDo4ttIU
qz0jL5pl6hLFSeOifK7IvD82L8WI307XUMhTU7vyrby1aLmwG+C0Uc2DCaDKy0JjKRCCXwgHs6X6
67wWhD/6+pAzB7YtVpfsKqz5El2Odo0QJd7TFpDLgQyBKz2Ms3wf2SNDy2NkGKBO6emBayjUR8h3
oWmHr5KZLk0PHEzGEefe+DFsyhTAj7NHr5xFVk4T6F8wgjS+NdQbRc7LfhQzvgGfEbkOeyCYhlvD
9VTbqwQf+OwfH+frcFYM+wMo9MnssmeimKkBAnoOlaLGZoQxnKdtQlTMstCyn371YHtBsHdv2Vqn
5GksRSL1g1nuxyM+bYPzZXWS035g5zefM9+HNtY35oafE3aRnDR1mJrk29t08NUz1kRuNaEfK3ZL
P5VsLchgmD7dbWhYusKX5AjbVmiR8W7tfq7xIdQ14MmcoZJ4DSdeS/P6JWuHSuqI8v/jvEKrH3xB
rBjZMKm2+w26WRI3dpy+KgcRUoILbBHkDMZt/Cpa05VHiinmyfKFCbkWQkbZzyEhj/0TdyThoons
yUXdzd2Ka46AsaRX/jcOz/4Ndr8NRBkrrFs6r+XNOwfqoCQ6aTO9EMmINgg06anvMi+pOdqE7xgW
8ZfgyMQkx+I27QoXlMV+0Tr8P7VxHbYuVSzq/6jtEgODhekvC5J0NAkj/9isykgglIUyPvJMN32R
ErRwjHOwwAFKm6b1Q4sFEDVFayXrASLDpwWNpxT+hGJWi/KRMeMXna18Yn/sidSodeYkn9NYoH6t
9sINy7x1YwPpUEiAPazJ6SXImSRNKfy745tyYBPyp5IeNjVIPGbmhXqoCxcrH/f/sdHAyOZx2iGI
vjDZv9zEfCMRsHz8kmjdhX0jlQ1pYYpnMVFp5td12GB7ulWDXIYdvnmFxKoCqlLRP8ndRCr8zUss
qlUU/p5wKAgZmIMY+maC728ea3Pl5Z0+dWCERuKoTV3DS3yDJXzH21jGWaLcoZJcbMWN1tBYee1V
ndQ7QxI9/n4/kkzsIy8KCdoyE/8KVZRcyqnrsrdzlekOckrmWCMoYY3PvyXYcQuaJsjeZScVnzyl
sdWRcG+pRHcmXwk0yHD78XiFbSi+ytNGCFHOFMZep7QQH7jMSns4kHx7cmOg6ZJHy35qLzAcqfBY
b3krEzFtT0Yp/mqhg5W1u/FdVTFV21T2EGNrJj0wGuwlE+qjAUQX4MxAl3zsRiRexwa5P5wN3lar
E4xOTKqQfSGVd5t4FGB3MTE/tPNbSDUpwBOWw1sv1FPQDxLe2jH95aM0nS/ka9qWAcnpV2N8CFQV
OX4veXnOiEbD/74g6Qe5N00bstnThiKABDRwFn1F4fzRFMK/+b6M6XZnLL/LFcRQuMxuxarczNT6
4durFZgRwMhx4qPEZyOGPcQ1Co/cuqaYsqBPly/lRbQWv0e+8ZhONL9Lj9TgbCKR0Tt3YpzVrvec
orgZIb1hFVU/0p8CaXUIVDA35tlwCWGahzYl03DNAE/JoReCrEgqBpInke3TE6Er+auc6JQDuDk7
FDyySYvZows9jPjoAwHeXwTxQbBO9jTLcKzEccwm/xGVqEZZ4vIkhGkLSGu4cQ2lKj4L+fTpN0aV
fvC00+WAIW4WXEPdN2ORabWwVyaHZGJ3ypMIgWCiqGLlpm/80G2r/xCVhwsd8cPiVAowJOO7Ho09
5BIEMHe4Vita3PoFDdXaJfeKBnK7kq3KKN0DNyi+hlkE+wza9XJPyF7OZP+Hfj7GoZoF9GY8A1rz
ms5aRnIgs0q5OjnThQY9TkHsLnjid4HI3NZW5m+DoJ8DPGzZ3ZySAH0LNMvTM+p5IHzaFKG+cHvZ
2ykKa7GZfHNfRWWsK3LqNTxHvM5L5ZOdHEXp+a+Ql9l7enTSfWoREn9yGigOhBualVRlu77C4EWB
k2w/Bacfs3zfGa6HmKYkfZ5Gp/PlVfkiTOVyHvvO8TpyefAJPWPf3KBELymY9jFbKgSXtIg+WOgc
e/iMn84DCAmRU1Qk7z7dmMTFwv5sz2D33cxg6rbUkhUGa259ybbzfwTMMoPUX8QDa8nFztJEHs/y
usUbSWhTVhL0r6PfKFBtl7fwvHvl3a3eOzaKrKoCe7CBmfUCWzRUb1MavkG/4QMINhIqycQP6gGt
UQNuHdMQMtvsxWxIhsnWgzZYqTBzMOsVD91X8wwwiS9DK4fBmJpZFxhNzAdPYC8ALjG1oHn59iR6
BDOr5lFO51zxex1C5VnXqTJO5NKEMT44RwQ5vrVPaNN3VEPPQjwdHfmaUHu26jQXE98ibIiyjPx1
4zXNrrEvET8brFteIH2iBCifJt5/Q17torA+nRVR8wZGe6n++zYgUOT+2qkVtxbCpufg1Y7n7jrX
khTIr7HrQA3t8yz/8CLiPeJO3F5NY2jTzLltdneBxTm8Jam3ROu5glC4Fpp8Kmj1vjDRSjHu9sXM
MXVuk+f2bV9ge2NbOI7l5McMAbcuMtUtYVh0uoMjNBtvrjGC6JIMo8mFHw109kdf/01e4La98u4X
tkybmrBkohNzzyQLu5Fs360BaI0cwLoAdh5H5nLlV+zKHMmj0MI3LWfWJdmqlNo4m6oR16EZSKEz
z7n1I/nVd+ldbRhO6S2ZyTf0YefUT8e/bbLcsIlwKzm1wHdV8bYW3URiSyjCz3kvokjPslh/jhJu
n05YjuSWhPkPRQKj+F7yrR2Upt9Cd0KfD+PJHMtz9IhTYtvbbMoCjRwpics1vBJKE9V4Zy565ju9
/SpiFi0L6KEyaLY+evhNfLqmm24vyVZWStjoccCNwXnQw/mU1LD6bxldnLSSnK0VirWSPFwQBz6V
r2h5qmMYWqJaL8ELvojBRYOrB1RJmsf43JEUci90LzW3ehg0NvYfUJovEkQ9Hy3d4MgOrGa1Z8ek
L+5OkN3LJYQ6UxYU5tbjpsCjy07WX0lNEg01/Jg/QRUcu6LHHqzN+w0Z6phTRNlz5IMh4pU+2sMl
l1lYDZPuulW5x6z0VVK2NqGicC4Y9C8Jv4xw/hsLpBhuIzz/C4C8XsH1V5pdyr9yeLjtFkCdJijQ
NZqTeWzl7WKNufcDA8XBtO7luG3ffmXOrSYMk3xBIEYO8hUvSUCn9LgFLpjUiIBtahrrF9zBwO3g
v6aHVF7ZYrpOPX5RHKAuAeci8A6Kf2oxYiGESZaC5zQ/ymRQXgkvXQmCuM2bY1+SSi89aFdIJ/Zx
yLrwJea0qkMj70zAMgku7QVYepQFvKbQTpq9zccV5pvSqwb4zI9zzzIYDwNhd4WObUob8DoVEYPG
eVgoTGiE2xIsJE0+wblDQjbxzNf3GC3d44H88ZfC8auTQX3tM8rh6Ci6SeZBxrrD+SAfFNckN0BW
Jzi1tscrpsz/Z/5Lo2AH12Su75xom/oVacJr50xS/Bnx+HYvGUYkJOWak8eUSH0PgnCYfuYGR5ey
pHBLrvY72nifLeTsYGLZFThuSn/mrZk0TDX5TYravEno/RM8Cm+QC2O0dAKD3GIdUTjAauBW8OFj
3DVgvJXrs7mnVb0BX7rPXwBhLtQK4GOVh0HAvDF9kxgz7AXyw/Opegd+qsjHveo7pjrAAphUS6XP
ZY429sqUIlzC7wnZuSVANmQztfTSfyiFGZhszvgnm2z+behZp2eiZxOkO1OkKSejOfio5dZmxLgr
Q42mb+OUq0H6k95CTwHdOyTa8AG9VoTfQTYtZUy8ZtFuKPnEGsiKnztAkqFIPFyMx4oILJuWKOyf
3Hn2yCbCgYZ7PTCAIltecg+jB3G5SiVhVze6K5+4sUj6BEb/osS/zcZoDv2vJh36PD+sUdvy54CU
LzdDhqa4nesLWwRPjRfadJGie7ZeZ2na22PvIbrQY2NC58rfNQITYs8YuiyjjzJqvZaNLvUnKDFB
gYKZhYs7xgtRqadJHntq4s3fRqpPHUwwMEG5Uge90DuvGE8ChcuLzLJA7Hn0QaFKmxEnqI1B2vkQ
+WcDyhS2fojn9Bx82gTTjQXOx5a7JKkFIJ3+U/gVhp/bFoaZ7DIrlKmQ7K/cJXYEvtq0uA/40rwe
q8hEr0eSgLgNbc6/QBUlILi3mJvh+fIr7QHBJn+PJPNWUEsHT8nLboF5xMSayD2jB6BmWJuaKeSn
hS8TU4OUz9RlJACpyxZ/vCXRQJY7MDH9GAPel9ZpQGApwdphIWq0b48c47fcuKzrR7oQ6JUKGjP9
Ei9typpesJ/UVx7vx6idNc4dgnb4dZaJofoRvEEE7sy4T+RP722gIDHNZui6zjExQ0MfFema236D
bBzaty4vOfIE0+2DPy+rUmvjXd6CQ6FmQsCJE81s/RsdbzSVcnE5bSN8FxGvK0EiyQMTHGzdbclT
ovCZrMU1e1zZxy3OutRU5WclvGHaOE1mg/r7LR7xK/cExtztS7ja9KlZcaCsxyEpqJqEs1SOTcbf
yKHjpDOz/v6QpprnuIIilPrw3YCtDJgZoYBbzkmmd0JmFBxmwZHwPv2a2Asgxjhuq31q4HXZ7t7Q
npDIOIpQQ9NnMXbbMdeIk+58gG6+U1C4UoqcFczHhtAewQiSf2XVH+XKLyfSqy/D/cV5yLU9I4U7
bhcFwYE63wry1plszTaocYa6UKAQvoxAbieiAOQYz7Aq9GH/xMuYsHNo1OVXjxg3pLHfCj7MYAWp
ZmcWbE1ZOfAzDZP/N2uXRaI2Illi8CFlXH+5x66wyYYpLjVcWbRULO3BOQMTkeLlcIwdWCw2gUgx
xibYfjJzN4slqBMgMFsFaeeQD9HJbaijiiYotXgRerX7HjIReNtevM3sRD5Srii/cmhDqoReKWud
IRnFlXOurtGBM/72iAhRJmykLQEKfAfn3miVrl7HS+dyQeXRe8LxU8wPZDAl9tdMMRb+0cLmmaJi
7GE1vVqcxUnhsqpepl9BHtKhGuZ4BlU3BdPiRl4kWQLTsx2GJanoJZ+Cr4x8tLhNUcNhm/HAPbfr
x9GAo5EMPWg2VOA1lXPRDjyYiyl+6T2rC3DFaOqpoSX/HWv3VbiLm1dRt7yG3ACXrSqBmMVkHdGG
0GpXhLpLkCumS1m962mPC8VcktpcVC2kBdx50Nsk7Grw9T07qL7yNY36I60dnGeldl2UnYaJRwiB
uHl/G2Sop0yRaKHvPakEqDu0yg5omAs5QDVazqV2XiAXVp3kw/gPjrII9eoZEUbFKWRDJE53rJ9Y
ELiivVsafvZYV3gOQCrx4wxAWWkX1UUwyTQef+3/8fXDzsG83+Bn3qHwaW4oGkJ+qg2kCoMaKtPF
g+pz5WbTzVSYswJ8zRxpA03XiuXdR/V7KiW1JSx6KNMLllHH+BUO2uYGTdsOFkMvtzhT/zgUXfdJ
I13ulKFDGG5nw5dyuqyRpuCW6vk/ERnvKBXu9R3Adre5isoPWm7xUzoZYf131Y7Dc67WB/SRx+yr
n3u4OQ9YWXlUMkKdRQCCxszi813GTp9aZQ3CntQ3knJUx3GqiCt5HJM6jwBwfL+DgTHdA7J2NZTA
b91VkY0IXXcQ++ujeeySRGQIGJ0M/BmJt4St5Svu+N9dXUAkU4RMEnZxOifFSSrM++Ce+6eWq55F
Sp6+B5mO1VUqJvhnomsmHNqu1LF00/y91IoRBC1cIyW9pxYQy1or+IZLJqBD3pQBVORatbfArAtk
C/uLssDS9/uHxN6y2cIMcdetM6Q1Vg/qN87JHoU15pi5vw8Y3dbYeWxhXO3pHM4P/B8sDLzXvIgc
0BLga1SnflIjot7X53iI7LnCnG4mCuqY9n8xvqxvEDc8orwaa0PPkU3q6jZPVOM6luMuMnf7p+VP
Rg1PJvFxnirbUM1DV9iq1SuUQdfgmDseRU6adetq3dslQhfUShg3aMPbSP4yN4cGiwhNO9CZmLVA
UtUeyjyixyhnB2BMwBK+LvUoYy6bhw4CkyGmoLfnWHfCCZnd05sHgVGxhYgCugeCEzSWisxjaG0g
W9sR/SFAXSHC9/JGzjS+8g3pS2gPKJUevwjuTWR7lKXYhcrU6u6Xmeor0qR0xpllP4F4SbbQLtUD
LvmsDYIcLTZ9usbn0HwAIEC/AB6K0PiTfYpybMkK3L7d5zbH+qO8d+yrl7mRopUMA+utSkB5jaPP
R9ocFVIA/lDp/tYldzCJwOsIPSPDWzHEdjsInf5WKqb/inJ/qTJFee5YjkhKe1DDEWlIKp4qxmG1
ovbRsJPiFE2z+IeLa65jmrg9lDmWQdd8cuffQSYEei4oBbVs4JiNI4f08wS4AyDOeAf3Gpg/R0n5
Pe1EVniRMtkUer++vmzSjKqwacHUzqDXv8SUmv+/r+iHoZkplkMijinBkKzjx19NWoju8UoJU0Qy
IQYzLXpvhMW24p649NfqoJseUFCQFPap0XhTuF/NTS7xJ3XokS2jj/QmgCX33VuUTalfdxvhR+z0
n5motmhyxdCnT9A62CVwak75TiUYvkQczVRmoQKTRAd4UNGTZiDB1PtkfBabyI3bt5JHMcHgbsKk
l8VZmqhHkLOPXDkPyPAAJsZSUf26pNDoTvaKM41SADmm3jvISosgqZOUQZEy6+Gyi264CVwnaIyF
g2Acjv1KrxcCsfE3Yt2MJBO90Ko2FwRWizmY9wrJffJ3nHv6JXvtDINsJYAdkUVkRoIFdieCGj+N
Ev0Jh8es3/cFAB5sKKzV6qbZNOWi6HyfVywMbQN/rSTqs8MBJ1cvPCs7+6tJNL3g2HITSrgQCSSc
U/2R7njWyViC09KTYYpTdL8C9FOg1oxTMfOc+XOdiD/dK5z4kRr0JcLByNFuW9TMdFJdBi8evmY+
E1G/IC3PBc9cZu0V+3j/FdK6QW/edvrlRQBd/Wt1U8NF1xEbYUxFw/dnd+S67vcbu3Ez3dMm7/a0
i3tjztcv6b5wEqNUvGzxMut1iv9L48MPbH/qsjjFTx6UarIw51mDmhNj7a3CMG/tuP7pn9E1y0Tl
7Gtz/TQuVUDX/E0Ex+M9EtP4v+gvcxqqOp24qHTaFNHQtUFHmN23TUpc3PnnSKXw+CY1slRG52Tc
GWtildo0KiqTEmHbKqr/kXg30HN6ViJaJsMBjTAVj3bA5A1+vSaMlCboGX7Yg2uAp8Sd4GRiHlAq
7bz/aiVNFa2oH+EiHANQ94D+rA==
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:22 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FVbI+W2ezbUB5aUxmoiFOMYFcgtf81isRUFomy4yepmXwmRsbrpDVPDWpzxg3vL9
XL9TW2AnlDkUzOhSrOwly1wyK3w3R/FVaOGNUQ0gQ5n5HKWQVWwxR4fUKtDTK9G+
Rpmk0g/bIPG0ZBSyo9zypaDStjZer1rqkIe07xZ77NM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9104)
iKxRuqYgvcoRQbK8B700P/lnFj/oq6ykOqaOmlHGZLYpXJ+2HH1viP++rQUBHHRO
6Pr25CqxZKT2S3Ie+NbT6e+iR6heSyJpjv/ZNlrrq8DrMdo2AjxGNarYLXrKDgFn
tZWkIQxV8khPris1hwt2MvpCWJ3yuKgbIKqU/UjsyomBrBeCelBqLy25kki/y8s/
vznplD8X17Qak9AIeSXPTT0EA1rQklkqzT+p4D6or7sOJfEv58itW48CEEltN6sK
dkJyZ6Ak4DURjWuwWSLFtg8tKfr8NYgjJ2OEhCRhb62Wga6hBMXkI2R7pNyO7MW1
SpLqnZ/2dfp6eYHP4j5WbwiEZPV29vCbsvTMy7vRcVviWG51kvFNuHbZRJjkMqYE
/p6rHCd6rf4UXyXXOF2YhOoQzTsDa+dpI1yEZpjscpRiyY9cXJDSOTHN/L0RBlKz
i/iVhmEL8TGt2b/cdoo3OtQ2mTMUNRSXx20wtH9RyhZ1wdyhtwIEvEEG6xKCKtEq
Bb4p4E2tRgA7mihHTy/Mg2byUDBSW1BAnWs7WgOwnaEo0Mj8u0iJCU/+XPmLcZkd
7zVLORBLbI1JD0zNel5RSwZMZKG9kYZXxjG2SAtuzaQHiYVXH4sVizYQzz79X3rU
mmjJqXUccnJNv3xmI7Yp16FN87KUCxzijHTYl7RUnXBsQYCdcum8bNw6g2DOzpTV
kLh2bmYbWFOMRC4HWe/ObMAlG00WHjXdVVqnm2Z3cXyTUxFSnQuRYjanDqngc2Um
gx7jq8uTsUDu4RdIHIwzJ/2pzOD1kj6SkkGR2+Q5n5FXUP75uj0Q7VW0rBj73kBX
oyCeCb6FMuMxe4LLrUfpjhD91584G5kBY8b5IqiUKkitFybLFhoGHGQDPhXBEZlC
nsuSxqM1nupm6kHT0ZFscMM2J/00NohwzQadv7M2MRrxno1QamQOOkzX8+7nJ/GA
1HUJvYmFpBB3eo0yt+wBQ6DbtJuRBU+3VnKWD/UhgRTHAdQAuq4pw6dh846dlDVQ
6CnJcjOBdLhkRTEU1JnDFQwleyJkJ+wR4klpa4+rLsv7mc/nS60Jb2kBIf+Qkta9
MpmEI0FCtxs6d+kJ+itV8ZDT/w6zQnQINh8Ua+khYEM9okqke9dUMtHYmmWED/rA
kq/Ruj7TAYtfF6Trym2GLQwx+eOeJAqf5b82Vrqkq6u3XaZhVNymlGSQz5NUIrTS
w9kyDdhf9UMTVrV19R7czd2LMk44E6y2nlolEkT24qe5thfeKEx18j3aFCVpNYqZ
Ctt0uewjAxssal0msR/d0ZHgRy7LQwZFNHNzpP5wz+94YUfG/t8JkMZBO+S15C9j
dQ85HNibpQzvXISmcadlDCok1HAIkBz/d2yMXmY4pNIdbkncQGsOP3WcSJ5Z/XRZ
QuRVrQOXI7mOuMsgCp3mzOu3Rv2QDY41KgZLTZqZn0kdNOHhr7VJKttYofVsr6me
h1BbdiuqnthWAjZ7WiqyKCcZR1M4QZCM3aj0qujP9AzwoAJdulAGpF8GAMsrzX0H
AdatxVWhMyrCRFZ1tfSQ1mOKhpa3OAlQtxonO+p6X3uwec+otjlOVO6kUIv7N79b
7NWJBSmO/BGA2dCp1R02T29wbQr3IhtAB48CRQYhR5PseOL/uZFfkbv69r+vnPVg
bQwrM1lI7ysSLmjibJaCY1VpRP+HqWskvw2IAUcn5wB68X7dY6qai8iqZJHgLMoO
I9v1NCXMFgndLlru57FjFQose/PMQ7xZkgbgyaADQe8MHsl7Ip0qePuOvI2R1nLB
RtogC3NDdqI+0mzfFp5LlqStZUTDtmPj0S3sQrbXps09OVpm5uvvO4RtF0SvC0wC
W89fEnxbm2TCzbqp6LvbufT6xw/65mHRfx7ZOTBXp7hOlsMpemj+FMrje5r17H4n
9Lb0RMwqLn0b16L7fu93vAd2FPPvfpRyhjZ1occKy+FIHmtBpkT0GWF7lqXN6O7b
Wo5j5nUHx+H+K3FZIbW7DsZIkIYfnVpTQRj2RJRKW14fyOnlatZFkP6VYTepE5F3
bmv5nqcpHhDDeqQUHxp91JGYrfj8OItu3l7Md1pTCR6oMAzpIyUE+o2YfAAF1IOB
Z07aCGpF2FRvZuGKLaz10V6DnVx0UIpjN3trzKZeRiKEKryDMGrC/1qQN0nsB4oz
dlhGF14oJePznEqztlXRzJtUKNF5DZDaoBxZwiQZOW6fLpP8Lq53oaIaiLioxJ88
lU/dAITWLxO4whZpvpKvTUasNorTu1kw4Rn2Ho9eaVaqpZmfJXKrs1ei7ZdZikwS
hW/kS0UZScsEEIpWXfkSi49tGxk57YRyxy7xdNda7TIcq/fpWCWO/CYMYI9fq9x0
Mu3qPrAeiGgb6WGcfVgrNnza2ZCYUdZauvASPluN5JkrWq15Lrsx+FkzuiAZtT8v
k9eK2EMR89uWSvHgdiCyavAbGexFkltUyL5Bd5KvhlGXeS1IxxwpXyuadovrVkEy
StioYmGZgzUI5dHclIlIIUiimW1rzdFdwNe+lTSw827fUvZX6I46hA+u2nS1HIXc
MtbedLMmVD3kWFrAkSnJXE8Yy1h9MnPmTw8ZHu23ImR3ZZjMEi2gNHuAaIpTWkkN
/4vn3SZmZnLdp7FCRAREdt/WN5Tg9rnH+avHCv8mUAIy8zBeEoyO8rUiDhlg5qJo
o3yu2sEgQLlu6cTaAHf2f/xHlk4MK4xAehX6Q52cbXaZbvDCq++mKN0QpyjvcA0A
pqf4dQ8tjKfZVcMijOXOX2hbCCa/xwxjWCfYiTsWR5PC0xkWCLWRQ3ZceVUvZJXJ
9rl64Lcd8/LADWQyM0R+yYBnO1YcBJuUUpaMiUbaUkbugDDJS/HxHpAZwb5lwLWl
NpEets59tVY1KgU2ASag1RfVx5NlbDqkagQf10lgHLga6HzyP4G3nHymypL8QuoC
G11oD6ZBp51GPv3AkULkBYyojt1oHJGO6wJXTUKG+89mWkiVVhSpDnGdI/chMxZ1
fr04IhfXDGvFMxu+wvno+kyMVy9rWujnaDsw6hOSjiAv7Un3o4zPjzXs/tVsAU/s
zHHJMeK2/lIVgqM/xX/YUsZatZc++exE+rYvXShLAbK89eY6IE+J899cGamMYxG3
p0+3pISl7bGLMIQ67NZxWJSlH4RIb5oFjeMj4jVaHggyNMipGCHTHt18Grt8Y0Vz
tQ5VxSSlZOTJ5kfXpokIb20E4nXy0chvYuNgCVvte4rNc6gB3HBLcc5rn0aHYONK
uaM29QFhfK0CNvtA3ULk4Ze3/8TiI9OI5V6GXxeBhRj5mfKWnT0WxKpAcIaUElSF
EHIHrSqE6jg1fIVSjQpY8SQQt665NUiyFxmXYJT9blSEX+X9Kc0VwzmZ8VEyWM6e
uLUkLivNC65KFEIeHzEa+gGntPgYm4gam16ArQAg0R/+dD6aZ9HGX/aPNbQiAxRD
eS15yhAL3rxNH+03VFKFMIKnWk1RNPhayyuhvQiz3jOTbu0K4aaikX3oE1+EZI74
PiDmqOjdElYx85cWLKMDYe8zxFkWcvwQFGVY9q8j4WBNQZpZB17xX0MOxknxqKlq
a8kCGT5QjUXZM7i9vDXVhSP7gbZfdb+T0M+fEJO66/P5D1fMjiBdixfTtSIbX/4e
vBDoiWWDO79zGbdlpkkmLwGxfghqYuazbXvDEparnML0LfGAmHzc7u19+Mm+KL7d
LzTZfhy2aEU0ohVsHeGlH3fkzjTF+ixthYRKPS2Nf+FlTimaCS4NBPLu60UWBBPr
RVUAMIORn9if8ke92CJsNyJQb0TkAWo1blbi8hb1FT2rlGsd39WOyul2yTi+LACk
Nijfv75oypbyaE5WTyulzIW+ZCi12uRs2Ts5c9nxWFsWGlRb4inUAKTEIaFYaEDi
8zkGXTDbn8tFZMS8dzB1JA1pYTjjtEjcXQz8g4p1flbKhPJgh4FBmEkUfQAizU2f
20X+QNIDeMK1sNUdeyUoMIwIez37qA9Prp7Z/Ct+5rsbmu5sCVn4cMfB2wRsog35
PIzmsMqusj8e2JeQl4fGKxqCseagPSblbE1H/exGog2HR7VZxUWomGOReSRjXh55
yZItw8VlrbTnn7ftXDAvfcds6ze98SSAgM/68gOFXfEgIcbPhTIwHe2zbBOzC9Go
NupxkIXMTsk1HweFvX5wHYmPsMflhlzErI7r22AQVPF8vXfxmZSqG84TXnPj21Vm
KzE+FCSdJFuYgXP2qHIYqPZGUbVaTA4Z6Hv57ss3MsOXfEzx08vpmzWXBH3Bf2CN
AEK6wO7kzBjwLhHgfPcJpE+Z1BuJsqFGhlczpDGeMpE5OJP8wsKsk6+y5ko4VtWt
K3l7mhiTbSJ+Hlc7KFFhtHVf3tjeuTWTkOT81yhoVnHlWiQa13yF6+ukYUvx7FwB
pRrY6Hm81JUn04WtEzdR3aYNDnBqxhyWumnHm3PP2OYI6FwSB2AitmN6EoLVaZCI
qp2ycVtpgUplSFtwvdhLFGJXZ7FkEZkdP+EzZmQ5VS80A3Gbaf18kz2V8D9GvtHl
bq+mBIYy9Mab25lDZaqpkfDP8rsZLNDE5TCqH5Phw0QmIV6u86mM00GEUhG5F/b7
L3IjkUA+CCWDawP3/R+8SpNVaAwmnDtZSI5T2Z+IuhzQ0+QnJjfy70JYtW+A4F2x
QA5mOa85a/pPiK8rjVpqvTuLDHx1wS4rCQLpJ+xxThXKLBswA2ztf4KGaSiMlGR9
hkqT2Jgjddreu2Cd5G/FbP9ym1kGbJl1UdEdk962iIARc6Yl3ACnckTTbHPx8oWB
44v6cuU9JHu9dBVkHRRfIO+pV4pkWk8C48lI/u8HqNIKE3XMnqAuk1XcxrlSqNUp
8MFvAbEr1fp5+whzHHMIH8hQi93WIoc3r3+CHoK5W4tKm0SzVCL/8/JeDw9szzuU
EFbiF7+u5mWWwr8hpO62UaaCE0oID+tA6OYu24wgcDBKhU/HOit5RFSFbqAYbRdP
PtrVP7ihgyNvW1y5E8tLMmR+hMVcdZ3abNRVOFYymy1gouPd3QEPyiC1d5IT83hb
zhQ7GhBk1rL0CIwY7VQV5nRmAg+CupP1vqF1INuutUP1fnBv6UanPiCrYsZYBz0s
zB09QsnsNlw0KcpBz3hlHChYuj1L/NoADoouQXZQ1ENOEnJOp+lULxy5/bPL1ulZ
33z64e6tUfMvYpyJXkSQ6p8HrubwuSVvhDyLqLIJ6PrRRdlkftzMEGcIfUnmmqeS
qEylW9dqndaWSpuFuXkgEAYLv61FiV0EoH+VwiP+PtvjYVFRuhVnsvbmhcpT0cjB
lxbqwfkEPx2tSWRYg/7HbtzUMtqs6Dsbmxz02jL8Y/qLqMItbtxTJbNuPpPCHUmx
CPBPfJSMvnvw2BSNNsdXzEbaWJjsmf25AZ4xhlebd4AqNFhcCu/TszpZSey1qi1A
TkF3wGKLLW0IgVl1Ek9DyohpstFF8MUnAh/N7JnMb1TNlkdlmwSzSSIzA3Qafu4a
f4ADw6ZBZ52qH/jKVDtOgdHH6e7R0PhzLvsGyLO+apkH/Xe1TOZwzbty6GKLPfSY
/HJD27xR3Cj32pnkNMEbnI2SVead4WP4SLomZPpFUe3kbxYeWflPUr4r3zajoYH2
eGEz1fHss4TAtbyI2PovwMwcBz84tsTrkoeqiK2AWnVuxUxZqD9BiDHZ5M5X8Kx0
/Yk+jHxqFHsuxByB1hQPaKvVvTobwAd2SxDwA/++OvuPqyLSLevQfroDQVNPYK4N
caMyJglyVGAIg3Y3inrtUtv8cTWMFRMBvnGcXrOdF5OG4cw80gebapHsiuezPbiQ
mAkWvUkdpyrZ0EjmB5eRM5MnKNkMRU3LJ9clN0XhVR56e1avEMAYBFzi7+wXPMHj
OqyYW7cGjwSB920nw77TyET8NMOypP2vqVYdJJflNOFQ8B6XV7nsVU/doP+ANdNW
qmEGtVMuOm7BFOtxaYXJ2okI2S1hEeLX0HL1p76o9V8aA2szXGx47PlezuABMNc7
u/fSl8XUfNAcpMuYQTwpWLRB8o9vuHNMk8C12OOqs5Dup5FX5axEYOCAMdPhhvnY
IfWL9ONXPmCv0J7/M3YUs7IeWqE2IYLDUDrKS4gczP/XCTgxE5JmqOhFeDAn9lcS
Uh9xE3RF/Z83PZ7HMtsDsAjJaNVmQ0BynrObQTQ27ewv4qj61izPuuVABxEWKQPR
4d3o7c4jI/qO9b78B/UH6hlr++ZEcvpgtyrtxAgT551wtUIOhd96nFUS3VacnAbN
qWfOj2QgSvt1Kw4/BjS85sL6BjggipfpsT36qH7FOUrdW41b0XKai2oOD6bRmmhH
Wsi+nLLKuQ+7T3cYlPfU6Ls1faoEj9CBzDB4Zo58jS5AwpncpMkH93K7ZA1VJLYC
QVCpQoAtg3rTCIck2caBoL4R6ioWi5pmOZx4aH3jR/LCRE+0dMKhANko4Se2ijUC
jU/GDG+mnAlAQ3d3UKvNo0C4zf5cO0sV3O8FKZjwShqrFqazcfK+GcbMLgeLiY/4
AfhwSQrv+AtDpV3Gvk1YVxoVu4aWKcF/+Y54Bu+nI7pxfbFyWDtR5+BLOOfSjEra
WfsH8fEGJc2DukchTceMnNvbJB3G31BLi4Z/EUwoIGFVjaW7VGkE+tuLZzdWn3UB
jsQRF/zxuL+oZ+BahraIpmnc3t+AA6zcDuU0ucbUlAGMjUdlc5awZFqxFT9Myyhu
vW1NAm5RhRiHXBBs5WyU3LqyUcHIXg2ibRGmzh2sH/GgmIG+0kqqf1ibq4Ssz7ZR
saNHE2GXxNix1sgQ1BEwg9U/AaXJPdtlJXBPiLB0xgTFvxWpnlqn2EdSsy21lawZ
wTYdrY+98f4xvi9N+Pbdek+r2wvmmJv6DndJDMG/5Hf43LcreaeWCYR9Baf5ue7e
xqi62Wu85ESs3yN6NIOt2TIbJaQblJOwHYnZa8B6P8Q/eIJ8iN3oLezmylDWxmih
OehiHSjGftYC3vSlGSnqySLkFJXDL8G1U8TwSLXWt2UL5YxQm3RR+rckD00z0vo1
dLjXPZERGSsDjjc+S00mhc1RUHqk4gP/ur2HNja3N20DVHw0VYROvJJRf7ygyyF2
tUGonFrUbTMholIsHgW9YtzkYVIzZKOWliqH98ryWGbK/HC19LzrP/taTQkGjgyh
ZZ5uHfwOy9YyXijmUaqV15xVRk8/vi50PVrYGiJ2ZzDQDIBJ+g5vB0gCj0cnLtO/
lf5J6GASq8nWjbIpAJnEP5CttGGD6cQEFmkhX6ThSq2lpHov+L5MdVug+ix+ErVM
tYCw2mWdG492tNqoP8sQXE6KuvcrsqqKL1lUWhi55BFooDmS6OGsbKZchUhuD12v
er9k8k1krEYllUKxzm4pL1aJZCJ/39D+90g4z1EZaUAO87toQPXqovijQ7faQd6N
WGLQzexZhtyQ9uoI8S8GAAjtJKmqL9DirrHFCKDHF2OETcWkzisZ/L91HHjSzwRV
KbdY/aYY7iFe/oJnHkBzZ41j52CUIFGDsBNrtlV5ZS1VWgF70ue6nWo07zfHnSy9
8yoFckWh8wANmQTH/6zwRLZ9xeeEToIbAvDIT9KPE1+aDX+QQIspYD6ABffS8ABT
ODhWyuY/2IZgFzu+fK+mQkcjp9zUB7KMvaYZ15RC+xP5TC94ilCxTRyZmX6IOjAh
2znzQLWsYP9fQhyLrkYZKNtrYrwb7gx1Q2zNUHmcG8lgh9uJXsMGk9ourZ9QbH1q
5z19mrvAUWTveBL1l6HKplmJD6G/iF6KQRVpeRa/mbeWTgnQEikHiGWkqstGmAgK
5pCqxeCCm2SRcAR15Z6CpuSL0Q7MW+8CmKGkzZ+G4RfzVnPZ1KJGtYts51ncd2NR
WVOvofi6oIFg6FOe/wnk/eioeIQwjZIac+pgomvJc+lx1kYfxin7hMAHttaoolle
+2tzmFV5+PUJlSofMMoKMQr9nN+TQTwYqqucwZ6FkqPjnWjdvb9fWbassTjKFf9d
9YQz0JLv8fMofMXYGpl+Pp5+smThvP09MPB4JBCuB6Add9kuGVm3N5lh0mrOS7SM
ZVmJxbjYsmVIBlD3oMPUqKbHl8cPe+jinSBBOjRL/fN2tGmeXO6ymgj7hnYlWftN
czeKV5yW0AxFNUxcBQGEqTJPmhh7GqEcG7yhr8zb5qLRWAWdsoif+iLO6U1J8q5Q
IMsu7yjiOe2a+zGTrjgimJvtFkD0U51i3SAiq/08ELfmlolDaQC2B5W6ilDk/53E
cS8V9BITiz+LpAdqABTeeQsa5XoWscibds+8cbUjCnxxjcSSRvCbyDa2OQq4V5VE
zYIm+3/xJplWZdFZs0ikgmvcnt1isu47Usw2rU3MysE0H3asSEZwCmLgEl+5KPFH
cQ08diycavcmkCWpoB+CV7smMrth+P3HX9VGbAEw/ET0YG4PMrDd60ayKM9bXu1p
46NHk/wsyiRuAJqDMfCg6/G9yF4sDV0Rct3nYXmyZ1iXKd6eQaf53foERcSw89X3
cLvsopNCQgqZO4OJhgOCi0k5Kyhu/efW8l3u5gVev5TfOLDExNYfIRUWOOYPF3cz
lBWnCjT3ovHxQlj60if96Uavy0W50TC159rwv5vU18h9yRjHhYKkJ6XDV8EqvHle
U2g+AFGFt1S0zlVoRukIJGE++aWu/avnm4ahlGDnL7ENlbE+zysMTZDQtcAXfhxS
5fLxFAoCel+hou7CBj5k2G557dSdfUwMGm0q4SpeKyXMuKsOFhUDAGum2MHdJJLR
lsRtxiXAKKCjvsxxb0sZcQnum+lizpTxLiYMXovNOedj3uoSa8j+w41+BdSodoc9
oum3pTpXp7W6QzByRZMp5nyzOOff8IGSjxxMjnsh+HxK8kkEPpNFA6IrxEm/rwIf
0IoKQuan1IRYUmE/6vdOy/VMvXcNONBX5f5b0iRd9kmPQDDm94FYncgjxrsIm2Xk
JGST8OzK8nQSKgEkWYPW72NKHCeruApEtp8E3Gs3js9yvcyLCcn0Y2GxA3veW0Yi
BpBsSCAAJp9PdVb0ozrl7Bd5Th69pG00Wx8d6P187wQdbJxTMSYhIsQw3P2hoUJm
KyuwVdcj6yiZCaliV8+x3CIILrH3ZBFZxJyvkee/UTgobcvOyLCMp9mILkgarPQG
dSL47pe0E35+hAztpDZuCc36K/lkbWH7r/r9whknqExLyntAOrq9cTusMUUM9jSo
muXQjyPWtO0sQ6QzolrtAIEYCwoShTBTRsepihKE1IvwkwjEVRDIv8NsTsimbqTF
qyV0/Zk234hfm0SsKQokbBN+yMGIUdlE92PrLShwoHucQLYdHPbmiJFUBH7kHhv4
TF4SW893PyG2SpNiPHbdt+vud0Q9pt6GKaF3pXGbJt1djcmfJ9rsWWltwmHuQC1a
wBIERRn14eufd1wfZN+oaU7ogNJGH/r62Ws8iLyyE+wObIhiCnIjK5Wak6XR8KMK
YhAN8pmCn+rfmCgHbL43TAHiKys38totvSIVv36yNLw+Ni0qs8yDSAtut9M5FvJ0
oHHYEjP9l0O/ZhEtaP4uadZqBlXn5X66wJXSZeCJ8xb1nVijErU5OQpjWNTYC1AC
SUyqMcD5NSNh3ljiCUZcdRMv0X1qIe1tOY9Zr6ioU3Tioc2itttTb0TiZy9FTc77
oYfEj/687oRWD3c5md3kHKnA8DKmOnr9pYUgX6wrcqIzT/dAYEQexh0Hp89+dbph
Ky+dmn7W7pUENV6rWEOANlI4AYckNWhlUtW9+kBQwSMhpJn/Hjfv0htVjteEzJcm
BTsdWMMgWXAQmNX5Qletze6Fd8eD9LCYHay+0lw+Z6Y6APxLYkM77cL2eQ0jsTbV
fvxiabOT2KV7bcjucgHkhDv+T6FHZals59+wpH5HqsjJ7V2E22oL2CGXDj5ZTLvZ
OBT9To4jM2EjjVw+1ll+KlmzZ6Bnz1RmVV3dNL7kiWS1l4bu4J+1gwYDIY4kFdTR
HQywLMhYxvzLvlrxBMRRCOAC0nfijpOuRvyw8bLjbNmCFRaY3Lx1p1PAJjeaIKYf
6xfKJcT5V4IqAvuLN5nAuw3mUyVxr718UH46KGQxCWrE19A40NRWwKe6WtBQWPzf
VQ0+fiYqPdHdPSd2Dcm/naAl+jKtIn49A08RShNhvpSnjO7/+rIpS/WfX5/+GOvg
6aB2VHNaxly98H2iqFM4OkMbnnsJWJ5YxnDrrr0acdfjpkoGyuch4mBZXiGlVwH+
nj+8M0YW1N5tQ7/6fAhxSmA3ErP6lrZfglrBP7kZuHlG3FjND2X4sjUJQNxo08zO
JFbgy++g0NYTH80Ai/AvAfADpzu3IBTowOp4+9SAGuNHPhxdKM56+rW6U2UcM988
/LN/pp6m/4lbPVcKPGD8cN6Q1AwxUNIh9h/MJ/C7Su/j7RJLwy/1d+f1MdM/3Q/e
oktkb3TskZ47AeRr4qEqNn0LT+Re5o6twcWB2ZBpEnUr3PsDX/TQcAxuCN+nP66l
qifMwuc+75kxH8ndvNJPWqRvhFk//WiguHmlU+u8Q0Y8u0f+BwCmJSe1FVZIc9eu
yyJK7r1rc9qa3/ff4sJxSDYLCgB6LV94/9r4NEkTlNyrx0Xxyuw4idS6NzwctyYq
9kMpjBviAFnggli+MZHlpYh1Bj2NV/b2KXPCx5B8jaKibXZZtkYJxvqnHfVrV8t7
EAg4LqJ6QiCld2076IGqSad1dp3wrqetM4inIXy0HJyu+qgUA9pQbzT1N2VOvEn/
C9TzNyH6UIDklLw4GaashHuSeknfsJV/e2Uk+d9Ds2yxBE+qlXcdgQpQRiyPlMSB
WsGeIfJgGEGH8+ErEOzYtJsNTvFcHgUljn0l4CCAyhpwVOumQI8vd/M4OKt1TUId
X0x8H0HZgThniB0zAJ7Afp59to1t8RYKr7Hra4CNrrhoCgZaSFuWH3qDSDN4+k+g
6d92R4z6Iy0SAMIq/CG1lz3I19cXSNArvlaZP+iSxKTCEKlbKnyWWKKAWqHbMJky
/EAooUCiLziGZHNVIjUv4gyNFNwzHD92FsqjnnrZr21V+yB2p8subWDirgm2qr6O
j5GI+bgHjX8FzfUgLk04WipQhmSQpAYdK/k8SsQ1Q33CgQVM6L2yWTOxBV4szw41
8rcqrbd/5FG8qz5CYvxrabgNgyDahZBmr4c+6s/AYZZVAPFecjrsCE8FVTcjGLMY
zvELvmyfnNp61b7K1Bggb5SuOEo4XdHs91/FZfE4qZDjUosu1nHWFCuQYvGnRKOu
T9pJY15ubFIS/HYPAd7wM8KpeRWRIZTT3wIqY/myenxGcAi63v+R1wI8ZTLqIkCo
0lHYmB8j2ap3Xb2AtInpcfsHOORcJZRLIASCVj4Xkmvq0WwUNmJaqe8Ra+REpUTl
JrrBVg4X9PvybAnPSlVcDlQiQQUV01JayGyY67nny8yAT65Mn51tV1xsCX3AkRiU
6I/dPkvINocx231Zw7jT8vxg8GT2mFY5PE7ULFUToqGXcmlmXTQy+CyS4plbRr8/
7Vt0+HCOz8WrUK9RfsejCuYClBdhC9b20Bycr/QKa4EoeDPhaTvd26TDGsGURCpk
FntkAjylG54d6fFRE5c2k6flGI7cKKxd1hXKcSTOfqEivENeJZb/PQk017gAcP5z
od+vJkqVhUQkObw2jVTN1jcKPlziWwkllRDN6HXZCqLX8vQS8a0okJzwxbjV4F7Z
yOaeuk3yDXpTz9kSbW6gHdE6LAJciUaFCDELNXRPAEI8S3HNhR9J4L9JIrqXdBKb
Xvkf9tVKOjusA1z5kq2utk9/YImiyp2DRYD/T9pfsV74mw06NcLoE7WkTUONbEaU
cbLOSmn8hoc+sUBcFigeFyx2VCyfe4/+ISzFhmh3ueMtRHCPJ28g3LoGQ3MXGrxO
1g9tdgjwBDEt6DoxECIotmu+ZZ9N2DPrru1+cDZT654V03v/jdL+fLI1h9fpNjHR
/sESydLwZqYxW5BAeciAFhJlwl+FHQ58AHmOBt8fkZKsz5R1voTh2YVgJ/gknVr6
jILDstqd01mFL8brMmP74XVA4HhfJ8ga+Z4J+Cs8GYDwHqT6ycXx0nGPTQ9i9X53
7d1e9yaPSdw7h6YZ6+tE506ibKDy2y/hQnZQgruYexc=
`pragma protect end_protected

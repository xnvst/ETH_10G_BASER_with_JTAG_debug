// avalon_dc_fifo.v

// Generated using ACDS version 14.0 205 at 2014.11.06.21:36:38

`timescale 1 ps / 1 ps
module avalon_dc_fifo (
		input  wire        reset_ext_reset_n, //   reset_ext.reset_n
		input  wire        clk_int_clk,       //     clk_int.clk
		input  wire        reset_int_reset_n, //   reset_int.reset_n
		input  wire        clk_ext_clk,       //     clk_ext.clk
		input  wire [63:0] dc_fifo_in_data,   //  dc_fifo_in.data
		input  wire        dc_fifo_in_valid,  //            .valid
		output wire        dc_fifo_in_ready,  //            .ready
		output wire [63:0] dc_fifo_out_data,  // dc_fifo_out.data
		output wire        dc_fifo_out_valid, //            .valid
		input  wire        dc_fifo_out_ready  //            .ready
	);

	wire    rst_controller_reset_out_reset;     // rst_controller:reset_out -> dc_fifo:in_reset_n
	wire    rst_controller_001_reset_out_reset; // rst_controller_001:reset_out -> dc_fifo:out_reset_n

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (8),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (512),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (0),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (2),
		.RD_SYNC_DEPTH      (2)
	) dc_fifo (
		.in_clk            (clk_ext_clk),                          //        in_clk.clk
		.in_reset_n        (~rst_controller_reset_out_reset),      //  in_clk_reset.reset_n
		.out_clk           (clk_int_clk),                          //       out_clk.clk
		.out_reset_n       (~rst_controller_001_reset_out_reset),  // out_clk_reset.reset_n
		.in_data           (dc_fifo_in_data),                      //            in.data
		.in_valid          (dc_fifo_in_valid),                     //              .valid
		.in_ready          (dc_fifo_in_ready),                     //              .ready
		.out_data          (dc_fifo_out_data),                     //           out.data
		.out_valid         (dc_fifo_out_valid),                    //              .valid
		.out_ready         (dc_fifo_out_ready),                    //              .ready
		.in_csr_address    (1'b0),                                 //   (terminated)
		.in_csr_read       (1'b0),                                 //   (terminated)
		.in_csr_write      (1'b0),                                 //   (terminated)
		.in_csr_readdata   (),                                     //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000), //   (terminated)
		.out_csr_address   (1'b0),                                 //   (terminated)
		.out_csr_read      (1'b0),                                 //   (terminated)
		.out_csr_write     (1'b0),                                 //   (terminated)
		.out_csr_readdata  (),                                     //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000), //   (terminated)
		.in_startofpacket  (1'b0),                                 //   (terminated)
		.in_endofpacket    (1'b0),                                 //   (terminated)
		.out_startofpacket (),                                     //   (terminated)
		.out_endofpacket   ()                                      //   (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_ext_reset_n),             // reset_in0.reset
		.clk            (clk_ext_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_int_reset_n),                 // reset_in0.reset
		.clk            (clk_int_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule

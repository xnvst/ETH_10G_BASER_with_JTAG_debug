// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:26 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NGVJBeKzXL0moA6k5MGOqQZvowAPAXjjFWLAsF1NFUoYLeG+Tm0f1hbae38CEz9i
aKjjMutASBwe7oaCk7RtShsJLSN2eJ26Q/XE0tlvZukshUGouudPxsWnDbmapXL7
tP7kN7pstAQQj3tgRega2nhs9iKLA+akB4Th7LrsrWw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12576)
3uChC9ZyqLwA4iXeuL0Cp5i9PtNEB4ezfthZPVUSMkJa+keAZV9WB3OX2PB3Xl3v
l0T1ZYlbAuvbYlnl9L2W6DlSv9WKtV6hEeToye8Dlb49VGi7gtd++VMskhGERuQK
/7VlfQhwUeyaV+QSMIvkpgO77/qqZsOSNDuFwluIqlyUMb3zvbUYlIhaCd5aUzA8
bBLHESMQyhn3dS1E063Rt+OsFxbT3RC1VZjaGHdmGDSBy46l6KE+akCl2Wct69CL
+SpeoVFsnwJTiq6d05g5QkwmHkTEZ5AC6mc7cWvFjWmi1ZtUTbWB1drPMfaE7tGm
gTw3MQnNQ+2dElAWlsQ5leug8AUPhGTLWDaq318F/Ujgvoxoaotb3PJY5QB+Er2k
fWKgLKJGCVUPHfILEmQ1B2fVAUtbZ/Yg8todpljmmL0q0pTwg0m9bOY5Gn2pLMqc
pg+0jn/OSQy0Wv2BBduHH834C/YrzkC3McO/MDJplqvQ1LAFFzThhopK7flEPnD1
8KpyKxMp7Z7qsHvGqVx2ofNpzbUspoNJD1UHoSqUXE/CuTsHEjif89Gtcqw89CIH
fkvWNxCsc7jGEshMYwA6enakE2JT0/HIes/StEG99b/CjVk4JEsoycpE2xKK3H6i
UwkAqwyB5gQD4FdhYXLf+DGqi7XE2Q7R5k2N8BLPaTtTI7ZWo48Pqi7OvI0gvqj/
RdbwUW42fhRv9LA/NzgMkzvvvpDaZRRywRV60Qj6vFmrqGvk4FIGE0+aahM34Pxz
ykq073EIiN5B1GTegn8ruuo3HBSkoyJvI5icqTnV0nt5Z6jenGAOBUIONR7Id18Y
1brIwGsukonHET7nXdKMNj8gcYlEHgE72ZjsHlpFmUlfqzAxt8beIxnN8h/qBSN/
IgwUsNGrUTLzggVW5MXHtvg0qGryZTyICw3quuarB92Dt3R/NE4hqWvFG34NtzIO
Ho63pG4PwYrBwjON2vznYWh6zeHiICxB+M+TRzcA6CaMQSaGaQ4hG8d4O/RRWOTs
2/1PyMm0rqgoZsIVdBbWxwJb1NkPh9Sr6IdXL5nW3dK9ys/87E5g194oLoMpPFMj
v2/mNo4l3o5tRC7VTPGbOHUCAVMC2WrWJJcun+XMY2KcxL78CurblZbc3cKSRLx/
k/c618jNub2wk+bUPO1CYWG2R+BLAkDvO0s/rsnPJ7WOx9OxQ0tjsUH6Op0AnuK0
F8JH/C/G/s8Oooj9k8el/25Ca0AdQF9/m6dXXOYnYZoS9QfEhajXz4p4NDdPfVkP
b/V/xermrrhv6INom6Ommrnd4uLmGE3HKpccOblPLMb90gFE0QL1HmSiwl0fdn91
Vh09SekzxveHkDiUJdP0YMyIGhiGXFbzkpRJNGje/SfFKAEXKSm52OWDxkaHOItp
mpdOKrtIylQeaQJqCRSx36Nvorpal8M+/hfmbDo0Ss/4JwVRWojlQEh5zcaJDZsP
YApmKzEsdgijlhaa8qJcmeU1z0LQuoW8bcMKhkj+rN1Lpmejw6r68HaTqDf/W5fZ
s7VfOMLiL4hmXTpoPJFhJonLjwyy9/LqmWowrh4Fky0iN1cP975W8MbKG8xAfWbi
LL1GB+JJYnlJk1cXnL7pXThvQe+v8Lhd87VfUPm/2RlKztZe0EC7iImxttol3XM2
Vbm9dKrOGNV6VVUv3ICLmgQlt0gq2ZONfKppoBMDPYb5PwMXiSQn5kMhO77jd7OZ
Sdm1rcIb7WchqaFLJlrJGXvrSAjQIc2eIeAii82UhJcwk+w3z1sgVNA/G0KEL01H
Qp0XCnv8Ufh9JV2eSmyEH+Iqf28g5CrcFJ9hKep/vMytf1VjBBFqDuykyig86JAB
fexhUl7x61yZF1ZSWf+I5reRzDBZ6qg4s2gvCo9cPVl/q8cSp6F/hnKKVgXfqKYu
bzjasQlFNuvojo0e/SLmHSHNufcgsQUY692uKC4xDJ3rmc8+w45NzOJ7Lby7lgKP
x571DX7SpdXVv9SFQ62NaFjg9aKK7nTSvCGjMdEgyaLE2AAHsBywUt8nAdBKWHaP
9H7ziz6wHJKKVwnNqpBqP6BnACJbrsHvChOMqyJhZQOuJ1pTvTHKwmE/HlbJg4Uy
NWAhgDwYLWnXpum8T/JvgSw6NMLLDRrQHiiQ9RJJqc6wTYSDDmYVt02ezUKs6a/z
xc+nrGo/AcQjr4DJu9TXElYKlbnsIWjG+9OpXu+tJsORsfS6cVREUGdqk2VjAukk
bf38gLyJM3WgHpZtlpBzuSJjbdHDJ+QbS8YGBrsSfq+8NiivMCF3X4yJzIomXTjf
qr2xLCv49tiPRsPD2BtVOenJEIZ2ToxZP3Fw/vv1R0vkVQ1X6akR97L+md1VEpFq
KcPCTMS7tnrAJKsTnINHxdGdxTk0I4TkptKIQWFdNYNtAaiGIuenb12QTQLSWWol
DDf2/R1xzRv1SHV/T1e1jYpmKoiwTwPHmQ9PTYBvdIouVLCW2rO+QpzHTN4TjmJI
Gq123WST7LMx0LGrkQ4Sky4Rm6b0yX7qVh/1/cu0EvXoo3YFjEMQtLCFLo5mWDeK
HJmB0/1hsZel3JiZKGjyRwokHiK6/Kw09kiGYEmxVqTPK8dx6JVk+HiVVli8ZUyl
fpv31cCTlT3JEizd54sBx4Czt8KjnVYa3qZN5VPTY2grd0MokoAEE/ASmD07veF+
aaoPHNSaZdIFfmjalEq2qqNujsLa0K2TLt7iqNYjwZoNtRf9s/QZrlZJL0jPxKun
OydXRniUs8re5FtjZwxxGf8uj0Qn8IMUosA3OaCRs6YjOYd3wJc+kStM97GTbzBF
mnWGZHREa8PeFJwNiqzj76tJMdDqRxpfPFglBEU75PcuWHkSZ0arfxVHqh62wnNd
emQLcnYl0MW+23VTRK5P8t9TLhCqplDVr4FCVQtj09AFLdEZ24cyJ0lNvvWhiZ59
TOtlx27QeUGFrFHTupKUvmZvO+oWE+RSbNdg2MlZ3Z6KoqCkJ3OYvzsDZVdjVY9Y
1u/1oYw/ygI2pdVTEyUFeLrzlQuqSMjmM5TagIklrtpJf3Jx3530R35IL/ILvjLx
CxUGRElWtnNxP5CYnKrWrxTjDv023lCoDBxyeW7rIF3v4NmNwVAXVFbbwnYZq6hC
uA0uYZZGBshePjR1VkNEHDLRqq94E2abecD2FnGwgUpOdjgJ8EAMiiK09SZi//VT
8F4J95mokQroFDigPOXr3lnd8ZszclgwCnnWl319N+TWx6WrWu2rDiPv1vUC+sPv
G5JINa2d+Pye06DpjEbcJiu0W4ZItLYfshKWhQAWOOsKecdwHyJumVq/EYGRcz1m
5JKpjMhx3Ys3NYBwpXtK7QpoVPbg9DAsJyfANKTi3lA0rAmb5KczuRyfSfrPvHJ7
wUIuushLhiZ30yMoOSgitooxBGtkODWeoHDmhzYTRNBteeUXRlJ/0sbJTABpi66d
eZHy4QPMdkmn0YNM5ACWsMR3YtyRwV+GouxmyMhESH1GzcE/7wUXkShUkhYZEqoh
5o9bpn3x6FbmLmlmFR+UoWnjZSRxCS8f3Vm0MRARnsdJm6s7G9Dvz3YbN9cZSacz
x10xJdZgucsWjsnjGKmeUczroSHp7b4+8/KwSpnYLhyvxkc76DUrdLYXTapihHPU
1n7oe1WyUTrL3H7bTxAFVuSwBWfKU3oeMEa+6ghDJWlBeiuSKbSWvHrsi5H7f1E3
9/JgjMhsrMbVqr8PAwxawP9VQnS/cwdeNy2d7ubf/DqcqXFruFJTA7rY2Y8TpjXT
p1J38isHY5lLTvG+UN/XxvAH73BMbFfBVRyGNz0Uy4F6DxUYuoWcgJI0Gy4EMrq5
TuuIxP781C4i30yLPn9X17DC+qEUFflYUvKeCx1KWaTzBNosJEXxcVoAm/TEUbEX
Wo7onHCZYCHvN5u8qX/Q9ZbJ2pcaaSiKo2lETEyx4U38zJ4LKSG5qrHo+skB00Rd
mz5RD9VjhqkUeDxNsBAQHyKBFkiKRZHEETa5bg+jGXQW72gham7igGo9lVfpD0kl
E0oQkppYDct/ClbOp6Gu9+2UUUmrdB2Qtj94Nwm+KUyMl03Y/qKkJ07dPf3a0CxZ
x8Ea3IUziv+IMTcGfK6Mo1OLKU/+B4sN50nDLAuerivoEaNzFOXxHseh2iRJZ++M
UCUFdPAie30GHy5ZUGx8rbdz/+tyCQ7wESRtgcIs8ygxOkk5Mcc817eqjNX9yCnu
7pI4pjngiGHzqNGXiMvp6xdEZr5i5ZNM3CdD0UT+l0qWcxlYxa9v6Wo55XNNd0l0
aB3VZRAWGi1T+qv/b7jur8mPCQBwz66WLaq9ssHLxCGTEftzwrMUkGJ0mw2wXY2a
eUnySQ35BtUpqkFA23AiKocgakasyd0Nm1N8Td0Y2uXB+VRPSpn3Jh1WcXq6DtIO
DUNS23T7vHsVnhkG8OSiYxuZ6fNrNyPZgo1M8ij18/WezC7YZnAvbQsjaUmVCXYV
pqwstovd8msNyG4QBnYe7xmAQ92l2oqaDH6vjbxIzxlY3JVnxXmnLGXo39pFfTLL
REMwT4Nr+GGW9BPmu0J7i+9/acNtf0HdIY1a5SVWyARgPXNlnU4n5wQJg3lcsV4Y
o7YEqViU4M4y0RmGOjPbEaRUGmTNt+OpACFAUysWKs7S0cJUlCzPGAI+H8BDrsRS
/C/xx/G1R/xZNOf/xbnQ8W8PipJRI3x/Fz211AxsfDmVHE+ZTObfTZoXN4315yKL
4yqoC2Vk+QKGbZ8BcSygM8U/NdyJsc1U838cjgTaRkc8vfDRDdXVXR0beLf7X116
LM3s8NJYQnDLfXJnJaI6x9ZQV94D1AlzziZz8qrsscfGo7nQf0CfSQ8nHP9ySP+g
Ef+qfv7vKYzjnEFIsBm/A13fO9KtIizDt47VYcP294gz2vJXWm5rweRz5dRuf0hx
+esUv+8xTUQRfvYaqNZ1rpNncgT1heXLKkUiBrDuLe73o7t2FiJViKLwbGJrVxhu
jPDziSvSfmlAOL/ruA5RLgILPoV2DUTlSG5qLBpYLx/6b3qTYS/w/dno+liFsG6b
YbETrbqHA2KAISwTFesL1IcpNQXZ5YWPpVW9UO5FuhH8yYwFfK/10iFyQNiA5Ge0
Kfkr+hSWajjKXGFHqoC7k5W8FksOJFxPYdZ5/eEV8fo8r0OGvNkOaXovFFwIfo7s
8y9J5vYLRnV9Q1xQ7DZgn8y2BO8GnBJc0qotEgpNFXv8KbABIdLwoQLbb6Wde4/t
1AwnPrABEbNqfdqPLrRC/JYYiI3BXWZyYGYA8hD8AW2FwRUG1eeYCkOMgI+t1l48
1wMEFgga2u4oEB060lOS5QGLQKXhIErlMYwoipT97kOmg+h3/HblSnCuM1SAYu6K
JSUsWmjgQtzV3TgG9IXbUgzQQ4OpxZrqiQTxrRTdC7GK+rZpPVGBGK9b9p4SD9Kw
NX+QpukMx3rtVaQru05yJRAp9L5JLnk4W6SucfxmwuvoW3ogTrksBW2841h782mz
nLRtDfF1/s5yUhU8mu2KIlGorMsfEP0ETKx+EHfRxnQyU3NTbfUr9zPgvmn0Tral
BUz7OXI+n6H3nR7J8gxvjwewln0jkUHGSUk62sRJrU0eaL9KumrmiBaYFRy6+pws
VDEERJFQoLQ9YFMnsN90kRePJY1w4xrzWiC80zNNXnylLcSOq9qo4J3h0+/sGqXd
5Soo28A4t7oOEXPS1bKDGoHkEBe+kGRlJxJsEaFNcrbjMvyaj0kiuPRd5RBXJ0G+
p4cp7Not5Snj0TWVTIDfD57Q0g14xxGYNv3THzLcnpEHJu1aV/LgBUJoXW6DGFPE
dcEyQK8QhBjnXo4s76VSleaBHdDCtQ+M/TXev5ZdfXruCYbBXbw+WGYwd3ZIPwTm
Kji5sqNfwL10L/pl24jkWmRL+wo5tyLNGVExhO4ohr9d0goH6hIDbbFXKuBZNMLE
CIsE8YbNv9PfT4eFzrfDu5G+qotFwj499efBaMpdXFn5NPuKE3QaBPPrXVl4vP8t
8xEIqYfgxSNVcw02edtdyqb1/zIZP40UClJeih60NPFoZIzaGTOyr2RCM/lYrbJY
Cjq2U01S27YvvzJGNbh/8UhYsbgNTgweMVFbZsKJ/Oa/0j5JC/RE+TfobKGob6Yu
LAkPXePN3LK64CzK9uGHYoIBrpI6QniR9O5NzwaGSNggRlr2AeZ0OuWP/qd4Fn+c
4FLt8S0EhdLagOyo7tfUk7D5RdoiXANm/Lb377nAqXSZ4ki2FAQuyGeYY0v2z2XJ
Or2aPNySqyQfefwfsZ7lZ+UA7CcLnyyFlyneS4H76Ts5cfgoftJzkuFNtfrj+WaI
eerkbZvoSRVIlOELqkDN8Z7JCg/DFAGZ25o2dtLJ1K2rgDpkefDfXOS9nUiYTeuy
sqZxQIbqs9FsTl54mb189E+zENGNOAttf9MDtz7PN/IrZg+3Vht6ki4MHK+Ce+oT
Ge4CSCYQkiX5bWNs0I8qu+VJ7qZ26DnPiH/HV2zGnioCzyMYwY6TBGfCF3s3yAqo
PzOM+VevPaTUVqYKVrbHcx1zFYKzdhktAUsaejnm5J1Voh4HgFVde5RFC4hUyxNF
CWduKTKXB76Ea8+j18zASHln3z+avGnIuccWatHWrNOazDmpM/mnHJQei3RuaA2j
OMm6hygH9MqDgCLF7ALNFpYsBDlICup6LYgI8F0siXtEUjrMcS5EyrODnkgIYSbD
X4d7v7SSyz4caMO0kkgR+egHxlkvJstiRrrttC05DBlBkl5HI+1nFWpq7blEUNpI
rIdpv4G/ko+MlwBCMMTK8Myt6AupOzdoOq9sX7eI2Xu2QLkXDw7AI9b5m8RvTBUG
UFvlJF5iV6jB94LXVLsg0XKkHhk6ENmHahnb9k2WI/bCK5/PfeGYD2/AZHuM/EhP
zCt7uXaY9oJ/B5jYLCWkqos2qpkP7Us1yjHnE/GsLIFBqIoT9B9CoCBkgTbaz+Vy
X/MexoGZhaYDwmNoKGOh5qQNu5j7nqOL03woAWZqGXMhMTevXHytSECtTanwSSkG
oZ5MN26jDsP8JBmet/PwX6wqDTkWKydMm5gDyFpC3Tc1l4opnK2RIMmAG2gSH1ID
kKGYzdpjVXxi+Wix2J2moWgBeEgWjRAV0CUcRf41m7nFL64Wuv4qxXi7KJtzxWYG
3zcZh8M30T8kVBJMB14YQ23SnEDEYp3qIOwZeXkf7yK15C7jARouhaI1M5qWYnAm
l+Xc88XWsX1KLhxoB6/3Gc2zVWSw0bmt0IfB4iJqu0Ciw7pZnwvTmzHbz+QFErhg
MIvYJVAtUrHHIvHcp/6jrX65au3EJnJP5kdIj1Lorg3dEsb/WuKuDYqMAS9KPx2+
Xjpo7Y1yM/ups70jfd6Pr/gN3MtaYALMF9mUS59hqwEw9AukzAmGMjfmiMFvsMHz
qybd0CMAtgDSYVovPsJqH3v27t5Q6Rp8ohj8dMjqTDB3tIa6XH8rEpFAx8O7TSww
NaLYNIhGzuua7UOD8obNpU1uXmtKo65CWntM7IO+MSxSg3rlkY2FrUCuEy/zYfFU
b4zo35RnZ0wd0UPAEbwiZoo1UK3qCeVt+7IgwS2LUnZv+I+gtllH7xBMHiLatd5W
B8Xckvtash+LWQGitkExBhR4OSb7CDvHCwqFKX6Tsl3+vj1EhnqR52LIdDIQWJPK
AOxaG6U6gfGHnYk5O/HdRXBJXsxSg7N+2rneZGtRQxBMOHx0MxbxaEhMerf+OJvt
ZFWNS4kqPHrpPiayDVZv7NLWFqPCM7HP0tXyqZgM9xGbf9FDmzESMNxL2TBdgQQ+
EPRoZeeyMDcp4ZXW5t90qGKds2YMemh1cZ+tdQBoVao8MYjf9agQlgKAt34kaNZe
kTKJ6lzL8iJ2cKJnBSCGyQvWEQzMZrN7fZIEXTO8LDOhJn6HAe/6K0X7xvvKwr/k
MDckvZeLH4Bg+0dEJqXkzAwhNpeoTanFItc2nIRFvZvC0JAca3Y02LiXaHqLYOo3
CFNBh+Fd392ERyPBuEROf3A8rl1+s0CBOfyGF1IrLPnn2DeQsCSzZ7Ub1GyMsHeT
KjXmpNKyiGe8ecmUtfTNNLWvl9LU5q21PEHDQ676bq6iwUy5tw6KJcV4L4CLHfxb
eoAkCmuCvccEhPZP9IHeCrC0mPSMiY1jH5L8DchDMkJmbVsw+ofgbwh+9McFYgFQ
Y3TCVg1lX0e5w25rBaNtMFAQqvMdDVE8+sbyCh4uShg27hj59vlJJUceU76CYlf2
93kE1YWOyaept8lGXP+qe0cu3RDuKT0JprrK35zaMdUbZDWQsryJG8jvVey8E04e
+kdFLEgOuu8U4w+L97H0aC4NFBgCh7R0/hdkifqKqsqyIDn1WfBcojq5u3S+SPsO
PyX0llUvYCeKzEQfwWMS8v4v4+i6V2FVXbjQqjvSzoi+naoGKmUJm/3rkgLVgvVh
VvDnzmo/lRAoILH3pOedIbbh5qiarGed1hcT3+KYro32pjrXDMrTnSN2Y7W5Olmd
xpJMk8qhCl/XF3neQoom2QQuQI1h4+Z4abKvBI1nD8vWH4QxIuU4gd1qqOKHY9We
HUvh4b1Imnk1P+7tI8kbJWx9vB5nOy+7lPNCNtJMPODscE+yR01N/uDtfGKkFORR
t/tiDirS8F/bdrO5oX42QmeLttZYjFLySdpgpyYxAtS5J3omb9pfgPL27duPiVee
S1lxz7mUqMOBfoaOk6uvtotYtYpMCS+yue9EvbNf4ltRXPkMnuxigVIK4EWfQxYr
dcZ3X1Hs64dIqSw1r9lFRtfCymf5DUOM29Ad0ZERSlpWreCcEXJ9U8yr4/UPDxth
YUG+5F3knyNaBl+jNTQiGg7tcxLuYr51Ti4KajvN5uyH03P+26fjVVLOydj4BT17
KPDAmulFtPpp0Dh6wzZ4bRj1IAKowHdfX5i+Bu7fa5EvGWTw03Lvu8490m+EmueG
yImjbX/XSgByoknlvOny+8Bwj1XoiLbEFu6LiWxhgUNg05IMq5vtEauEct27XL9n
Tq53DoRoHDAw4pj8/Z9uwb99a+VgPCowcferVwj3WLmf7rcvAa07kC6eOWqSu2ff
YWJHQY+THsexlnbC3pr5viAq7CTedQp08besRd5k1Y7zYuiPcH3OGtHdQKANqzPV
/KbMeEOrUiqFcgrxJy8wNM6GXWlAvFPpuyMvndbiMg5LqtJPfBSbNpQ8eyEALrkl
O6zsZ4EnmgjDeHEWj7qtUGX6WZvGW3MVj5CRCM0PFYnDJgDti9em78XHhP38JwJG
Pm5cT6LE9Vnbsz/xwmwkF/eK9bYNHygIyHks1U2hcp9gVp6rsH1kupaDvVJiryfz
29dAzrnrm1DpD512Ok6AJqnM9l7Yxu3wxhHdOrPfI1FeiBF87DeI4sgIorjxY46y
+D+o+W2jFq1Xr//ZHgAPS+WRFjc7HDt62/d8auddG+xfoxI3VQ4s+RRUiiHbZ0sK
7aPA0/ml/znhfRpXIfZR0OJMciFYU+TGHu/B5tuqzau1cFpJQCfE910xORPTnBN6
9o80eryVBJBsv9ch2OT6FjSeKPVWPdSaIRXMiktv+ew55l6VgYjDcEzDClhIY/d4
jXblRkhjOQFlkN66Uzq6KWHBssYetsjpkjmUvbEfSztOno8RyipZMamLQjjQomVL
h+ESuLMKGnj0fhT/doGHEEBnqOsUfIHmroERXvAjyNMfOXsviCWiUhmymuS4gkRH
s9k7YE4+JrSjRSUNbYFIAA9dClIrzjxrxUt0wIoQEHUUlAP1f+Eh4A/6OKi6+8rF
TAoTjpx9/dsPIBalyVIKVbz2ta+Jl3SSpalHVC+JOyltIH3EmXiFF0EbeptWtra+
iQOmUXUyuQG7OTn6qKnz6ean7K+swv6zNpzNCh5q2CIOYqkIvjPv41Ut17NfNQui
C8j1US6qzvUmr4gYLoTT3DF9Ine3rl9zymlAaJT88chGgQy6Vk8OYkM0Il2YTuzc
z5Y60cWmLtsMaounSMKVy6g6MrrjYxeCxGxN6tVUh5BipHvVbPNG/UNTvbs9wpRi
P/bxxLUBr75g0+EPOsMnnCeujQoTIzLslWanA6aLBzkCwbkToGvVKt1aZRTnnlUc
T7+ZJvPJ8iG4B/zoGou548ORGk9cSP80u5VuBvkFxrOz0+8TVIvRh0LYIwmDp2+F
E6qsrJbtpazJnZ1nLMVrRI4w4+WqEoR0kfaguv1ZLxElEZ9VKS9ooEHcuD8uPg1O
WZFuSarZJk66OYn2GHR9vsaMap8QvdZLBi1YTgqwoPD6MqH1fAcc6sTT15rgNvuy
t32I/z3bw0sFOwpeGWn5y3FIddEwlP7K5Jvyzmja5NAf4rIxb6ICUuRvqfd9yf3I
I+S0kULqs8cUyaFZKUkBlBwl9dIF6k//+lt4kcnneFj/zbsSZCz+4x5UvspfDtvU
MOceRO83Aa831EQ4Ks4R1sOXyCiOeo9tfFBgziZxJET55nPFUUQrYSLOJI8aqAEH
wGaCYK1K/gut8cr76UwHq4tGWpCRA5CDrIaKZ+Jk22pcsfiP6IW/jv20C2aTSM5B
hF+zYPJhv7dJYjSseLBpAB3rtmA0Z+GFg37UBmCxzmcFMCaSOtvC2HlOjuOywIxc
YDXir9N21GOtUldxf/aZacuMNi2LUj2CCaNDjMDxqZ+UDJErlrjlU1kN2Zan3KWt
Lxb/AtNVfKA+xHanbfRTcxB+q8QETxtinoDKhSQKs83r59CLXFJfhs8KzHgVuqFR
GorRjWPwcaiSQwROdNbS0wlnAzVNkYYZBwAicFTwdZSprgYeSx0CWt2dWSXsgIsQ
v54qraH4+yekKKOEVUylqkELl6Exp9jfABXZg3Dzn49lvlLqb6dKrhxjlcm5jXxc
sQDuOR64A7IYnqG7R+OtFtTK0RKArNqycrzB7wtrnBo5gKsSHU9BthBgXJoYC5Eu
4VdRi980U6nnj4JdEs69Kcz385wNJgBEs70cCQoOf9EjubMNB9zuOnqvvEUETIJq
GI9GtRMGBDvG8LadTpR04OZq7OD6udJXnHUPOVvycjFL8NfLU3pk20gYESvYN8KX
yRjbfZEYGUHLs+hJf0Scj0oR/60NFRHYRDJIrsqWAY8WAfYd2Vz7Mh8vIw6sr4lU
KNNIy8kgv5AC4T9QSG09fkyCSMtTwwa6envrtbA43t9/day62ggxsNqv3XBxABOO
CfZxJR6ptGUMHh9X7cjvbSTOgSQwCf9/UIz3LtpfStv+2Nw1umWrWE0K3k+OYrz/
bda0qO5U2ajvY/SXnkR/aIox253Bv1Bjx0vpp4yneU8z2F6Up+OxKJcbN/0usqxH
zus/JA4LWIYnzVQlOPqMT4E2z1dtIRVRUtFOT9jsw0KpEUWXeRUyFh70Us2iz61Z
Iucg+VgbPYXdpx96uGxA0DKghUT28bbecJ6MaMyInoM3WTY/BBJdlqVvlToZjWiH
Hh/JfyCbgzDuKv5xbR+awtjEVJ91iJpygGOU5l2+Tp+zFf1lB6d9RJ08BxjTqxNd
XCUCszmWCc5ASN+/DfVEoovnS5C/RrQZjWZwr+k4DOsVNXCnRH8LxUDdWGBXj83K
c3Dyk0g8NxBEbGbIpJ2tuGH4iYf7s0HHkZHr39s8oyNbzaaiNSPQuxFW54Rg9Xez
RCBaGHz9m3cnC6wuHEJJQ2G3i/AcYJCXM/OK25988sNqUd96GvkiE5/7qjJJBPmL
bJ/T/MgNWtTGOjjK1eyjl+iWyjl0CFPQxXc6nwX9+AWCNGC58Vp1hEI4Jnw6EhUp
tdszBK92R2HL9BnIEez25NyXCMYg2LEvVq3zKemcsvNNAwFY4BTxhAhwKcwviRkK
h8iIKaRLqWRLPc0Eji2uGIbmjuP0md7jCnGBhVfD2D106hhKHNcMiijkZSQQDkfW
v0UTNHGAFVPK/Yz2Bi4h5PIHv/uPW4mFNhLDBGOsu88rgGHJzmE2i1m6XkIT5eg1
L5fJrDR3mRmBgobO+hvaym1svrbAp5w/vNJOY2ZqRPPQXLyA3IGUn2hCYWeaT/yS
TTK7dznxtNLMbM3VU0q+dJBi+/ftd0zdDFHA+bXRiQimpleA/D9xgjFZ+KvfGX0d
IjbgqL+khh4TecgRdf555e8atIohVbYkzKjrAFb4UxMVtZHA7BlViJcPRdrO4LX5
kuBLA4vlN8w2qKjhtQYorruMTfNrJTMZSOAN9veqGjX3ZasktpHFqMNNqpe6SYIh
xz7StMkfu0xM9DUTYKOPl/E/QwaINQwFKf8HLEQa/BF4uwh7AL7igq9dXJvmhNXW
QIzzjpU63wxJAZ01mfu3auB/6uWTDAXUEdr8Pxg2eGXkzz80qXc9I8F8uH6MtiCr
F9bvnIKoRAgZQTsD1snW40sAM7EJoJoZ8JWAnYqW/aqMdKYYxba9uJDrWaJFKJVZ
P3/ixYSjshYn7MuPDgYZPV0dYIqI2ZNj4JtEGhA8+BK8Fh4PQ+pmjV5XozytdvgP
cJqKoWiPweVehZK4o/NOUNpNbeNPKjRjsGrfFaZJZLqYURM25+AYb7bnDIcoi56k
ovn6He+sKcj3i9xVKm/oGDkPyW4EPWwHiH3FRjLiDh/PXNAkmVdWknOo+d8Y0dzx
qwpQztFl2iUBc3XAyZtunx7YPbLiIJxBsfGFL90sylLqt43ngenSfuS+Kum5MOi6
FnUH2CCIj4xhblgh8dNxYv48I4BO6OZVqApjuZ+WZCcBKcBOawLnod0JJx1zgwzr
M9YqP1yDTGCBO0HWOQ7OOsAqvGJJX9vWrDQkwhxfh+fMKmNRCYq9UHPPHQevjzAA
0rhNjU/e6NV1AG/GrGqUHs7nD1l+Q8YfUx/p7KmyJFh2PhaQS9vfpPTUrlzblFmI
FmV5+ylWZPFRBRScpAJvCR7/dX6ldKfF2v7P81Rjy2V8sgraiI8b6ZIu87ehR8q5
7ee/7Qvn2d37ovhl4rg0iB20fgJKqo6ovKdHAbCkT0W1sQy4YcEqRRd2E4F7jmrR
ll/wBnyBjV59AoAQWSPwfPtC6SD2nh1NxdstLYzKWr2+p4YF94uIimC+GknxFb82
o6E6JQtDyejw32+z7mj5HP5NFcxMMTgvkJJdAtubdxlHMoxFOr3blDI//XBqAnxh
6ZAq62axg3mtEJb/eWl+3uphKDJSI/cyhHE02S+J/YyfQ1FMGPv4PJxTwrKljOCL
8jMk/rFtfvdNIpk83J10oUOcX3SbQWfc/B4FqNMjPM8nXSFgbA/pw/SppsKXU+2O
huuf/lQPVHaJLlQuB9Pkld4Qdq8ZHGaAsmBfe6+J1SVz2InIMvG3b6390bIg/zrV
DzRUjHVZmjJ/hQTC3GGbHqPWzyVUgRdMhn5g5Uy40lIOgVICuGeQCXNZGXtjcOpg
7NV9GCeIL9WpPeLhjrDuuNyYQ3nXco6jcjTAF4atr48683QJiQFSbLed+ji0biLX
JhbgvDC+q9bSukOBZK3WbS+ZvQuNNV/FuEjZBI1i2Jjsoc3i5t5UdMumkL9m4hFk
fsFByo62SQxiCxiqPoCgmgMCM1N6BrwZ76FhWWHHqteQGKuo56i+1ERvh0MSEYNc
PXD9XkIrThDp+mbMuCzpRNfxJda62OkzayoWgccZx4JqG8MY9RpCBto6A2ZeSCnF
Pju2D6+XYIpnhZgO9oDpmG6hje/Aut8im4YcpVYOSV03tzWiY0yMlojQC6ZkJwDr
FUn0CJeZwWVQfVmDjeWhJfOOmfara4Q9N2VLhZ0yWRNDpPQDaJKVZpW1CQvMhJZj
Uy2IIw8BSZlczFx/R16BY5aa0UIiMQMvECYqVLB6P1HncwjVsFQbvFfE5JoJacDF
erT8W+9VyRWBh8Ii8P4iUcmtW9QjBbZpRnzIaykN8Zxad3lPvA0zd55dX50Rafu5
7c3mAK3dURZPJz/BTcdk5QTOFEujcW57j/5kWN+MbcfA7a82R0RapipOdgXKqBFL
JsOeLCkhF0PGQbPtH6kdMMChVwLgDBaetTR/YAncOt2qbPgJk27kPx6oiuRineEO
3gpUOHr7PIU5xOss6hfZ3xc7S9aa0rHL7GP20/mbqr52jZ256kSyKahghLbr2G3r
F+/G0v3JonFo88iq7iee7BWojFPLTbdrg7GBEnTacmXhhHjbk42rkLi9VAQGUaZs
g6UnWXgh+96xgdKGDx0Mph7NdmHV8F4D7kV/HzKZsXvBBLeurjoP3bKE0OauAIC+
sQpkwxGsJVhNf/pCEtu6wHzzeCMxO9a7v0U7AwwjGHlalfqXjLgepNpp7QBpJzJv
WBTKCC93G+DjJYm97IffUxryFQUEPJTyJ5eR6A1t/lPVbfnBHM6eDGmH/laqxUW2
mIuZ8tWL5uq9FUWWyGeb41WhVV5KJyXHPksp3dYiEyvqtf/GnEFkMFmD3yA7kMw7
Zz3KOtDjZ0kc7nX3yaM3c1q693O3E++TvBIH6ep5+ELSdQRwe9sBj+AWIyBI1+7X
dz5r8+k4b6HYlnz3UZ2+XA5W1X3ILULmsvNsHTsucf3WGFrgMytOwcDuGhZOzMwm
3pUViuo9A5DlKip2J45sg23V054k5FqsvOAtm6GiGHNuywdAhlJ05Qo3VJgsB5cg
aMu8PqkcUI5UguliKxyoCG9hcO/XbE31BTX1VBphKsJ9FSoC+G0fGkNjdPXlA9Ig
e+aZjUl8v8BjgjzmeQ2ynxHHFj3jcb0OzpSOGqk7Gqwj0NKwazJBTv7+/hFUPZdj
rcK7RlLbcVlLSfqBZjuIfrSEqK2t6lyzRFb/IOdb7+3oJPCqbaQ6LAKYBz8iZTfO
GAzWcRTZuSpsVqftxopTUfYrBREASGlZWCazkUhDr/65p+yPan0H8Eo0UgmqR+WC
18tJ2P6bEcs4NnqL4oNrE83k3yDxM7YOK+AdSAaiE2V+BbiJdUulcj/y54r8thy5
LZZ9K09rUMpBe/1XOfV3TcYR/hFkzWbnXgTcX5Bw58OYfPX39mHwdQVwDXW0QM1K
Tzibqc7nc1ncD4OpaUDy4sXCZS8UpmkK0p1/tCj1o3fNHlus1bh4ncdhk/Mb+jji
MhFV47A/oud7B/5plvWrrpSU+KERgSuaB9NHbiBViPLWzml2P4Ih0R5WUTvqfSy5
6li1v1BiRxAccDz2vrhfW8tqS35J1xLr2c2ZquCZPAEhaND2haxdkR/unWF6Jl5v
NYJiqJu57xo9+EgDTtSdHYCRfNOu1Ztmx2SRk6hUbSyY1JPoeZwPRLKHd+yONssO
3qq1QUHNI6u7aRnnySRcRpxJwtk6Noac8rcxwvybaS7Jax4dnSooSiXJi7J3PGFC
wxPJ3OFjEbmMNfuZd2+ps6gYqmZqEyYHmQEwW+7u6MN/5hzzoqU72GCn4Rkh8XCm
1dr0MRyWqQ6JWicUt/cozZrWhH+zJmkzOH2w79NOQgCiXW3BWQXBNSaZuQHwwSYY
hQ7766lZF6xzRArUgseOcoseQyj+FFI8sBLgBqxZNI9q31CskOwAfefG1nPvaafa
45Iu/E1xySyMk6zuGcc5fNfFDXLbCsCq2ZIWuCUEDWU/55mnUDYsNsQG1TOchrN6
/m0BuW6oFybHScLmf8GGWVJyyq04Jl5z8GjGvDM2Rs6LPCmuu80qoXJaIzjNYrWU
cToRKRJj5YtR2/2O6aKO1eS4Rb/TXwdBLeezUxVdvcMy+kfldvIhXK9YUxd9XMNt
FfbR79cbyJBA8iFamzcEy1swlPcD7FGHYJNkX+QX4RCGhlYyQqbLtTtOaSVSThrx
DqJKIM8Ncit1l40Qf25VsDmbBOKf8kSBI5fSTrpud/h7bZhC+ykN7zUwaq+A9+sv
7CcBYQqnCJWj0LORUnluGKlJpjHIAAZFEBM5Le2ngMf9ytPA/g8peNZ8gdo/47Dw
tjLOVzRXkGavAyICbuncPdVSNmzjvUzsjnmJkuuzu5kXQCNcW2AYZDaQjregGsHV
j3uQVde6y70ZX6Vmc6Xdb70qlOmxs/ubYO5JQPZWz8BfS9GUF0mJWd7ShFl93EuX
L3mThrSubck4UmpOHjp8KHrOdQRlVIKILwfSvZnMrPCM2fgpW9VNXi/3uK8DthHA
MTTb/RER1inVez8CrF8UVMJC3z1FPoQvGxYoFwKOGqpt5aOXgHbtIqJEhEnnRoJ9
66egd7bipGCUAVts0U42UnJmm4DrvikRjUeBJLVQw2LKBJb3H5/dsexCkuwYvMuJ
AcG965KHeOAr3axyGF3jYlCiM4i3l2o8HHJPf2F8gPH3Q/hMstnZ0l8TzFGbYzNj
ykFBARx+gAOiUVtOWNFAR5vRGMbsUO9DNWz7RDY2uuYIEulPRlkIeUNiHB0pujTJ
pXog5pK04XHjONp6cB3GWs4smzXHyIOz5wEjmR7oHCr6T+kAD0Wbqlbn5bIRG2Tm
YIAn8EnExgH+wMLjL8axKlqWrpbnfQUTXYLIa+GIV9Fa+VuZ8gQJdiiBZ4ya7Dip
7a1cdWDroCN27mmPyaymroP4yO3Ivbri0t3OVTGvU5CA7QSnt3nc6EeWM4VCWMxI
8ryEBH07ChT9xbO5ES9gglz6FrO1tuNk0IRpV16tn8maZN/R7fAJ8ucKCupc8rF3
M/gx7vDyt0LzrQbJFuRKS3IWpFL5RjkKxSsv/5Kitvu6+MKI3irGrtJF8cgG5fGg
fhVjYHdmSt0S5vmwEuTvwuTjXCxIdEoT4f9hXSYfpaREyEX8IuX3au5zGdr6l3OW
hGDnjoZWVYjU4RhCqBUVrcMwJTFS9iKcXgy7EaCWD4rPybx2BfW57GSWDdBrTspu
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:26 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pWDcESP+XitMIs2J4wPr1ymN+rvupLASfMV0VEYWRtxTPu8864J4m2Vj5X+bgkKC
nQ1XzbkwKIhxugdS/cmelzHkAvtfgYf2r3nZ55VaBOUTxqbMtr2P2y/1qN9BU1iI
Lk4q/R8pEd95nd4UaJ4QRKeZ6y8XwgyQdX26zYqYTgQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1632)
LMGg+gU//jFjcFVgDvz4Z9cBWbbWrLSsRMbccPn0b4JflBHDXIi6EWMlDeoFkhlT
uMOckTlDWwqJW5Twgqh0CGzXuGRNnwPHV7DiZfcxxaDuTfjGnI5LU1gJzEVCCGRm
C9cO6MrepLIB437GErZl4YWVoQxNsyBK9066pI8rhAMtVS5ipCO2uiNk2PI3R5bn
EyuCXEgkMC4+UUJ7DM8PhyIx3BL4OvdxFDCN8lkVavkwM6wF0IW66nGU+EOc35ie
Um2CqHpOEbDxwOVEJcicQ6cpMmDOdZ3zdNZWbgwuOJ1xCG5InE8yG6rbXA439FOs
YkeLxKVO0jfy4gayqHUpnIs+1MGvAPMUQe0GcRmDIQR/T+dsTuEwDDHgJcthvm8t
cby3SBVvHymXguZDLQk29gpzvrxHiSspLVduPFNQ0RAxWyPvCfyEAnRIUdEdXQ5K
Ay4YUjPm7WZLIeYV/tT9dGpjO1l4fZId2G7DLio/Gx1/Aot25BqjjHlfw8uLRMEH
S+aeDZk8uxShrjeSheAzI9qSsgANzaeOGEvOy/3eK5sHX7K37JlwYdD82mdV+nAQ
GAl0djAaeUyfW9j0NyQ2iZXz1tG7K1jCiSkrINVjxW4LG6nO6QvUwJD9zhR4yUc3
5RtKTujRfk8vlojzUVFA6Kv/8NxqELW3rQ4pQ/Dp5kfuwfym9+gZ0qNByhd/is/u
xTMHE4F/6Xy0UGq3gM4sBTsw/dYu0rvRFc1XyxOT4WEGw5ZsFr2xt5LhVCPdHgbJ
VSgO7zIiATQFnZCgZTDhk5XqqHulOVhnPcMIe0tjirQhSJEaGyf+4LO4brZzvO/t
HJLfOlGeFGaaScg/vtf6t6OxuoevIWRcp3lauIr4UABmJ4AgaQhWD5kT8bp4fnYz
jGmoTPAJMkBUjYbGcdAI5A59XZ3vhfTlSq/Wb8ve9ln/Fd6324H352S11Hz+X15c
szHjIki9kKOff86PlTzQSHI8WObBTgRUaeka0q/gacaHsBpm7pvQkqXCVAMwWD1I
NO4/w9KauUP3EY/y2+opb8bM+nuU9iOwEF8o0u8EH3NGQkkYr703zMD9htjbm1/I
OAgNVI94RWHKge0SNplSK4oWwvQdmNZ6ivqqPmU+uEnz/hmpEvGUZOtUmVU4pgWS
1iFJ3r5wTTt++5pkFTmAxUkw+hS3SsAFDDl4mAYv8gzfljTuk+wrC3kP03a/zxFY
fYlPPbFgmwx/vShSz/Qh3O2zjrTAizswKNy/ScF+WPpgESbRkGCDXG58TkxG7aaq
TJCmviEVxbUmmC+jpus9u0SOJJX7ol9l1Z1/UFfsPKSQM/4Xd96JjEDgXWDb8oZV
yoHXAMAqNRCCDwW7W2tGKnCHZ/pZpSCHm+CFkGpr/vt0l32QTP/ux/2Df3MtWSFC
GNIzva6sk0HIwQwVOzqG1Vz7scL4Xs6ixlKZWThbany4dnqGYdi78YwuSCgAgHhq
FGSwutwMWcaY42F3fqoQH8MJFtUuazgAKD79ufJpfbOrv/MMRyV5iXYPwXPUdZqk
FeePZw3MthJ296lmNIWLPedlH3dsMv0KcBrVwZ3Lv551+fNSuf6gpoUzu9mROubV
UOymObWGvafkBmIOX+GCi5r3+ZKat7IaZ98WT8TABfbK3X74gu80im8hT0Fyb9GH
PbwRLqamt/XdVXnwMjhIiEzZSkMg4Tbx6gp+teucUHJQaXpqltqMQcAymJTqaClU
LYSurVJHP/zZwyq+d+hN22U37YSBh8hN5TfCzmWN/2ZVtk9J893F4m7kkJq2WkWr
DexKAy92pC8oCXyvcH+4KMBysFGurNBnm4BmjznoPAV9QSu0b5rSHzIpw5LSNydw
d2sA/LObfpac28GggRxGIgIUapm11IHC5rFtmMbigUEdKYc3GQKCW8RSf6zIb0Rq
bS0oDwgLm5oqEWSKTYYSu+2HQz9VrQ+74Ws+TvkiRwSSCTutw72XR0DJdK7XqfF1
d5zFyQtmVRwpdiyFsg+UNMEtRNjrxs7GderBoMwCIFCjJTdddHASN+PVFFvR4Zto
qZDz8Da2Bsw5J2U21JI+KNt7c0NxEJoQTyL7p0VXrzOYvuXQ4eNguFBqkwo+E5DI
v5hNBZekse/srrKx6h43/qZGZAZiKrFLW9IMSZnCOO+oxleOW7BN7Bjz4ijQilJY
`pragma protect end_protected

// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
l//zd5fpj7ZzICItb2sWNTtyqJCRikKIeL+6gzeuzpljGx/Be8Vtg5U9XSbyCwtjVST076L7PFZ5
ErDzgHtN81pwT7POu11zvtpC4yXLLutIXwpOyYkSiTdVOHfPH+z7L8SlYCCfRlpPx53SYTuSXEMg
k1vvHSjOny9KfQppSQhcquuYque7JlkJWzxFOD5iv2FC3dYIah4YyPwyBAHQ8hX0ZHP+7XqwveFb
xL/JGWdacCftDnI7wZIUfiUcrQH/81374utooj9VbBLVNhuFQzi0edwuLOfY4OxNv3i9b0aMwuOO
RsRpKDPsnBb68bNv4BCHKmyLHIp3SaQaWQsspw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
qoxfTUZhyrfBiE3smNSJ6vfrIX4PIXk5kIWng5ewJAgFUBmfu/CebaJN4G9myCeUQRWYi5VqQCrB
BfO2EQHg0NYJh7VNIfIGZ7/XE8/buAtmT8M3Cryb7XUrzt8dhslseLK1cabm8W3Vi6XJ7fG1x5SP
+FcsVuM29/0bwr8ddPbss1xGozIu4MbNXBe+p9EFUX3+XGhTqR0GeBU/XnROmNaB7N2T00MgSW0v
Avs3w4xbZPVUpkkUg56vYaOSIrKvh1NfVWrk/TPeV4cj09Crz3ejMVnT+PpimeBMrJm769KzCvL1
8c7j9sphKOMIvDlbHPFfO00rzuC+b45nQdp+Am6uzWHmLZ4WMtX91rll+3d6AJ76xBpywrY+TSBB
0UcOorF/6ZHRLmnIxg053IQIAqbsdFxaWNox7qrA+qBJIBlCHZEldb7fnQlc4T9wrXQv+rwCJfZe
Om3v5RDXuzDx9nE1cMp6Nxdv7X3PoFpi5izlVsRihXa/tuPg5fopcMwC8Pmyp/iuHskZ6Fb2vXxG
N4kB3mXyaaD6w9edz7P7XVIWCgpqCfPr6tKCjvfbbqNbOClfxMwrTtjk/36T5eLYmMrz46pJXTEU
r9Un/evBgbADUt2IKbNk557EdGBhR++H9lGEvuwv++v9ytSNBYvHHUhVek2M4VFqeoMBAncEjO1k
ASsFV4rKW/IhNF0J6MHsYsDySbhDGezNI5/k54cBMOnA21OoJzh01Tz2ONf2lnYl/DDdjq0IBOJc
NOra69pd15aocs58WdQi8Cs2NwHNpFvphJkB1RE1rviIKPq8pc4/fYM25zgcqb/ODDc8FiGE0pqi
NoUBkjfJcAak5trpRWeDhiO9anvRGijydl+FTUtLsqLCKaGBJGbyj63K4LBMAZq9GMB4u7KHruWS
vj1rOedt//mh2hFzWmLI8mjFyCeWjTYkLQzZnn4c1GqYkHEI56wSaL5ZOOmghAqR8bgj5/IpqukE
qWoBh285K8jDR7dmpPl6QirZncKallE0ef/wD+mwdQEMRM+2JgMZYtYL4rK30NHG2/cFrllNj/YK
n2hMEUZ6OKFHfXLjtABSFqjZyTiUO4xmMgk+cpMCWNAYYIN9i9LS0tdsSmdjt3HMTiATgFkFhJqU
ua5OMianjnFew7MLW2uCNORsf40YByJZ5tkL6vryYkrhx5/0YB0Jwk5x2VJfGCYXOlxo4cbsLPFz
8MMvJlO+tmSIN4lGIkeHnTX+coOBbFwyPWtiGrYFFsxi1v9sT6PnIqkVvnld8PItQp2+SpAtKRwH
kbHJa1vjg015aza2UgyZ/uLY0+NnJ6dKDEN+vdnrk0ZcvPmaH2lc/0rbujH9/9POt7SfqFYjfkNV
B8K1Z0PrtDuVTGobveqddPnkgH5felvNdTRPPwPnpS/YmYIZDASmylW6zJRlj8y0BNtHau4sViJx
YVwpS668KtRZFzfGXHS4fhgD2ViafcZexzhHx5+fvWrN+7jsMqgcZYtd8tfaFFVD3aIl635UFc44
2ko+EHG6eBoMcGg2y0IegrZSgk0dSwdE08ZNHnNvhP352Q+kdeaH3LEyqrmW2fLuOIdzNP3DFJaX
U3fJxJGpo2aV4v6oIho/hsxJ0iRz4nGvpoCnt46JQhYBVhjNEHPkjZj92JVIblQigT3l03DJvWDa
TWBzs4RuRixqp9Qq6JGdt1Zd+9F3Jnoyrqs00tROlagZ3TL3ufnpfdqn/P7QJlnqzywHIZuHyxXh
D/7w9IdftdaCtb4yNmPnzGMObSPMQhQcFfcT0rM2ieyQG0epOk8zALh10qZOlt29VMy9/n8xMy4z
DywijkimfSBCGzTnMN1Qr4K6Gkkv3/RARQQa+lXUcCY7/X2n8xc2N8i1P8YmJWxIRerFf/zdkvPv
sn1aieHET4/YgdvnIpy40OsU3unmjUs+pfzzeQYey4VUfayuT2OQ1B/8iktyyRJPd0U+RQZDPbO4
ajVeji/0LTsMAzrejkeKT7IUf8CI4o6ikgRrJdiwCiosozFUsWNnfn+VCMEXvGupyqVQ4OqLLUB4
kFvJAyBHF6Q4NyqFWobuwtl4OIgbTP/e/w+vuKRjIEYGxnc5tX7zo5ohHeWQJrKpYcxibFNIFkU4
HQTidz2lfhOtoqGCI7CXzB5sGtR/putawvHaDORl57XdND2LAy3pTJgvtB5wa3AVg6Dgisl7wVfM
J+eBQvUfmigQ5dRmi49ux3FPlLvt773xQVtLfLsFrnjxCUHAuTa+W3ADbpmhjkhXHCpl3XthlsLF
Gh/xheLqrt7W2hXnCaiMLXateVuFIDj3s/nZJn2xHm553QXtVXPguthJYQLuYtl8Q4U6I0MWVc5M
NjSI5wRI3ITWzWSS+Rhauk/5fm1lealbhtShzqSOQSCUED2lIvdGJlHerzdKBtWlAE9SwXhmaueq
9XYPVgufR+o3+x1MZjVkde6s6aMRf9bulFKUQJ719EZgTbFCjdpObCLEBzZ9GJI3YF3zxkum74E6
dYJivE2Rg89Sy9dzcNCLVVniVrtrfi/LMPdA8OUNjtPm4BrhSX4d5eZdiR12VbWxKd1w6Ft+RB/q
9ZOKyd/N0Y2KlrXft5euvSyudH9EvbpFikzMz6zVAxw8KSB8CBiJtg60XIt34sfMmwZxklSty2FD
84rMbyiLliaTlBFhw3F7Z/sqM5bh0geawYqCBbicIttvwfdDnyuE6x5wrmqXKxYepH2Mce3+nZrY
lBX/iIa4aZNwG52llhesvy2Wy9xKskzulnAhl8XLJLJVdvwVEgReWqjrljtv3EAOQRbAeUWWdq5C
NgrlY0/8knQCUjApBVdOa/RwuIvj5lkmJYm37MCsacnbJ1vJJT3urv6KlHxQYIR2sZi1Yras6Q+6
MabwsipCe00R6bM/0bTY2UV65slHwvE5gZ5FuBBSHBfLhuwDwkOk15IrZqE0xRALA00Vl+G3hUdp
4VglgVIiFFX8bj1PRIu9AeEZI8coWaoQgKOXpcIEpyGvBUTfQRz6tN9CewXw6hIsQ4HfbcmKsf/r
z1clqhumgX0dNsc3EvXkIykWIgncaBjweDGmQQ5ZZIk/cNAoDqJuWSVeNi/85Ug4OjjPJIgZZEZV
Mad/u/AEzb5JGmd/Z0JsgiQmnu8UYWDMgdvbMTQC606QsDSC9hfDZ6ybPlVchyFoI5zD3gbni3zE
QWL2FL0vbfQIC2sWOQTCvgb+kQMRocryz5+xW6+7lGe8GvQ5MNXDf5C53lWvd7NUMkqHClI7R+kV
TUzbww6Qp92ljeKQqp6WVu29pLqviYbvRqllbhdb3t7cJxTrqc+vfl/SSaXf5QOSSBAHN+DtHMbv
+f4KUlN8+fGbOVmxNBV1V2xRcgdJxBwUYRUly70+KGWKEhgqvO3MLzVgk+5+lIgFpoLFj4H6mGj6
0DY8GmrRH/a3kurdoRvJDxV5QnScwN4RK5KGHQ0qj4lWhlFDUgvZtP6O8wx4DQw77vzG0r2zUpR0
mSN0SukldE8Ci8wvnydP9HuBEundoV1qwzbHtg1sT1/rgsCLARn39OUZaTPq5UiJg7Ns6rlaJiHf
c10k9fCEKfRrrsAdoNonh9mFZXfYrctAeqsPCAlkAoZkWE0/a+NaaxtfZwznttu7vdyT5XFKOvcV
tH9zTZ/oCE7I1p0vr/lX/VASnfokfamFH/rMU/qIoYnrsDJgrb0vFk6WYYuddnufo/X5wqFxSg2e
b/fBLiGcEF7oDtJaLygz0h/IiYWn0YOTPFs4yZx5WW6eGT6EjVLTsBJQeswStU+Waa8TtNZRB6cm
pPaUARyTauJloXCOgJKBUcEhYMscwdiXPMTIcoJpLlDA6AoSAEpoPbMqhzLyvK/LVArt0oK1RIP7
II5IZyeee16Xo3xAICTSA8vvuKDi/gIknu9WBNm1lsxwXv2wri1mMO3RShQ8ca+eZUaMEvAVqfyd
X4Dg0I5ankB1IUATpsSxznzlaDWtbWDVDnq/kn+IjCgrhQeRhNTjSIikFdgIK2yd0Pe4Fwo8+/Ec
q+e1Th8hxbPxrncE+y57zKpfP1qrpK5gF+EtTy9YiQ1K3mhbOPq7OF1pY5QpVc0QmjlX4V42cgKq
1BOsy4chFLk2IcpSICzR0z89WbsS4tVp+WR+7LHLvdvhqi+7wJ5KQmpN6m14vn7PLl9RVnoTGHWb
xyJbjMO9w2kuddiC2N1ofjkCOVqJfsHwW/YxH3KOi24PGSVl7i9KnsXvkuSWpBCdoyFiFITZHRQw
XRdRIklQMclZZPJKwODBO2OwjDmDLzbSfmk8HaJE7FksTQh3fWQcucKQcsdQbljzroQK+iowstd8
75PYrWTXjtKZw1Y0yBXVZa6IBMGtctX+oLQtNEqkkarKoCB68tMTRfFO8uwCXp4n3OKosebDzJnL
6+TS9Bgn8Oahw9dSsXjoD6s7fs/lOyxghy82ZWsXvFE3F9pvd0RJD9tDRr8/S+1W4o27/xYWMz+y
qZNts/fzjGDuEShBfsPQVN1tUvsfx/4DyxU6jY2UOFA026AHH4kXnagawaUpV0IQUU030JwB+8iC
CxRyZSmsD7anelvfgawZuXItGCbBU/k6+6Rlya2csv9ZG5nX/ETfqTXIAtHEIQ7RSzZ89DbPbXER
ZQZMvCnnuuU9DMxgKBzYYlw71eSJZrvDYIdyR8fOjrPtJlyLNt/Zlj2IWWG69Dd0xwXs+maN+rrf
VJxfG6E9UX8qHEDZJB6mZeNpAW2xObGhD3Lse0lS/EbzCCKx/Zoc363nmrnR2OAaK4Hl5jrNGD+g
VgnRAsKSBnojDqxqKEa+dNXpJiqg6Jza7+JilRd5zkVLh+RYqzJe+SXmsiR5Rn2M9VHVx5vhql2w
+f68JnEOerpPQMeNan7ktcpkPxbTjXX/SEGCPZw2lMLnLslhjzRbB+xG6bLOOmrO3hX4wLD13gQs
N6ZXzRO/4Aqj7tAvgKG/M3LzHMJnG0EcoNegXfeaJhzBqZSqI6t4LPEIa/ER0NvsSrBucnLILl5S
YkZhtCcQ//n+8them8pn98iHe7MxnM5wrYaGAUDYeVRPtCCoXeCAmEsaZAqBoplXr+YVkE7MJoUU
gTMwKRKHSjNqY961uVasJ6cjX0WkRXQboyreGqdERTIt5GLpyMk35NyTFtKVDnOHWgD2S2Onri6/
Okwp5HFL7Hkui503oX+/93hI/xMHwpMalA13jdRsqDtLKtVGLxyy20j8DgtVHJc1WQ2JfqwzCF/k
5XWJAoeKRO+VmISntAhjY0G2JPJVl8zgxKwyHJNXZ5EwTK+lMW4I4k1ppC4P6ouJjHHMBrKIfdes
CR53MqNtzTbg0hrg1O1Lxc8kEh6fVGr5xHtsG6Rb08L5qmGSC71Li63HnupqC7SX1j9tolpIUjy7
yzLffJEr3KluLEC1ig4aXdFhDkXjrT6z67p5SWvNeoYiC4aJTobRSH2j2KXEkaswu1hbiByK5dLv
QhKPCKzttf07YScPzaB8QaUbmxa/d45YUneT6znf3b/gsbpOJDuKhKaWrr1ZsXRBSkmmQn4iWU48
aBso5hqSkeMqe8rTQzIXdtvvwj+phoB6H/zYCH6m6C6pAS8FzSQghblfVMPyjskoV0MAZqFXHgg7
u08YnN/KUwPmkmUk8pdZ2wt4wWmdJlkKejGtnFfz31vF/WQOz4wX3iGOGcOj9HA54JoN7krbk8iF
MUMsMdsvqq8M61Aexd17YqZjFuO5ppufXZnjVglIfqAw1S4cl14uvg6Fv9l76x8ZqiMm1o+YNbyD
8fqyucV9w+KD7hI5Ci+4tP8G1lLfHngRywZZkvaLTuiFsGIF0XYzxOGn9VMNsOqrX3QXXgaYCdhR
ply2xqPUlCVUGC3YSq2rD34VkyZQLdEKbmEo0BP+Rv+2cyOab4+x3kInYHMz4icyXIf8qEJl1V6b
EkfAdksXsQzH6ySEB3+uSb4Dlk5FzvbHl8+68wK/FLZdc4OdT+8sNjbfg6JXVitS6qqb2a8q1SCF
NhXoBN9cfdxyax1lOPWGj9WQ096aztYW34k1PpaXszf2IOS0L1jKpfS4wT/bQGNrqVk6fmvxuXiy
HG0keZOJs7VKpUd9hJ5GCPoBqLWIhKSz4mzZrR3/Mtq7w9uRfNkMGy30Ya5VPlS1+90apQwNWssF
tijvW4VGfE/6kArMb93wDcKXNrZ47BV3VLhPyncrtkhJNWhalYiOF0G0jL2QAbZv4r2XOgWQBZt/
kLdiIpy+MZO66kJLQXjUb+t+9XkD4T5JevQ/H5dpZbJW/0dx0MA7l++FLOU3RS3PzD1bRdYe5xNX
nWKABqvfMScSchRp5Nz+otxvjk8Q7/3UlHpUtaCdnQardLw3Wr/fi/O8nKx5jhJGcLMfAJlvtwTt
68emxrQUiPiBs/0e0lRGC78ond/Vxt/Gvganc8tU73q1t9ai2lu/9QXqtenBwzICiRiZY4e0KDoE
Msvo68RzICXUc/VESozchVXIhvQ/ZIY71doLTfeh1yknYklbC0o/SADOEGhiuTq5rtgHx9FjpCwg
Q1ghcbnbSZv/G/+56KSovdwbHmqywHGBJJv/n1xO6oO8OMc19eld1T88H/DP7g8wRWlefoIhc2Um
AvMEXlgfa+6N2SQD/SyGwQksYs7kH4McikM0AjFhphQnk5pZ557oHSzFkufTP7GDQ898QIfzPuI1
8oJbi9QxMfb7aSUpPd2YpIAksCxex4fTp6wAUNm1gWKFzayWqRE50RftQ7TH8hgCbcqS+VgUrwbM
nKgqQnlSjEiQmCabe16jD9zgdgrgwVvtSdH+c2pOVtPMgDixs8erJ5Su4YsWFNgG+l2/l5jE+U0G
8fAnJkqwPEQlmFztPyoy7G9+4Ng+Ok83RT5vk4nFNj/0d3BtxD0HdIbaV31eX2Mm9Jz4OAfL3Mfu
1uyFk92NTSe+o+EGR+LUl4Nnbp08S7RBEShj7KLMqqqNc7WNzGT54kFriGCOi3nHxNwdlDuWqnHt
88jlpgB0mEPJxL9C4OPtAlBMk7BLkSdVdkBqLP51mIepvmcIQ2IaVJAb//QPjIiMQfiqqLUhUnv1
LE2df2UXr7N+2X40wyETJ1mhQ4DFlix8Vsdsk7B8jlUq0aPqce+UgDA7aJ0qVeUZesS+2/+BzDef
IUDZyOUpXAuwqaXqanr2WKWzLSCQyqer3TOPQJQhQ9tN8Gxx3WQRStJVX1b2kjYXqr2ZOKuCdckj
GsBw5pBZx3Y0yAR9ZJubKqbzO8cHFu4hsczmn0mMk0TB6xjXysGDsSIHxj0LTrhWBLAYI8pCBjac
J1n7XODSdaW0E8vpjzbXPB6uvoi0HVV36zef4b2JWXIOEe0MgSqfMBW0pksZ5Qz0RipXY1Dmp/ai
/mvZtigmFYJJYO+h81NN1iGa0JzWLmAmfDd8FlKTnJBAdbXEJDBo7k7rYfZ1ObyeUJCqxU2Oj28V
+MFqQF40uhXqV1gv3VtFEytxzZzJFYieAuhiWvkriJQS4NgR3G41Se77MvYiW0MSUTlBE1BS4MH0
hSu5+rKWMQ+7T1hYmoauM92H0fG0w3E832Dg05eyzZmTn9gzFz0T4phNngcB8PUIwRA3aSypxyux
kE0TGomQd8/PyaU/SGgJrR0YrIkf+psUFbXDolaXEw/WgBA8tsPV4O7xYpPc4hopL/SKtjyDznEb
zs35e3bZoPidlUJ62b1SGFlbl9j9R0Xe45GOtd+J46+sGzdBtN68vc/GtKu9Nh/xwy4TuC8ihXUB
K3yXDA9e331wuhbcCxjxEgRRWnacjMZmqtsZNEuWvfPeDWdvkGPbSi2E7itfKYH+ShrDpLa9r0ba
InEgnffAPRvesmrIJPUO+OsSaJaI8tbuT6xvU80BdtTAcmjFl9P9I9ZZgrERRlEYjWWlRRyYcK+R
+A+JNIiyeqEpx64utEnO6AmSOIbI+bwfDJXx5zE9IunPII2eN9k/NUsRCOF6mpfz3jImxOnDl75Q
70KZRxRr2qlUjN8UzX/lArgcqLqeuVH55HOnqLl7WrNKXQueYBtaKGaNMt9sLSKb5t1wKjF6aR64
c2lMkXYx4tBhWmzqf5yQ2VCJ8/ai73tsDFkZEWBLUk4zR3/ihGQenugzSnyk4yJvKFUXIy3LWGYO
3LHgBPOOD90ZFwbAzXijHg0d2AhR2kyXXszwOG356+Q1c5gAYwQRUtMisMyEiaXPC5wLA6c46xm8
0DeCxtmqD/MuAEP1XDJV5XA9DunJlPeNedgz9MKmLrg0555ySfEy+R1O8SrmUBI9gr/391nHj15N
W3Gt2dGuPStbSuNr828lMDqGKx5PG2u8o1/RYrO9W1VMWBByGUXhrAQ8sM7oUHCZ1Mq+Uc52kwhs
asQgsIXbHA8TvES09dRrg9jCCpR6xkNtC4SwrP2Pq/anPmWnKRQwP9tQrnoVAJXrW3h5peAUfNYU
8qWAkajNo3f+FQlLzMigetTJznuuL522/vbS/3JXR9B2c03qZjb+meKCdcudRvyxNO7+9IrSwBVo
w11IYS/9x6BNMlTv2TdjPEaUHZ34VNcs0xctUHjbvjqSUmAa0ZLCgi+e1Wp6V1TALSercMfaNx/8
CoY7YdFKmdawcuEeaJlCAkfRhNM/luHRV6T5fDIYCxyoIjoSXOoZ01et+qBSKrkXegt0jkzPkEx8
k2FrS263gw+5+cXfxRg8xLFJH7W87ZliN4Cp5no0OJcGYjJrX44PuBPHvVGQNDjy2TEhaa4aa0Hi
pBFN7Jvt0xBfxsD3BVuYGcOnelP0ZNmTQNmJl7cPMeFnjfw7gIxikRbD7O5Ltp71pWVzD++1clIW
wfHJHyzGSEgC5pfo2Teg/oQE1uZXCqLk0kV0YPZz/LgE4KdFkD4Ya27rGskK++vHzdkk6ZUoJRYx
Q0UwcISkS1N0FW5n/hggSczj4JpyfC302s3c1FrMbmvxhttR7GQGRe/dHItsLHejszkhvWcBFVcv
fJwe1Hahc6u4LwQ6UDOLpfWelpWYe2BSbsEfR1t87/HiQ33n8nVbbdt78tmYG8MpwfC7cVPuNBTw
TYWhNojuVXsnHtXkX14i/ZZdJRkh4eElh/mMTVWhpZ2zy21F0WnvGqblpivbJzNLdw20HCcbrZqh
Z4WaYSDL7d4qL5Pli74YPniyID79U29n189oBWZpopzRvvrlP2h89H/UT1iHc2J25qi6HS6VYgpL
aM5fAq3IgW79o9dTrKMVDn7269aWQK7i1xfOIdW6dxKpzSgchEr6Iqv7WCCj3P3aCX5hbqLj3FlJ
h9XiuM5zZjukeqzoMU+EmQ0+8UimGUpZvsY/RWmpudrs36QygxmdauJYvqtEPbrjzii3kzMwmdGQ
b7P2TaDqjzt+F3uaqbQ4nAgjVuRrW2KEb9u/XPE36B62OPGqVOSxpus6o48cKJsS0S+fzaIe/W4J
YlF1N8Kh/TCpyo4567J+lZNkxreiWrPp+DdHH6JfafAYHulDGQ32zJCunoS8IPVtk41vzUg+9QsJ
2Y/shx4kLQAM+543WdE2FQGz0Omzk8PLvH4lxHdEndBzDtUhAcWnBYwZTq8yeEYlyGPh3BY5lemv
bd8h/YAJPnuQYIh9CS8O2I9BCLiAN3cZQuznzJhswljIN+ftE0s6VR/YXo4Y/nBZOUDZR3TWwkca
bQUpan4vJgzDPOoxvvsGe8XlThIL2mS4M7qFVY/fwAoJ9oUNTCabeRDpIZAkOrXdA0m91aoktlL9
0ZqPZNwZ87xMAUPH0gtZINtiawkt875c+9R62DBZZabV1LXh/NReAd6uBv+nMlseSsmbBBzroyLj
DlqkrA1eVScGAJa0edkRnnX56J0bbhUNR7iPE3PaTdsrST6eo1NiHN8k+0H5rmgK0VtO8+9kzitv
m8ika9Bdcpcl0O6qJUpU8Qir+D6IJjUDZy8S0syHdnO7tVLmzQyjk+M+902vVIvlqmHcSKe35r50
o9r3MsjPAIl5W36BRuPt15QfCDoq07OZ/iM+l/5QNIviaes8/VITINH2ygOMAZ9M3JiYBc7esT84
0ja++Osl6gx+oJWyF+2QL69kIWXf5T5EfMDfApvx1HAxtXaGcBMpzjXPRdVKLSPUKifN0VSuSwy2
YaSvKw6vm06UO6B8ox+B3e/jmjV6TgwN9QHEgHN9xpwKY3Gdtl/3eXO6DFjwZrEF0LxNB7w+inEF
2JnE+7RhCm5PhcWZtnuQa4a9Xk8Ba3b0UAIJ93Lwycuo0Vm3sOLPfD556BZFM6bUYUTl16GvaHM+
Ihh2CP/HQzI7iT3qlqZsVwgzPNhQAFRjXGVjnuzEIUicjW8kTmkIkgwMGh2N/sk4BS2EPJnrmaIG
r334M79q+NZM9MjG7RVuOuhLx4JlYlLA1hAWEJXeQKxWH7t4skQPRcTd2rD5qE37HItljp6FPOIS
39yu1edPDmUiig3/TzJKa+do//LH+hMdzL29TksdxtRYlEMt6+AC/fNiHjeN6EYxoJ4Qc1WSllSB
JDvCt8X27+x32Od4/mrZU+JtHs878H7x6y8VKjKZlR12hJe6I8G/48jbCn5DX7FscOthUnVeJocb
W3EN8bIDFDcJxNAAy0ast6aPhd8dc3Uf9qsy7tTG5oZvvajBRDYiaieFM7uuoEYB/vMAOYLVnQ5v
GJfGt3OxPOfx3/OAeYRKSWdDsc01FynMmY6OvLLFjPE8iVwLmOw39l1wcPLFp9IFi+A5WulMAfjI
cfApq8DO6r80G8q23opRVnwz/dEdHt98KKPP1NLtZOcbvVnxNDNrDwliVSiUOiC45HumQSnStwZW
e3jKSjbvwgK4EhNmQBPPo6VsSwfvb4rmZUSl2GcuU5Q4iOFujS7G4kroG+N3qXGxp+4+xIoU1IjX
hFI/w3lUtbwSMkWe/3/se/usS4zLiy5vvNLpPQCirJR5pX0qYHkX+qB52BudhSzbqTVFrIDtI+GR
si0fm4oV95LfzQLDC3UNvuqIpBnAa5XvbONudBZKIWzmqIKlH4gys+QED0TKVZF92AKYkhnJzddO
IUcggRI1sGRX05FrVaq3ipEzdFBtlX8K4b6U88EwDfHsdHkuvz4lOIk10Frhsiy15SYai0axXk/s
3g/l0FGysf9nM5lNWF8FMhmLEYxy1NI41JkwBYrrRIQ29F/n92beCbKxmnm9KbJ0ujITXjEoKMLH
gfInsvK8M6gsOSQKd5dozxY4uzXrxcFjznxAiUT4iKhVMzj9TE/m4NrL+qaAczLIhGa6FvA6tOHT
zMzdtGTGz/NCQRUK7Pe1hIDuhPk4zeyd8pxzUn6WY6gt1IoRJfJpHwrNcvHUWhCyaXCt24SV8uAG
L55HcFQR5yt3MD+I34dvO3fEBe5x1XYiL2QK8h2Asa3t/Z50GSaJnODqIxrOAqnwr2DAnJooH1AU
7uMPqgwotXK61Tq134NIC+hkxZrxvop03HQiprfC0qUnfcSr6Wqjby4UgGybS1UDrJiP4BdKoPVd
pYUhbU+mjvth1xQ+Xanh2snJo92Mb5E8vnP2SnWkWyQXv/aY5FW9gEysA3CTVg3L1IUTKjcMLMBP
abpgpGsf8RvL4/6HoEPgFI3mN3zupwHpBNAsQ1f3GoFqzPwvtwea5en4xVJhaNn+LGeVE/2Feehl
t3EEtqhkgO0I0yuhYWyehaRgPv3LdviIyjHfbEdU6IRc6QU0A6ReHldlbYjvMGRQ4frqcJOyoNLq
1qmnvWU6leUhliNOsznFuVmR7v6ORN8Cltr/NPfZdrDu9SeunrM+ucIN90Mi8wubtNso91TWOFEl
mL92D9lBrH80ZK65Mke5vRl4X/IvMt74fLimmWcW68dk09gkP3JqYACAaBvMhtGoS9X1tN/jZ1Gp
KRaQzFRHVlk+z67BvfjWeRx8lc1lbwjryu0ReJ7Jl193ucdDlvhFleQMWMDWcg0YPjgbdzBhsopr
e8tP9GXA8NKHsU2yFy8tHcN662gnJD4wmiBIgQ+ztJMC9UDmVjh55bv/XeVkiLJwZhusBKQuhPyZ
dEsp9icrTTVyb4psXNJiU92KUP9B4QOOl/98i04vcoNhn9JEkd0kTUGFkIG1nUq2L5F9LSLO7uMO
2kElLOKbiz62zPkeILZM1T/1Uiug+/XH8YIdd93jjWrq6D3rrEVG9IXmcTd1PWYyVNowg5VG9xJQ
OoY7Gz5O9fy+hFnscURKhSoGRkez25rz77BZmHdpqO966/irDK2hldpQQEVhGvaSK+Ou0foVlhLZ
OV6sR2yAFmOuUkz06AYGUaN6EsaVIgXqX7NUSL273KTNhr4uUdEaUALESl8eABzkjU7C3ca9n2ah
ZzuqQMMOkD1y3buWIYdi349y70W/oAf+zUwgGR6iC30uI0eYiDD8SSNQcPS6EBGbZEATGi+gbN05
MUbMci5aP+jNC5D68k2vfWM7MI0YFVuQhfNaxWzuRqOPP48mQIjHwWtQUZq4g+5aDhk8OB02CdBH
CaS1aTYOnTJG9LSOeubclxMJ/sWWWrz6ubgCa9dQehwVcxjOtTG+9SJgUbTQZIohr9XP/niuoTut
ocsSLCSawzWfVDHVOGKyoGwMjjPmMnzSE/hMCVGC2ab0iRcR8SuSwxFV7N1cplgA27DpIPWHcRrB
GTcDM37nCFUseGQ8XEEmCNlxZDkYMaMDrerbZDAS+e/BwkI8AOSR3QDQNCVcvsRQbMwPWYEBC0Cf
RxlJnEIzZYn8fXnu3U+iu7tHJ9oNmZQ4SUYVxvPVNTMeNET3pyyLb1aH/KoWbE7Zx+tMzDQikJ4l
ccAsIZHHW4YCmHgslzuhBQRba/13cu8chSi2ROaXl58BhWuS+Nzt/jM3DwvEfor4etf6CV5u0Lla
u8N05C+2b+IkZak7Us82GkkVjEnKlh+7o9nW/H2Afb/E7/54DaOVv+w2jI/1YQn19ZQvUd7gmzjo
vvNXxMLCmPIV0s6bqgy35DD9m3pV38Gi9rhTcw7nqMz4leYUll8HOcAguiwvs+bYsCFUb62kwCH/
HeyQW83ByI8pT6D2E9ijemd6gCl2YYfj1MrzDWd+a9F/lXAGi9OxddRnEmoWcA6pSWv6zb6X53EY
cJyaZ0ZiL0rQNG7xFgUwvR3DSYkbeMsBbdb/DCufJLiXS0dlufQBdU/jw7AKc7jY+d1JudcfB+II
N+uPKHS5AS0gf5FDzXUD5QLCzZWXOu9EhgW7AZYOBv6zmGp1cRX3N8E/SfAGdj9Swhbi/G38I4hz
bhcJEkqCGJFwu8QYDNDRA2JQCylRkuPFmidz1SuvfQ3APmQRgnTd7K2vDE3QVJDM2PcV6hEuKC76
HmXphQcipA1+/J7fnIWjq/snjDVD7xokSG3eYdoMns2Nm9iRmxw9Vy25wDfxVMY8BZ+wn22354lR
J4qbItfluAIfNDDHY9Fn0PK+1gFDV94gH4KwHo9IRzBQd4P8wePznpoeN5+3m6W4/iFpBuFsCg7f
WbSA7V5u5MKTTZ6uYPjrRZzYib8xFjfk9vIIEcqI9DCsELDVKkvp7UBofndOB028MQ/aA6Js1Nag
Lly7GQzGP+nKicDmRd1mi8SvG9w69F4XrJQ2EPaJSw4RXU7Bj2SYwON5MfGRl9xEBTf1eO2NPEcY
hnWAtOx0n+bE0PbD33hhZvRjcdmnecDP4gYeg5oz2H2D5oiZBsVOhc5Mv5Dv+Gz9WjCb0h9HaB1Y
ttC+pqeXVDxFtjyb1JOVkziNkOoCqkcDydYO4EEYIJWcls7IJLRgdCy551roqiUf12jshvaFAxzp
lBdM20h6kM40Otuk6a6DMzaV5RgnX+oYnunBZqTame4U8KhsL6BclJhWcSbAKezmGf5NUV76Hiqc
uD42EtPlbiJBJ6D8kJPVEBSyGYPqMon0oVQxy4NTfQjNGFja225/a4UaBQ9snINSxOb6oQjDMbli
VC/r7qNZkPnIRJ0Hxm/O/5U3cLIYS8vZRJxw8Dx/uM2A4sl0GDxZ/ADTd7ZPyJIbwyDQzZBM1vVT
dMKlP1sDTKR6DpBaBsEH96n0eTDXL36Lxv9VRsZSmr59abf1wPM2c6fabx2wnj+eM2AfvGGVdSU3
4IP9Guc/uXP94IsVUGWInAwdNu1Tu97zK61Z9gIEV2GZrE9oZho8V7uDubF0Mn/m1eXQybnroWtX
LVEdNQteo6ypGgonFguT3y61J4aShJ4ZVu7XA0wXwoyWO+K6p4Zkj4EqC7UnjFloPY+LuOxkdn86
qmjJrzbJcDaBI6C/uMz0yItgQAOX76A29J9SlzFjOHoiYbpu3HryP1Cy3zm5Pxa0yuw6cWqSgEKa
05+xPv8OtsBTR93DtV1CFt8YkA42GBcAzrK5zTvI2mpq6PjO9sB0hvuJbxAy5HVLHl3xjYfpLZnm
qMsRalmJL+363vqZDQ6Fmmhp/ChJ/cq0fmtYFpArlmp0kZcd4xq/ZCXMHGOl6pM7nGQIoC+aBFV0
0/bJZu1FJi3Yt90NxkPAgvRRWqBvyP/B6aZqve2D6O5r6tEvnDHk66LzfKLDQwy02oL0LhoCNtae
+o8bM3PSTbb2cOvUfuQt5BzIgXztbzkJcHmMlvGr4gMsnsZ7tJs4LbVs7wFP16lAok6tN85nelIq
HZGiVE447NQhbi7r/waiiiE/g4IZcgpvv+VJXT8aWrMcwFFYthIYpJAzXlEzN7QtkZlYeyW98C5z
YtiyaeuWNY9/P1ibw3kHB0WUUyPsd2Kq4U15BMm+LI7w7oqVmoSPg65FQbUzAnv1gyLMlq/yTODY
rFYDwZ+3kW74MBntmhZwBNzu8o+eKiKzx0ZbAViCoBBbsIScu+9E5cdxOyN6kmoLjKhEPnKebP7V
VfDleJhU+LSFDf9Mdu6EwebO0+2gaiMObwF6ZGcjxYyLu/i9Y2nl3FlRUu3noFpCus6qTqbS9/rO
geN7eTx3bsPdYSqHJVu0QarkCMCKJFxEro8q7NBuCnCsrer4RbtbCJS/2JPQRPamMGIGm2vA4p+8
wgq4iryUwr/LZDeUQcfBjXJ233BCe+vC9rR3VcNP5/Kb1+7zNog1qI1wknzBNEG/lCXkmEhAqccy
3Xj10BUgn6kRpU/CMMIlyggOdOp68wdYPGd59+tN/O15003f2N62ngwlWtTM5odOtD2T7p+WN1Zo
0sIqXXCnTwX5HaDbURG4Fmch1XxZSWXUiNHdV0eoLhlz+VGYj2WTuvGLGu6T6u9jjI1ZiJRVoy4X
ANv3ymXQzh9LK58K0vfZp9jKaMR+hG+R0G6mmmz5jVX29uBGsbdqkeTlt2+pxb7eJggcTsXg8csz
ACg/is8r1zFgNsLJO3F/tAQokaHGPlTy1ZLvwwUL9czpeNOdWPqbaCu9MBxnpQguRGFVx6dgG4ui
OpkxqAslkJHfXlwA+W0F57PFeHE8JcE+ojDxxaBoY3lICJm8sfAd50HhH0EVdKxJ298Du0F+lvSw
eg7Jxnj+PbXYc5KSi9CiB9rG+heSHjDvhMVv4eRL/QBcQDpfSqTwLoAVnNprNYvBEehfpEhrnZxG
pZLwNRMydqH+D4sCRpGS6xG2ZS2rGo65W6fBxdBuEsgA7aMuZwbPTuhKhCDTd8zxCIf6VXFY0IIH
hp0tJedl4LiK71AH02Hlu41XxbssBBfupw2rdnUd5DihK/jUyekhXGTiN1o1+Gu1aDksfP1aX4Vy
DYY/FtxMdtw1nV1bQZESXrcANG6AUaBp92eA3LQpBARHPcOn83VakiJ7by4KU3bkA9KjVzQiHr5I
bfneq3Silawe4fMja12e8zL015bYsjZKZz1SHDdVaBxrgW65GxOMN/s1ee0070ZjUQEMM2L2RYyX
7V7qK6zX+T/F9CI4OcL3fHvqrGr7cb7u9YrU5J8YV9ETASTGfGMsuIsL/Cji1LaySFS9A5rxqPiJ
wZJgjx4jTSdJMDFrX75+wtuQgJ9cJpNzIJ42PRTQ+pKzuFzY94RABmjm4vyUXlGNPUlKrsVWy/ul
yslGStvzXCbYN7QmpgOG08my0ESPE1XhZfY6inX/kCxeEb+lOR+TG89bBCBb2T15MiluPdCNxI1E
vcpqI3i23DxJP1bZiPd9xycYfpXhY5WEtNE1yFfFP4XfGHuqufrPpXlT49LiOA0QsXKPj052TIJF
zXeQtcVZ3hn2gBYOLO0cQA6R17JNJF2h3iNLF6Oj1yr4IZvoPJF+BUnQgH6vEHW2Lig2kfYErPLe
uQKqbZHE1bvHKJtCHqAqw8tA1AsAERcvgNqHHLy2cwcogjL1637gbQlkPH2f6tPDSJaqJRNHSJ5r
JpRX19KmPRODom1b4sTkEHqFtA/BarsAke1mZSL8mF/qqfAj5ACwOpwgpWH07umQcbB4Ec39yQF+
skaLyPPnD+3Hl8iP1s3gKmzadWM9E5n8hjuZIrv4PV/nUchIj+lT8hh+JT/hS1yb6hCbCsd+o1aE
t0babVju0UbUtStojQhuO5wftn8uFZZwMfh6G/u436SBdMeEnuLTa9//LleaVCAgYQUtW+UEsJcj
tXoKtxM/l2dSrBvUx/a6gzOB3B11Su1oqpqpYL7QdpTzRiL/hsEv4Gj9CYF8DgCCmzXoJjoGG54I
a6vljLnIRhISADd/pj2cwbvb3KDy6FQxmeLSoyNHTjnSwLDUiCQyOHTmRwiVL9ZqNcu7u42pL4gi
zj/jIbwVeV7v8dTBAU12l3JN/WC+8Qg0IFCnE4prEScMCW+ZOxEFQR76TFJg5M3GvPBeyA7Y69fx
lVMsyucs0U5m+ZGYolObksgGQWhJr30vOqMitEBI6zE5CdzNOEX/ehCnj1DDjTl49ymq4xMCCqdG
4aezuaanrKfwGsWFRbX+sPaT/CyixI1aRvBRwLzojaRHhA+Qb6WGcl5wjUqfpGN/2DwkY/DMMyrv
K0d+TKixXce9UmBQZrK21HxUcIc0Gdig7EeY3V734Ul6BF9hQCAbZfiZerLlJAZSfED9qDUhIq7B
2bjmGnxiRkoU7PrMdEncUuhCr4D2qciFapn/bMisxA+M+GxudKsYu7vpLEwMR7P4+fsILmECLQME
l+7c3hAKUj9EbDarSwCHmxeCx7lWGJuaUeEs3/Y89iRI3Z/V3yGb5E4+AqZC8ilzlLDzNsIdUhoP
rTrlaH+Yw/5ZQTNvjtWh0zHeGXkWE1yFnB0t3FJ0dM4hs8+QKNvKlpt/Vf6IiPnW+uIFzLOOR8ly
BbJmWEjhfkZ1wLt0YDC3l87+4r2JubqBOryFTuRxuKMaaKS25qVhJVw8nUvkHflBQM5HCchlt8GD
YH37YPFLs15E6iXt8YrcDhmEQ5NsGCG33r/a261/iNQzFhQLoBz7skTlQ4EV6k5RKUWKGzRN7kGf
wsvsWpqJOJigpOI+rQpuUfRPGi/t0NH8iU2FCnT3Itrs6YsQsyvMD8P2qreoHnszqlbYwR0lC6y/
rE2WPqtzK+frtOWJT6w4RnlfV6zUWlK49dyJODndv4KyLuOaEeo5UBPtL1L9PmKErf6VLNqhvrqv
a/EDRYljnzOivGqy3UBTxDAWyzU/LoydvUlVT/SsKI5znMqE3PqoXDUrTDeW4Exps7qCrynjvpOw
U9xkVXYCFA+3KCSanxUX1X5ULkUpyjxj0zml4NDLJ9d7ro224jQZuS7UWb0l49Cclg9DXRlTCkZF
lzDXGjRvEeTCi3eDj+gR9Ez691bT+1mdSbCyEFrkQa7+XFeJL5ui8HR08Fdn3UmPWpcWV0Ys4wEk
KV+p8T/yuJcKv+bs5yatxXCU7Wy/+dBe5UQPm1oS9tIHJBj5BLoedf9uhPxYdW3ydMhpaTONopBL
eeMqYcPlnqCTO0BMy+NxLpstuASXCpFnZsCU1CqVAeIVlyEEuarNKoE9lNLhKo6j/uGjMdLfKiO2
l04eIwibEE54Al0kuEnpJvv2C5E+kIWgCC3LbmI2IS+IQMOtP6jQ6GGkr71SlwMyw/LqihdvsglO
CRcgiJh3DmeHIibwUGIDkiyj7rRUW0/AWpx/gRMQ4fUSe+7SgtmYcLIo9O0eFG9dSyLfBhGdX+ke
1nV5CVASHs/q1izQjbatG6DwFH/TxtFSDFJGF6nIbqfKmOuLEs6kVov8p5oND+D8SinKLZh67Xfv
YeoFeffg/XSZd2S3tEcVBAH6ARugn1bQ9Hrg9Qf8VzG91xgBLzqu6qtsTT4ziZND8z09ItOj2SIF
+UanNlssaTqzphCMOrMN6vvqew2cbCyslWiHzljSjVdRCCV4la8CWa6uphI6sPBg4Q5qfbuyZvza
bTJLzXI9Sto4qXWrC8zTbECuM/n0LQG3kzzyWLJek5o3G/tB7swA8n13PirMZm9oIgelGLpqUfCF
H/8W7dfCFyn1m59gowAnJPPTFx40/iCxIq5vOfkiPfWLl8gejCVV7sVpD+8SzQqwsLdCrrNDFrgy
gdsLmvG5lQeKshPz/bwUBDv4j+KrxtJrWpAw3ALtJnlIbzewo0VKDJ0BKillhqWfMEfwdQZlaEpt
DYwBP18C0Rtb+mfbiIp6tZEkioqU5n9yL4osYGThhNCE4TgurtJPWaBG7+/AhYTS9DYac8Fv2oiW
Q69RDakFVPwSvgxNLwq+KYAN+Ns7ZiN+7eYGY2uUFPWDw9K6+kUSb8Y2sxnGhWtg4OA8qsA0GbRO
Wo5ZSG+HINnRmFHDWuNhUcTDbE07iYh1mbs5HP+bJTrXAjKV2L7/N/Et/wcR2vRr0woug6DLDFyG
i6mponpJKKgAEPikcoEfC5u1Z8Z1b/AagD5ht+8HWYV1GB5LnslW5d26mL3i6boaniAhYLLmnDTg
4fYFUOc8OAnSU6cpmc/VXUsRQe9m94wfJVTuqyyzJ7fYsfcnnrvtDmGO2E044rkwCFxYq0jUlTD8
hdmQK1ZWMUnV3C6qJ8G0Pt6owkyXHSf4SBMJDVUr5A9BJ6wBJpGm1ollhEXxsG7DgTCIIYfn7kOW
5dR8oivBdtW/vKxbiHqBygS9J7HbMIQztdYoda1CFXXbFU5+bvNAZ8dGqhZZeopHg0VQLLCP3XEH
qb7qXA0yOKqidvgZnHJVRScsU+8YwCyGWCux4YV6aFmX56V6daAEQGcAIz3HYkf+GxR1RFeOtvHx
VJd9JeLy5FszuyNE6gxfANI0d1Uxqgv7pZvsHuS5zntKO3qhIGO5/+XQAASaOdIHHt6wUWjYXEfo
t4JhmuZ1fuwjIvEmGzwkXiOCZ9fCkdHDEDQThAk2iWY6BK5dVKjOJiURqt2MawN8lvpugC+MfNsp
6r780Qhpl8cG0zj1/AWlyugE7xcqHt8XxI+hiD4Yz1Vob9kPZYUCCdswvU+GvEvpVZG0yRD6bmzD
HvywdS0QeZAoNhndwUu1DGI/CZWn0UXxDRdh8gslW/cVtDcRA6QipDkRdafh1aZLX1Tvne+QMIf+
KPcCJ0QmGJ3T/8W0usu+UirxXUjwLkEaq0tduuPYP2m2agEY3Bos0ERb0Yt8kAIoa5AjqrUWdC93
PAOmWmTjnq38OUs/4arQAzg1LYuiGNHH6ggWnW4Ao9Va4XShB3WvEVB1VcIqrF2qi5nNXAdFal26
gQxlB8zl4cloygIIHmFV/pLPVUie1h+e0dwOguY2ZXIDPNWyiAHhDuyGdtJsk6AVY9S4lM04aIPz
zi87EUTzRuqdgBUzQJG2ShWJ3ZzYQGhkI1UY42CuJEtV+yvZoPuVeucq8bqnw0oQRo1NDsVSVcV0
XEOnOV+lW3pJoek8YmjncMi5hM1LYzKX7LGlb/hcF0Sjkf2oNJvqLYWyZl7qZ6wvA6sToOud1rjs
wXbF1dhLdvzstDYZkxXFnPh9SPnDaFjZA7ByKyHIwKKGEFE9IAKXmONNHHMFylTM9pGEFWJ9HMqO
immHhy/7iWf7UcVZQJME4c4fi0yQ1m4MZVuOjDzK0O+VuMZHjAPmMdctMnH8gHqpzOH7hGqNX3v3
JmdW+3m4xOtYg3bW2v5Yd11JPPJIlVUKwgOcqJCeULfL+rx82MYhkG7ZR5MnFqNbBakfvuBeFD06
MrwOhh6jmdhd3k9OyqM216ua6vRc72AZcFB5sIA2BFpR/UJp+aSJ2CICPhGwCUij5xXvWsdANTEB
0iHGqJ+7GKFwF3l04ArwN2qx3pEblfUWTfSO+Pd8fwFmAehxf74t2Mh66pYacd3ke0SeHXNdMN8S
uVfnm2Pn0EFrV9jRIGGsBEARYTNFlKQ/+njVtocHRXbKxNC+BdtCOrENFzeSEwHmAvNJDiXCFhXG
7LHjCdSmXVRZS44Surhn4hcwo2AGx1IguXl7O4xHmdDiY8K/RXtAAbT4Si6qTYMN3Wuxw99yemkQ
xR6d4AuyoAYua9XAwiIWfiNMfKo6/jV1yl8pgO5dAmzIIV/SXkjLVOVZadTbQdCVLJn1c3BcmKGS
9TDO2HFhGRi+Jg8LbppFzfBlj7OTQvPjTMROcGD8dVkq52oLuKZOMoe3OvYncWeYj+2VxAQzMdQU
WdGzqoUE4D31LdrpB1vSQusDLbBA8Jhb2GkEEimouDxRREKbP/vBWcrlbOtO8Pf4Oc4ziVz2Vl2p
hEp2rdK/5XK/ee2jgbgpbpJrMQIuTXe6FsBDUubOtZk16vIk/R6IypayqVuWanciTEFFhGI5Zewx
70OIvHtmJOVTj2DXip7owikuudkv2H8Pq137nGBn7VQ44y9jktQeu71401+4Jzdxr1RYVziy7LrH
ID2x+ysIazZJ77TugRu8CZCn4WZqx5ZzLs9xqXj4nKmc0tWlM926Sld38BCEBEIDsCn5FvoDe8Zd
Oe6XlJGtozaoOszkeLN2gyNuqiUBKFvFYJxvBGpDI6cn94XZJGIXhRRQlWHPidDpJujiMfuDueLv
ggTwPu1iWbSciEzp4AoG7fmb1KoyhVsmUYJlNYr9gWc34/+SrMh67ileYh8Ar0fjhE4Th1VGbpMr
yHWERUA3OP/5P7dFKj3VypQ7wBQra20wv6o1/+8t4fa98VSuogoEPnj8dUun4hplaI3Epyk8Mz/K
jqu75JRdspqs9Vw75iS9qVUzQ5w/2IYxbJ26CP4F3xPTy0P8KK8/maheTazoPsIhuMP7N7KZ5WHo
loMVJHdi8VNa69m3UmEjCYKg1IreA9F0zMmBdMj41yFTVUVf8s9l0g63OKgB6qeqUuSBbufJwpv/
N+8gFo+++oSWEMmARFto2WgQRx93L+8rCqjRXEdhDIS7gYlvwssx+n3ohEsywthpDQZtun5Xwy04
Znq948HkhIiq4AbAbuyd//GiOqBjj9rRG9G0Hyp/wIVTNc6sZ6mYqPp255gmwVskzhQsHlINJV9s
veg1xtZLm74GeOg721YL5Q8BSB1TbvI8W+m4nyEWGE1403N2PxFMzGAzGFDCdoY5W551Yb1ppw6c
BngRebSkzMpT3ciz51kcfp8/E50Shu+/494q2LKFjSFZFUEu/MGG9JDU8znF+fIpdmMmpofqOzRx
KWTfjAKl9/DuQC3gLq1x2IdY5gD33KRXnVBbJdkNBlx4tBDL1FFSxUX6FdBikO1is8Cx8ryZI+M2
tNQPRN5KFILc54eqoGEOBBmdy5RBe99AjBjT8HfRSENXBxnPu7I6x4j6J2R1ccseIXOinb9KZPkJ
Es2juTeujXryKxSMk9nkhTYJ0kkylUf/FCGGuUlHyGz1qxPF56hGxGi+ndAtUZda8PFmwFEfMJWN
x8+WtkdwPB45U9WnbkX2aOxJVWRE1VMSIE6+2HSwB4B26Ii0qTfL0rdoSHA6buRIVAB+kW5UfQ6c
Ok6bL1twFkI+YoyfEnNvJ7NOBsP/H5TKo11lkXDHWNnv/t+Hy0Lp04YWhKgws9qumZ1aZM+LgiSz
R+yN0XPtmjSi2GoLqB/hxYeVh45Am1Ka9oUI/3/zd7C9AjeR3FfgZcQFSL1AQSgpVO6mc2bJtKD/
dfAKxgdZ/lZxkOwvJ+XKf4sLs8sj6kDuOQxbNm3pNKcUheXqY+IMrGZL2YtrdUIuS7zMFavdRw91
jpJCrVyY4f8+Gr6FVLJ/HL2YtL5LgOKMdVU9ifAeMk/UY6PnQs1vX74LiF9J1Ak+QiOuy/bIBe5/
XmNjQuJw3woHHdFyZjCwcnZGfAU/zdIZfzH5tvOuMEzHFk+KBT5CxGHSPnEcA/A9mdm5CYKMSTw6
XxdLUgO+HtLmIXJ8tJxClxiYbSsCPLRioLJPeFotocDbLr3GRfAFdURgoU5us4iESjYC+qkvfiBS
NGJz9L78RTa9Ewpa3hzmawOcrfXlG7h+VTzWqGDEEZm2sARpQmQ8UQY9ckHfCANY25cNIBOxLP2x
AhloQFALV47rYY/MHZXmyfrdD+udreV8TRs3rYqVHrxj9tgdkdG3um8g0g6gq1yJ9l+gu1j7HYkK
tc81UMy5X10ImcfIzerY/gdZb84Y/e/lmO2eOdF59CoqXZX+T9xpwhItE8+tXnLyIcVjGmTsTz3R
87E0BtjLMzws76jj5IedqxOQal3kR2XBKng7NJc7EWYkWmfkdlsDyJUOMxs3MFy2XmCUeOj5o3nn
WY/L5Qa+3agO8s1uxe1wyKTRNf5j9lif5R0kPlJoEJJRBBEjphNwS0pLQERDf5g9SMeR9loVXsbK
gzO5ktvgjwFRPFKBM9+zbapn+TpwR9tOfvoD9GwkbmIE8pfjY7nnMCD4rX3SqNFY6h1WNc71CVZ8
gIAF/BiohUaSqsgjeak4NwC+qcw9eDSttfkXBVyWYHegzqq2DADxX0LN1IIKLef92UfntG0gbXV8
fi/zuWNBXhPexPVb2SMT2MtBrzAfeTa1kegLQsc1Oetkdm1fpxuYaeF+71zbeuUC2Gu3XgcUnnC5
5/ZvYO5vQDU1U8ScMd0S6Zfg21G4lzb763E9eeblodLe47Ld7t4u53QyEJGKZASAezXxBJbnUYs0
UwYVUzX63PZ+89M77Qmp5P11bjR9ksfRXjg72KRbbzk9fNEv4208JHzUGBX+pnzNsVGnYWJepFeU
xDJxZQfJG8jSF4CG4R4vvkSxkEs9huihiIBilyqU8Yb2QNWTja8rsf9TRE/myC1p2hqsleu2xjus
WNOr5Q5+RTWkvf2Xf9GDOp6NNOuVAl1YxM5QHK4Vg9DE96U+xVI+jSb9YRPQ6uec75VidRBJ+xdP
U0DGZCSLYuW16Z/io+bvOjbTmbNX819JxSMGbru7/cbRQBTwshon8KWZrk0Oyz7kM2H7HAxujiL7
d3uMh/D1EQM4zIKt8G3CJDOG+LAVEWo3IpDbKzw2c+bT0hauKG5zKqd3/par3cKkR6H2KhcjtjeV
k5b4Sb4KVLtcqBNyPIutxGTXaIcmmTKL3tflY8aV4nQwkQA+kIA1f8qSlwC5ne34K18xrxWN8uSl
P4jHFYWsV/9MTw72/4D+r8b5T9jHB7eWvzCElpdeJM7WfcPL/XNZao3CncSx8Vjn0Wnl5dXOBbv1
31eFJb1GgXRj+mdy4IMhZjV5Y/puuzQvN7CaOOXIGHlH646/7Cc60lccdChTyxIpC2n6GLWJxh1u
wQMiQ/+s53aE8TOg82zxE6fHdo3VuNS4Ou7idmiwverabW25slboofsC6ci/nUi0okmm1eA+Zj2t
Y73dWr3DPF3RtMePbfvMk6cO1deZ5CNggbP73IQXAwnAEU6NfCMGslleO0LCm8hue2AVO7zG2fMW
K70w+lueLqtkCRFfrPVCHigAcZsAnNBX+S5iyqYJawDUprdZVDAY2Cd0SLg9mBM4mEbefsMKS7oS
aBNqDrr0gdRBwPZOvPwEtv9PhUSF5TPeVLWjd6qSk3cCRrKTatI/tA4rHOuVNQIHh/r6rLDBcQQ+
JAd1xii7ZHPyjzraCorW4eDRCwi4S5Z3d7rwwn/lbSs93FRe1RutnfMDYFeXfuFo+TGPQ86zz3+/
BaoGGAuXkEu9qMO+dFtcI1E4jGEmYsfEbLVOT1TXxxUoDEhzQPcSE/O8y5qkYY/SqilM76lB8zfL
ULv6VS98nqBo05PZ9+J5c5/4IvN7RIugMmdBxt7rYpWxBE4Sk/A2fb564h/I7anayEfXb+VITo9m
Eqcw0j4HEIemeCCL6OQyM9zVhzmdysa2ttn4QhwKRBbwTqix/p2CHOLjjfy2KBpuKlkJLH7lXl+X
knqzFXX8bwAR3Ubamy/kaQLwC80TS7v0fbxi8wRPrOyiNbmiMidz9sO7lA==
`pragma protect end_protected

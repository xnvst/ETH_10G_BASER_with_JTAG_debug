// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
a8TGaNbvBE2+8y/rwJzAyTeo3GkU0N8fJKHELfSIZZTv0Doq8VmVHH+yKgHwfBLt
kSn0W8ZNkHjMJn/hVr0AIqxCjmhPKbQMWkfNiAou6LdwCdN5hbmXftR5aA4M7q0M
cVpYID/N7woK+Kovtscu1eR1BBbI0k+zh+5w+cdKszI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12480)
zEFvYwClUPCx//EI+X0OAceUe/M56GveLol8NpLSezSds5CjHIl0kVAPVIpK5JjQ
03OCO2u/9wuq25vqqZt6/tYNloLD8yAs9M92CY13QL64NXGZbWDOT3OYZBdtgM6B
eGd/4zw6qHUQk8+Fpa+6FIwjM8GbVtEJypub3wdrYzNM1JaotRHr+JHRsMtI1rRB
iTWPCin+j0Kvi3KddQ89AuM1gdvjOeyBm+u4cC/heTKXQuE/Jah288kzqzv2j25B
jcZkOYrjWQ75snQPnPux8p4zQepOyvg9/Dsr8ywHi5UIqRdM8PBEjFt88OBNrzP8
kapdCsRdjdAYTFQgscwZpIg8hHE5uFnKYXqlf4tmYTAZNNVUnAg9HYgoVVSvSmum
F94+5Y+0XASO/5oa/TZbo07Du20FfEVtuAPnNXUJC8634MtXEHaYnPt/FjEHbJv8
jzFZV3DOKCT5aOCEzD/rqH1eZthGW3OhKLaV13f+4ZKZFs+9h/de2HTOqcFM2c9q
dSaT8aDViA+bQxjWta6xOHEtNk5KAHuKynuSS00HY/CO/YjK0Hs44+4tYOPVR/US
Jyiivs8ZyPBDiOFkaEfCpMVGqdjSV7yLYv2Ht2OX2S9vXmS6gV1tyeodU6CxoYKP
hW0MrUVubZ+5TPXERKVvwTRDzZ8bQg30oy0+fCfpDC6UU07ikwBciY79WeYxpeUw
QBpRqERGG5sjVpwulezRa48Y7h6km6Q7BAnp4X6BkKIMnH7p6K6HT5Ty3ZS5sb+W
pnH79LSjLDMGZDXXCT194K/wLRGxEXax8V5LbZ128XpUbex0nOf1sqNRhX1R5iTD
0wsBBTnm9utKIVCk4k4g+a1sxdsIsrRF691rL0NwYp3bFgbqf7pkb4snT3o7Y59h
bi4e0Nm6Wn6dy4pi39qaTtJ6drPH4UBvTAtfesPIXw6UghOUZ8swZ4cOP5ZlMvpK
36D9HtJE+mXRAdjwghHujq//GYh7ju9um4yVEwHxlaNuBkzbS4XjgBiUgIMOVO1p
GicLzJBVitetDnatNUILmzUK0rRK3kRcsSrN3slYBbdjj2zUdFHT7uR9oIIkzP32
yI4HRqkAl3xdnBV24R+tyGGOWHNH/1qZKkcF53ofS74T2UokN118K8DOWssXigU0
3o7egppXh7oA5gAY7BmX3xOyizoYqsDNiS6XV8P+cd7cs77J4gaL8TVJHEq9eLsd
ZWffl+c50iPqQarY+XRB4iHa0qMJfW01OqdZ84LNtMzoE39c+8tR1JXiMvGsMGvY
81G6wQTft48bjeVruqcld3vfzdGQuphVbbbtHQ2mnI2b8xTdmbVSKIWG6qKPDpRu
imAwJboUOsEG+dbX39By8QR0gAqV/QinjBD+Nm4CWvlzIYKVk8RNUtcz4TqrqIgI
pGPfXSS+dGez/vmZ6eU0riUU+iBJjLhik1N1o7xIrh7q037TiXfdoX+flq5ljly6
+IPR4HkMth8D6RLaM6u4o2WIDWPl77iQvnV7bbR+ru7q/7SUrUiH765AmzGFXGYY
kWN3eHigvEI4RClhaA/JJ3Mn/f/CpOUJ4Ziv3Z643xWvN5I34bJMUnJtZAoeROQT
O+5aPQiPQlOqCZg6DPqmK/XIOSKgPQp0c+zCgwtzRT2pSiFQ9V3h9y8VJB6boFnT
cMBgsq9W7ahNtpVHxJHrK1npI0sPdSqTiPkbeZU9bA28+ZslhmoR8o2GjBSPKaK1
LjVLaAQGS+TVTbuerFXtxht3vauWvzEj8mrt/sKy7T0AnE55x+MojhSNhvZurTxV
iHkHjiKjBij70BRiJlxfVh6h6rOwQ+rXOcZnPNyTTn89gb2UCxYznzerqEwXSC94
FZ0oT81or80w93h1ppBX7L3O1BSpIGDkDmd47uppPzEc7DnVqEfvqEXbfLASOM0p
YouPgfHq37b5NsWerGKcuFz1DDHglDUSErsMiPFFOrgbW4YwIN2Q281GULH4JD36
8oILR3vTRkjKc23GfNoUgsU1tVu8qmmRuIFtBM7lKqBxOINcgzAcwcV5sV+RYCDR
8RcHOyBcFMbkgsKK8WeOQvLblyQ9PoWH0LKacmkQF8DoUcnvJwIWEt5yxEQtG1V3
e76H9Z7Ulq4YrNVOpR+KbiZdi23CeBRM5lTC5KlIUE+CC67DbQYH2cI4JJdp1FU5
XchCDZTJMMHhlCMXxaXymQhurobjZ0SxSCEkHxelIfC8EroeZyDjccS0uVOAYeNK
76Ol8YT8OoKjj0IVqE8+4ywEWKLkzD2NVYL62ew+hJggInEzSjzwXgM8lpWDgxGK
Wtm3YuLcvHFobe17CssLdT/bpS8f9TXe0ewv9fnxx+K91sgnxHjHXxR2jMcTS8fZ
FdZNNcO0KHTtlna5l6dBtSqJMasYSQb1Ge0z4SI5lO8bc5o1927PUTbgHpYEC7xX
yjV49qMXn1Qkz/PTG+0RLMCqKXt0kDPcK6n8ciYm2KFpqXe2MJPp6mCTAACoiwgz
vp2OSdFqATGt3F41gniFLDlppfNoHx9HSzCqqdeWkb4kjXMtJ1Lu8dVgOar94Z0S
3scAQu8ygz06N5ws0M1N4NMhcOxA/Mtpd8ATJwBA/+qo5jJT+BsxohnIjoo61hfH
AdSWLdPGA/KVEWdEmUywXYIhyHnZ79TJPlfR4yLknkIhph2yDbyjQtlAI+HquxPB
MUFnZ5j5oYe01DdThElWOFte727wXMrvcR2lpFD8wWh4ZQr/P5NGAND9vFnPJ0hN
0fjpg3wDKeJXcXScxauhCXTa2ho5aTsxd1pgc2L0i/68gBKI/H81sCdJznIrOXew
eG3Auc1e+MDL28Diomk/elvhFlhtfzVG8kKDsOFcPSXdjo8NlvJfOIPmE3YtfxkH
UTuXmp+RVc9Ybd9ZfgFcr4m//SDVq8mg2YybAXdlQ81qGdWHp3rqOzLnMegJiS6K
R+/oGlgBi4lDd7Q98DX+Upn5U1uEd6TePGR0n+mXfsuPHe48DYHCrOn4GdgL8Z3K
Nf87fqTeItLSQ7dFis5V4jI/UqRVVCB7lzqPq29tgha0VwctrlWebk87NM3605bF
SXTxIWgwmj39qO74gSXXozaF+f3UfeEs+ryf70ebHPvDcB422WAqlMcKLOisR2iD
yTj+QgoAp0A+h5TC7cflNxlOnG/Pu+EIgGWxXwU/A4Xz+d15sDYjVs/QAVQj2miO
cYqpvEesJVBiAD8ELsUKMIMZmF1zBi/NJIjK/sVZ6p1TKfTZmksiAjheb8aMAK3B
thAf9L/NlyeFZor9DuBcErtLFSv9ivjZhOCDnRHIJoRhQDCEvnct1LlmwlarzcVv
NQGEoQF7z0k3stKWwR7wOJ64B+3oHRE/fa3RGH7JYvtfW4edlpRg3uUuy5oECxDX
o0mHKOEGmKK0OXL/2yoqw9x8u01nJaaS5/ONNjW7xOTs76OU2HiojcLO3RMS5Bwy
v20fVhO07a7nvI7CbfIyXBKZilN3vQwTFmvwfkyb1vajUEpj8SnwJhJYz2eYO8i6
Bx3yBZsX9eo3N09Q9hsMg0XcVjP6yRXb0swKxFfnKH38Ml38u+UTyq6Ecvr789sN
aqt3YmXcCg+4BzjWhpkXXPZENvQAtKtnpIEqMIoE6g4LA7BzWnZhp4HmWDAxTDSC
KnaMl/mV7phKfmfP1kuG+ugWkEbwZeSfENRnd0q7QBlK8AngFzLNadqyX6t6+lvJ
OfKp0XzkLTzoJiS4RgWbxI1jnfSaSWCvhQ93SBbXQSEIC092sIFodA8TXlcn/GtM
j8ixAuKlmBT9gupGL7V5iOhEXhtpbQO8mcs7qDuD0oYILLWn3cEG2VnajQ77Pm7Q
UtjY4qH3iW/oFTBKxo/SezZxVgtaAH7yEXlCtR19HwelwkEOyNdKLb372CZVwk6S
vylpXSCai7paUtKlqLBCVQPUWgQPJJ+8DkjN9dlOus66cKgfQC8LuNLhwB4YUdtA
9gTNToDAO3eRYS0TmcPNtCNYGgIOg6khjHxLYGFKq6EOdR5dR326IyF8KRC7fR6t
X7IYQJJsDCiQIZuKmmzVC9v2G3i41sLIgRdrXo+sqYthPAbBE5q0koZxYF+5Qv4J
7r++QhCs6G+CzON2jXnaBDzv/yDmBdL7ZIzDUMUst4VVkSR2R8uwlqlRgdIxPkfp
f+2+2xdG30RD57744vOzCZS7pb72b0zXzdGt0tlu/ca8ormo0YbVegH6mPuJlT38
t2CpWZKtAvO4sizuJgAFLKcYGUgcFfQBkH8HCwjeEtjorgtYPGtqmIXxN2CBUF2p
6R84Icp0b7Gufbksb3cLUoaUGO3dy2Yj4RDmaPFLNZNFcjQPEpFUwljP0LY3l4/o
w3yqlbf3UJ1C1C0BunLL72UzCtXlB2+/13aXrgF05z5CFHExXTAd20YjI6J6NAfg
YqQkGKapv/jm253xeHsHC1iiz+gNc+vseGWLHbb1K/7fupvwrRuPqi/AXB92f9pA
nujbcDW8wMommjgIBOX3hZm6l1pgNiv/2dhwMNiA7qpWIQjTrmw+RkZFcSlFTMm6
HN52AjQwMfPzRSIDlnjdyvFm0QmEXt9Cn3EYQB+SxWj4pp5ta4S81j5Rf/dLdb+B
8/D57P0Q+bb/wIEP3fTKGhAB3teg0eSvCHU1Jzv8bd+kMYvMr2e9udeT63jSwRlB
D1sufAKjwnXAIwSP0x4qY1m0L/vs7/Vxz1E23V/8UuQnceoeWupw08zpVhSNLCCL
A2KcrEOCBGEN4yRCRXq8WU2rMmlPN2ZJbojSYJJw0oQ+FSHPKcV3uAF3aPB7A9BL
WsYAxPWGKwhLWmBIUQCqn3P038ms+vh742BBEDMY+XoSe43ObwLUotni81gVupmn
P2va2zMMnYrNCuso7lOaXqqm18Q0YA+nLiSLflcc/Mc+msIlRt8PuoPuoxmPZFJl
tDVaXz3sTKaNl4e21c+AQrCuDu3FUiq6MnrG/2SYkkOTj+bzk+srdCvOJBraZPUr
qBGR2TYPnRLLDh5vbX+VeSCZrHgdzSN9NHcezsUDvmarBFlkvkpAoJxrYz3WgcGb
35V1MOhsJKiQepF7r1yjy/dAC0YdfNGLn80t9DVWFe7XyU9vkKih4KWtWZnchcFt
3f1anyT8MIjV7RFuNJAWhwvjOJGncFye8RDwUU8ciQ/NGpAyF9zoLpjbI+uGFjxN
dCNqZM3pUQ0ciWtmgXw/97rfeZBquNbJVxxj4cEj3LbEI8KNGqf3T8co3WjySB3n
kzGLQRCdASJ0KgSz5gwy6bIGf2Bk1QjwR5AT5TR7HZVVYxTxf336ynw31UlQEpdn
EhsZeC3sQxbJ+vTlUMii5/2vZQbbMLv1kq9Ukcer515711MMORb1G+fNfxfOntPU
pHea1mUctqc5PgQp/AjatbCjoRndmKJi/CZonfh168KvT00eHomKwFLl/eKlARyR
la5u3x6jDx+9kOejsA+LPzC22gp5/txv/Gvuf25ra/5yl6+LBElLKHgsptvk05cJ
gXEkg2Iutit6/hMWXWNxbBbLppJ7WBCgyPnnKE/8WE1hQhJI426R6A1j0exTNGrO
NN1hTDCkP/b3BBMSEa216MOjBdZN7W8FrpowPvsbQIpeMtS4x9FxyS6tv9e3IiYW
w7973Jykk9CJnqGFrVM3EXfg7pQG8Kex318qLGF9Lbak48T3aUkJcQ3EG3suV13s
2ccW7PZvnNfbblDfh/qafAcZSOvtJ4rrXOPIlpvB7FT1SQ/Tk7AsV0ADZOwzZe++
9jlJTKkfVVcBReHkdjd3He243CNdd2MEoZJ+9r4wbL/+2wwD2tH9OsWtR6wp9qoC
Al7bkXWzfeTlxRS7nqlmuunGwdCuXOqr070eKOPWr3puD1ie/t9J2zm2lQqGJ4TI
B1c40cljgJ2GDSQbIExzHrlm3pt1iaCJhhM56fdDw/aXVQUShmRQyFhXH9tZoP/c
5wYhA0AJEYpKDf8MXc3c8E0SUnXDwApB5wnGlAXSL8cDCiV9mR7D2aPbD41EZVWg
Dx7HHfKFeGPRDX3MmFaG7EoDj3kEA9h1LbMJjUhgfCN9tuGse3dqvSeHdHnn6fOm
OXhtMuuhSpXVehTS1qHiL6ZsQvtuodHo6xHsod8vl6sVe0EZdBvDiiLcuBJRU3+M
cvJHZkivPEVjE7ET1Ga+IGtExI6nx7HrupwwESAg3QorsxJ4V3+aVHpIaMwu1xMw
hamVTJ3DDtBvcXmrXw4H/1xmgoQCJk6TUFIQdH70czJXbWH+Y56+QeJyxyma7gXy
z+Tk3d2d03TUNOV7TbvConyBzfWWUrh1ns8zoFvRw0lNp1gjwMrU6en7i/gGUG1W
uX54lQ3YCbsIcw/PRlD6GmHqBeoaL/HZyLf787GuAUgnXfWiH4wfVkyixpIsY6u8
n9lQcrlS64bPaJOfFI8l+m+drz+/rh9JYV+MrrDkCrk1yOo1XTZ9LJjvxTGmtji+
vfUr3b/ttuJqiD8LAHp6Me2hb66OY7OoZz9XOx7C7+WEcXrUsaLdyDC/bXmzPaP2
q+1KwmpOCyDquRKSkMN8T45GOBpPDLRkvNa1yfBdoSrVfcFbb9CI0ukrZbr5d3qw
m4MdSj44ziD/4uRNAag7CjFJJ1R2cmI0B5QHVY+PYPgLIKMMJ2KFmeiSo2u/JPFW
SEINlCDl2N1zA7H/+aqtjuhXmF2bQbkwrtTJbCY7JErRXnqjH1L9+OceMxhUZ/eX
u9E466eSg4Hbd1+a6E4ORkNkiMoox2RXyQghw1G6ogjiSs04TkrWGx7Nlm/+eEbZ
Ai95m1CI1K1BwFCgalO73hlCMvNokiIyLfLfteaag0MbpK1AB7bg0euAPZ9TXJsG
1pYHMNSa/gAhSEPszxc5MxdzC6vojDaBusSQk7t+lnhfwBHAq7eaT9DRTtaeNJ/f
LnGlvXtNdqwvaxYGH8okVT7EPd/ZVd9sbFZl98glBBh01kJt1PDqDcgg8nRPgelV
WFIIYsDolYOE/U4boaPBe/sFzrFwSpWv9YqucMlS0c+7wFgrUop0QVB1J/vwWtpf
DPexOH9YVpB0Xi3R1jJn8zJSyyG8NK4IiuUljFrnv95Z1dHQ62mECTj3J9wOISQK
hjqbMTsKdlhMBqFVluf2l3JD+FsnXf/UujZcwxZDe5MRL0iYwBZys1AXEuFTsuhP
b6TgZmEvN2/x2s1RgRQSJ9hxHiICy5izJb5Xyu7swNuUbnALi6NaCAlT5A3223TN
uiKHTKTDF8r06yDapDOwKiyvazyUbd7H2sX/4ILedhNwvFa6Hf3mNlXEUb6MmdKX
5VqhwZ+nB9BS08xTXkTxC7XKYiPKRQktmQLefBNsg3TfKOdBh72MULwGShXtQ8U0
I6E4lBQZ1zwHTBAYQD76JPHlUK4qPd5Bkr7laceGncuN28Q0qOSJfLvxDJzCV1hZ
0PqwX2GnJMwpgbm0Z/jfEGJ9YBlm2TTpUnzK5KMq8Aa7LhbcIx7SG6Rf7cUE95p1
gT1V4BwnDYSoowcikVkbhRYmM+dSCHPB7IIXJA2+o1A1VN/OK0Cuhvyc5AUj0aGr
31DVtXHBUH8B7AlRh2mBxRRIsjWB0HhmAAjCgbcO1VKPz9rFpYaERW0WwOkHtxy8
cW/oRswaRmJE/xRb2v0CzbB4Xm3fVE9QRKacKE+cFnRNe7DCBWyTxW9NAdPWx1Rp
rj15FSVhVtR0PeA4wD0etzB7xm8nyvzjQWAti3KB4SJWMMhLv41fRw7+0JGWahYr
59ZaT09ZiAztxcY97pG+XW7z7Ruot31kazwoSOhHVhzR5HlSVwdWTEui6s0bAxO5
Q3rV43AbI9jETs6qOiJnxL6eZkkYUvEP3CBARxfVW+af9Iq+SHlxIPrs80FYSEJK
fA5qEF4NaeJozB5JIxvzjOXMQOO3bToXXm3OC7PPcn7SpkUB3Q044OryhA1x2jTk
6Vnv2bOAkY7yfEyp2x3j1lj9dfb9pTSREjFaQMAK9urxNcYiOpuIDdAq/BFeTBRD
LqYo/EUN/wQ625wK/Ohd7Q5ocdwzGrOayhYavW+xr6OIOg78RLoiyJjlN9yVeAbx
C3CXh28AzxPt2iPhy6hSJkTAuGL3tBDSXul/NCb5PqtLalJjWbd4h5rnclZwv0u8
d4vFcZ2xHzhuIVq9kSL9kwJro1Anboo8XFUM/E7Oieaqe4t7aAS0u07Av5KLH+IM
rnMBy6wNqLF1fQq3BRoOGakVMO5R1qgimBCYEc7LZR/g+AkgqhoghQlR/jZ5qOZ7
VmZeVAvhIxkMxzK0nbj9XK4m3eIFCTLYSYHoRSpZTsWBfsMvyAUzRqPZ4gEzYIZj
CLDm3xlsPNnqhEFpDhZjgIkPWID7Ispqa+hvk5uUqXBI3l/gR3XHhh6QQSC0FbAz
mogGgqnAD09dXCzxKen4Yd16H0rjIiO6nEqCUSXsUyIS5NTqUqRh9tprVezm3AME
vMQdZoJhOu0K4p9uOhdeqwb7tWIL5z93BUxTXSr+Qg3XgUWy0QwnF7inR8e3zO/X
rr2OckWTCVoowtuESyRNIhYKOAM3B8vf71GX4NMbR8Vbf5URlYVAFdA+rTb+mrhC
sGUsZ0+diSqR/ktubTJWpzXJiHMn2sXdlprDD64/HQgaW8YsLci0JqmjS/cTJh/u
YdxvsXWYsjrs5QirDIItklcgZ1Og5SEYOTt9E8kmwyA6kbSaxNbXo5cjtINOyV6B
sM5Hv1hqaiW32W1h2G0oIXxwf/mvqBCn+1AD8hn3H95kW/V91zFY14z3FSRjLfqN
hv9JmhLtdWr+hFO5UP/ErIEUiCzdKzk/Gp4+J18w0pGzt9j2QFZz/om5BVJsd8oY
IHT7Z2hycd2Kz2PaD0GHcl0tXOTIn2CCQYG8dgtm39+4D2IVIsKawscDodMlLI4e
acE+IM9OkW+L3cpebId5mVi6d0VM6d7hGxsphXWTza2LzJBu/WwVI+6ZA9x7T2wY
QBz00d9prZBqCtE0nbm+/gwKyHDo+QyF0Uyz461sEnXD8RKlNOHNWN/bbvS9xZjI
fUz33Oq7rnzFcJoxgWSj3QlN/ku3PMpL4QK6sTT1113KJpGef7e2M0gr36oIxWU0
sSslIhAX66UGkDHHhk1oMflmZcXGPF4HhNODjavM9lrxJ8OhnJdYnrSBj2kTV4eR
EIhkDqK0uhCidGOKqFpslGYpJzyVAGRhvrzDz3/Gho4jX6/bhTTDeif2QfkyCu/V
RQgKxpcU2H3oW0Mzw7H7LLNeUbGwv+/+oZCDZ7jd6rJQI54oa4uCFfMxGO+nXb9k
t+ywG6qNGRnVhtGHMq9tytBY9uKZubsnynAEMbBoEKXxhqvAK/x8X0kqyLL8n5yb
9S1/KtjqXjUSRqMzJ2LNv5OTGNP2/oJDJ3DX1fz54lmZBgqX9VuaQj42OqPcjR1K
J46iuRe0A5/WYKmnsnkZUcvZD3++TAphF4bbL5PjKozgpaVWapT/LAn+1ikgdvoI
i4H9SBDcVcrO1FRz4gCk/k1q5opdt0ezaBFsJGBomwd8JeQOnsaeP0XSEwo7z3Yb
lkOzu24uCezIsPjgzsINTeenxzNaE5Z49qcHKXvz8NRpTdoIQQiiPMX5OtM+RfE+
m+8d++sAS7BW+2mCkF9HQETT0WD5K9b+NNDJxsfHHaHuesicJ8C580p5R8ZHtz5H
K3J89zFDbhFwAwj0QHeyHcwZBiMYiX8BZj3AWD6TdJswgD2vENhDpC0LEWlyOm52
VOpeYh6yTMplYNj2o/29xh2dCBjkAfZz6Q19C20bNP/Aj6vKMUVWRNUge0IMKT4V
mFFJP+DKnBaAISv/1fqhGMkb1/wDE4c6xHv6V21JKrTkne8kP716XZLya6h3Hn+z
vBpYQ87YOrh8l0d5SOxZcAzB2zvhvBIQmWzIgiaHd9ypz7iB+1KMV8sH3F7XCJzk
z2XSG4RrKNxaA9uEjxBlxdvNHle70ZX8cjCXZJ6r4wbl8yE5Xmy8n+zZF6oYShVd
xKae02DqkxbsfCPIfhfZfjdzzylpAeh8tj4uF1P9/4L7Jhv4bXQ0LD0pGu/wwQrR
9T14lrIDkdVV1IvxxfxpXKgWX6ip3xNm93ljF2IzHG3T4MAw24hpPqGnNoWlekAk
p9LvCbtVRVTBgQxgogc1dDe5Hv6EB1ghvDuWUuserObiz8edYhhv3HfTdRz4UlMG
7nLtLDc89MltT+Gz9++HI0u4GHSpiqv9SZmL6TuZBj7iwFm5sk63sD5vKPO7jm7p
wpm9CDpTrOZ6aKisziygPRPluEWqxWP/lhHkUCC6lqtSboet/hcCPfzUO+eQ6yo7
RbGB4dcUpcuOZYJ/8GzZPj2YzrvA+hiXkPrCELrSbj9VcwqUuOmqA6KSBJW7A0z9
f2hGuoZTRdWWeuCWDMw0ozUOhJURwAHxRtqAebYQj0NZAVWvsCw/nEEZOeZPln5W
vb/g3kTafqhQIdfDshhoXfqgch6XTtJPXnybkCsqqUlUuP2baBI1Ya6aHfg5p8B9
IEYjHU/mfkWW+ZmCNm2LEJX5qHj84Q5H2DDhB65ii1IK8J96RNn3uo9XdcE/1079
isflDz3I4AnR9Ir9Q1iYfGib0bCLx0ELyJrNCGYdnIF1ocY1n7BQPW6XoF3VpX2m
EivuUHdw6/xPVLjp98tY6ptH98LBjcrABTm1qix3Gz8aEPNur0mfL9+TRibW+t8K
apw1SZ1XWL36djlO5Objpoj4c/htTM5T3MxOXg26IWFmMbE3E8Sk4lGy28kLhH8p
k/9VmOg6waXLYFN7PLLelc3jhPPgHiSbtxKy0cXVSXE3Bk15clYs6QyfglA0D3vv
UwUvR8fkG/x9FnVbRehH3ndUyEdslKs7oORVtRmJkfpyVN9nacdeLb1mt7jJTstp
18xvhQlqSncufOrt9+yZ15XhPnLeRPg9Eq8MT9nbkIyPIMRtbr37qqLKlshg96HN
s9r/VateD8SnzA+wCN/WuPe5Jj116ukwHT7bdgYaMKtE47aj/Q5MuqPuYycBiVNy
01yERuidvFPDvPcJKg0tH7r+wkwAZd5kzlq5QA9xs3FFZFb/SF5iYbd8TzelY9Ob
KDwpO/OO4tz7V2lVWBQ41pf2RoVAUgEBp8w1ADeMjKLVCOyNsqAgfOJFJnoLQgM+
rNiA8YYdzoAMiV6EDKklmVhDcioxAj9UxFcRUu/6QtOyiMYEfBLKF34hO7fYenR9
IUR2k/CwfAblHlgXJXBvN4ClEk73CDd8cMvmeHizaLba9Fwc9bYLFgZtslPqLx3i
ZrnHW6zc+pt4OH73ZJ+MB/xqcYbpKvxkXFO1UK41e25XEdivpKPQOUyRgH2MStHF
bQJuUhTP8Ba2LcX1TqJ+pNj1vfO6lM99w/LL9QyT3tH3ButFi7SCjWgE76VdReHF
macbqChNLKngYBF3gdqNGpFmNkmesQHu0sDq/Sh71O2RlYQubsl78hj47XwnRo/E
WSx7G/xG//+5cyHREq2B3N5gRjOI0c7+iFM8Neuw3QSftzDGW9sch2yiTEjRHok8
LFbICwS+gzlnMemfQyG+ldq2qzFt7fiNyVb3hbwwJezpPaFrZkY7qx/rGPOQy397
rExpSpxpFTWD+BAgLRf1PsOxcRRtzgVffgl/woTntBvIOSAtQJGeA2B1KmCI5TjJ
uMJ2B1dwcHH70LEzKElQNDbjy+0IViQj2SOt4iEE6emzQJk2IxAj9F3EcGEAm40m
WsHy0ky/gLR5lWZer07gITdcNu+SiH7/p5JUm4VtD+/hYOsA1IuMXd15X4Ewb6oL
X/AkPb4k6Fea9ZafIxk/ym7IVJbiyBuQKiCJbO6u+UtAsfEViv3sLTTx5CYz+lms
i1pvknzBqhRC3rJyBWEAKf5VEsunCWO4z1Ifw18VYubKXv2vihb2Y59qYOmmgpKp
vZSHmj3oCKDA4sgGMXDjWmvihg0q37KCV1iuQXAMt+UBd4edrD1sARu2wGwJchJk
SyLYnv3FYYeWR6YsagF4m0fNyvh6/pyYglzfjT7BrMjQX6ACzlKeUTmQJi3pcLb9
/iXeNCwGJ1t1vpBly25NPITFt2BdBj51hDBTeOmMtqk93WavkDnpoM2GfZ1Kz5KQ
3Ww9Mw5hR4f22PjyxQpOuaO2A5Mdfom9U1hb66EZAP4Lh458KREKEM5p4AXfPGn0
Sn+vWk7DZezuABbJ2HC0H2E33fgn623pKjCLsCGxTYyy9OZvO0Y/L9W8nEc4jtMO
XrJNxMqdDP/ozzdp0QLbCB7502Agyv4s9U8JxweLpMQZIRGVHMT5NU6/K9aqoFYM
IcNBs2Xri0+wnt+BmuVl6mmFisThvUeCl9G7TCQIxYx5EiW0VgRnv5755YAWy1X/
V5Oec6G4NTtB9VZkeYqqeHRAkKOsdDUmQIT1K+I5wQvBGjOos+OE2fQEyEw7HW93
XGz5TMtt2PmNf8is+bY0C8esyX9dYqR9xZvC6ggJOCLMXR9spGyRZYmA55YX9taR
cvM07hRlQt2nQjmp/4PerfMoVTXBz+3p6XpIE2v6y0+PnOoQ99fheGLgBgSX0N7Z
lIv0X36sae1WvsOhBNoKitZJUtrvKk22dVQGgddSh2lnOQ0P3072ohoNNS3/5fG6
hmZoL+YXShn6YEj+Mzly1jBLgvYpUSPUuiEmF2To8UU/FKIiiKLCizZkv3iz8EPR
YqloMj7cLJ7KL7faDUIft7lHOrxfcgeAaXP7/rH1u8pObF6YQVS+lws11VrWCsWg
uparc/5SA53O85ihPocpr9pnb4nD495PbaY8mBFtbHH1IDSIRLT9ZgshkcZpf1GB
spoikyn9u+5vX+cBZLDqZatxN85ul4R7RCk+bgRpV8mfDNXREKcr0e5xx0KwzH9P
bnu5rsZgfCQMqFIKQwhidkbCNssOyxk0FfxTo7o71wh0bJP/AlyBsZSrJTRsTFW/
5luULjOYNGXl+17BT3PhHlQbmb3Qj3qEyNnmh3m6JGSlVIzFOIYDa9QSqUfnJRNl
srRAu2I3LIJqrIThbnCMIZhRb5ktbjQANO4w2YY3IhfDdLIyqDq1JxpJS3OEYSmF
DmPi0inOMkel+5SE750YQ4cEj1ZjsxupndNMjCGcXsiT3Xjj54ojuV7lwvh0y+mO
smjcf1Sba99nOzI4jDok5VKsAlc2M1+BaUga2VWGAMV8iDaUaXBJaMs1qrhDhLO8
TCLyCvsXIfA5+DnJnYo8Sx/3HQnVcqucVwN8u6k5b+388EASs+qHw9pb9PRWbfG6
WDKZTb8SXiqsMVTpFySDv1rkA2MiomSxP5049uSoCNtm59uDpKruE3eTT8IJWyVq
1GvfODzQLeTtpnPsaP+jJV7vkk3FUARFC63G90saLIhTgGIrnXxXyh+0xVIMl/rF
Yo39bqjnY3ze4QsV1MlJjPAQj2MoAM/wrqbkIMIp4knkQyjdCDoKwFFpZK7HWMTp
au93G4g3ooVqGJo8IaKTZS0m7aBsMp+NgXSPu25Sc9Divrf6tLiOLCckyzHFIKXw
eKEclsx3xvkKOty2I+xIcVla4xcdYrqGTU/aq3uRX2AEdJ/X65COqvn2Gkrxgjcy
3hYQAFCu7gCJLEyX071WCUdYK/YzfSRUWCmKG/uKS5LLayCKHroBuDL8mlfNB7SI
JEQCoajp54HYKlt6hU7Lu05KFcwBx0KJWPG9q+tij9d4TjPWJQCfaab2H8Ys3cbL
f6QwAd5gRkI6URjzAf1wfeKSx1BIv0o8ummhF0dJQ3L8ejFm+2bsKeUR+k6m7pwy
JlQ3P93jY8jX7EbiiyTAQ0JIw2d5pc2D/8iXPM05nHSRTpHX4idFFlBiprKrk+P/
lx2MlAT6wO85fcW1ofw+hI7rA2j2z5N8F7RyegMvezlvFyMTonlKXmi6V1PctMbu
uL0vajtqEDRZV1ZjW7EiQIb/C4iKTdznHeX+RfLmH5vvoYtkXS2yeNfZsKGjYMFI
FbZLStBmNRpUEFA2bVN1TKIzlOwQT4gnBrcZLD47BAiH08SuuOE6Z7zYdZCNRVjU
RSPyJX5CtI6UQukAnmba6WQGvVSCsn+Ppuag6fPYmaNL40dYeiPKODP/5ISHZadi
IBD7Bbw5jeBPJypGjLf0xAOOVMUqWm43gWlB69oqIB7Z2t6pGeJTW6Li2drF4jD2
Y9O3gwGqveKX25QFQfoGh3gGNVAQ4Lp6FdH4F4hFh2eYbQwYv8IJidCLY161P3Nv
KcbcG8LYK0ikihFtpo/unTga2PZ8QxOLgR3qQv7mWDqDX7vbcLHOVuywOVNJh/yY
z3xZZOV/hTaMMy2H0XUAJD+QWxv95KyusEW3FnnJFUTxFJHQxxZDrsDPWcwZ32aQ
sdh7isefXAS9jyjYncQynLSRQPnr1BKe2ILgO70NAeto+q5tGPP8HjYflYobabxT
4TVGkejfUgxir8W/VIABhsRvQTOjT92PJD80r5Jmy9yn7XtqR62cmLW2QNLdN9nv
6HT9T4l9rynmVpwusn2KI/d8VJWYzKK7qeFbGjn+YhmQbdVTfCB5Xmgtv8qaoRrl
pNtGV9T5MpqMCi7yna3Itzmw3eEay+qa8maByiLMLCfJaK6gfbvy72RsLzUy7ce8
woiXyob5GoBIOOXTnT9OvbxzsdvlS1HUi5kKDgsmnujX4DKI+GRNOQGrUw47B3MS
NEywokCJ1VizAGRVzEJPXA2uJNC/8zGHrNQ0PtOB5Bie+mbr3wASeZtLeOL9QAL9
6PMnbTAGPZRUYtLZX0/nJnXcNYPjtgLvNwVYDsPz+R7CG+wPipnFtqqNsKThazdu
E5ajx1AofxEKD/+oqept9JmoQoWRU9IvLq7gmChvLUzU1hEqMZyQfCBDjdxlPGc5
3hOMtv3IVW3LyivNLGPAX/r/GPLKBp7BFsqpJtT9wFmjYqd0qbEzuvlC4PiUGgJ1
MrCC7cgPVbj+CkXyTOCYyefO3EpDl5WnCIriA9O5XteLnzLyspQQ/WLgHYC+o80G
KCoKcYrutO0hAHhPOFWxA7LxpdEM6n0iUB0EPuVmeZTIYz9DEYQ6yDbKn71s/n01
G35G74ofv3zKwB4/1AzMAsC7xDUo4Q2QvfBLh1/G/f7wCZSMVJ3IK4HfaYYyRKBk
/52Lg7uAgbtXMcEkqXtCPx6na6kq3TBRAWHBycAP3ePKrIeFYHpD6dWUOKGYlZn3
KSK/tliNZ8bDGYUyPCWSLDCDNYm7qUv4YLwcLnA5FLBG8jg3jRO+V9a8Jg5DrKHv
/7emRsHpUlob/OdMweV62aqEX02gfR429lPDksVA9lZjwFJBPBgculyq7DLvSBMp
YwKjl4uJDRsEz7or+UtX+kwUMtpiaYUAS7zYq0/dQMR905dcTUJTkJYI5fZfp+ZR
ZJS7cPRK6UhCVpNTGNZwfhgG8cWMpCkWNM6tjFrs8K+RvHRTXGmh0T++YlyMkq7M
n8zRVkZGdeCZzqgAqw5mwp9XatpGfP+FuWJKphyGUahsiyxxCPoKYensViP0ENV4
8VhvJBHIPBhqB5eE0METHem+QE0f5oVuhBo3HCgzFSKrHouzL5NoGL6/Kplumd3S
v+2DLp5DvvbzXZ+bpat55eVFfwqoDvP/DnLfaWdWH2G7pamyRkE0F7p3V2MgzCin
2v55mG0Cdjea9dPiHjitcn/uCq5zXUV2oqofJLM1foci+//SuOmm9hB2OpskSKIf
mgVsmOzmXKqdfq9lqVbarJKCaNfv5IDyms+FgVDFgp3RBq8ixN54elFHb0TvR59d
0lDlyGQq86JtqIVYzj8q8Ww3qZJHIQiHPGZbgZiCq6Agn+ZxzLPfWOV/mFbceS9Q
jLYVgWftYJTE7f4BSb/Yxy2K0Ezn20Mts6C2SswF0ussjLAzou9wKvEmSt128m7x
ONhAxmw2dvPKxDrfEPEv0NAF2XTIqVakQGqa7xaXR0yn9vp6I8eAy9Z8fGlASbsY
/RDm3kF1T3MQnf9LkerTHP8zywsPsQi0l7zNZ1Cchbw2xsZuvT4YFHN2gm4TOCvS
vFnE+V2JoC2cW6FGBDI82wqONuExrjznxTEnqEpCib0yEDY7TAhlqjqlRDXMQUjv
YIyrNNdlUgIvxxvGQecGsL68I+IL8ptNLxagjQbMtYTDlM1MyO3epXTaKjuKcqKo
660Yuo97dG5heixQZYxCUXpghXXglxva1bD0Pek4dGtCwhRRB8ettU8Cx1/HcVb6
NCY5FUv2iI/pZBSsnHAukMKIx+zdNEf1eE6gc1nWrXCXYq72cmSocEU/3hziXPaH
AXJ9lVbBJO0BLSeHfW569SxBZE8e33PovZ4yQcDjx2knah6AXhF6WXItX8FpXPjo
uVPx1i8Y8IJORQF2UQh/q1PNgR7zBozjnr15dhQLJcHRjrML0DsO+WdoHDfugBgm
OTO4WctR73O17bdVQ5rjtdC8DM3cVh6Mx5Pa7fYQJd1g+kkHRq+l0VCxMA3MMAiM
gEHGLJ8IW2Pgr+7kvD+uT9fv+S7Ez8fNux99HCQkq43k56nG6nx0Te/bssPbcWEH
uB/ty/HXMg3AjcmZ3Uy9aGesZqDjXqJ0EbyE81VcbMyz9Md0qrj8BeUnO1hcCguN
qTYmpRYuywg973kMfC8xe0ACmA2ptbjTD4S7wCmnKeFtnmgb4p/QEiI9pP2jfOMm
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:31 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QtIkwXTuj4CP5CeZbpCphQ6yQQTKdTjw2zIfZXc/qaR064/d/Ea3fPujcVLL1Ymj
RF2N08C0N667rHkCF9FKZtDGxa6bGN675pPtqQnJe5KgHJ1miKTbK1Q1miVBLqvh
IF07YZn7kSk4FTOJoUZky/pEXQrp1yY0UAGK/AKQJQ8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7216)
cdpDKf3E14/f4jf0cEZYA6nnCTMay/9bLhjB9I3RekmSDjin7Pm44fnsikgWKU5H
qtzbTejHmKI2JJ4+P79BwJINorVqCywqF8QCDrDH6dCQyC8wy6Kc/fV0pmfIAyuF
DPY37zWMc0cxI+azYj8DmXw+Gk/JNImq3gRk3PDhHC9R1lsHg/5ZG2lGXzctx/y0
upYotWBgz3nDU4O25lwLHHNHG3JCgED1JzTIIgP40168RifkBwsSjBQNsJ3AydI4
sEx3nneWAqJkBr8xIeW2YA6rzIWUwlbBbGlPWA3j0JgfohBqeVlHrpOmIHLamRMw
531+XhYgYYM98Lsbh4gWKLwskLUBOFCupzl8/tsea0d9Dc1PHCS6EXRCov8AWgg6
F5WdXvKTFXbepZFgKTAGq4mJ+5dKzMB2JD/wv9sq0GqtMI3beaIBxfuLpB7idPTN
65bgwCqNnR4JxH0pfVouHDojWFdDSTjK5p0UONq+YAfZWwCtahHFC4CR/Rz+1zq7
7LGYkt9EtQq1MNUctNxxsXLKFnsJK/aTFjmZtWzg16LYGuvbLKe1UbY4KER+U8G4
Qm0RTmOTdskCIKsTZkyOyMmFF41iQAaSxjeaXDTV1/8Cd4rEV2UXTMiNjyactu2T
H4YIxTVQWh3pBC/2nhN76nTAmOaR3CR+rAZY+ejbIIYFcctkiEdxmSti7uR161Sn
ESpCGNR8oFyK1+6g6mkILljhWoTXi7On3/qw6WjSH+JbruQkKkAk7lYUyPho2YkN
WzsgQ1B7SiTepPITfT+QE6hEDgya9+0cEULH6DjAw2SGt1DPztkbuKbkI9dcitdM
s96V8by4Lu8DTlY3jZ0P3ZxmIkPuDhUM1BiprHqcAOxAnkLxkblUfDUn5G87v8eH
EIFm3AgmFl2oZ0mVUqCOfrT+wVuCpAo9G/T/xRVC0wGCj8Wyt24BZiEZCF9ccFLQ
Hk3uK60yA3Zt3Z1MNMC5VRFtkcQ4b3ZrlKNgxMVwP3Z2d0CcmKpIwTxR1W2v9OER
xrNHtGPoI+1A4k84AjdDXXsIIdyKGp7xKpN5vL9Sw7ba08a5wO/Dk0v6hSGKHYKX
7dAgse1nnXgsZZq1Vo41iW6jQiEDWy0W0QRO+WxHxGJr25qITs4h48Bc8Q5LKuwr
7D9TGhwe2hG8o9bvcbUokqnVFJdnMp25UxKN/SDxTXB9Vl0W48JkVh1z1NezZZA4
ecTDvgLLZ0uPhwnApBIkbvnE9HJ6BQOvU08DkE6PKCF4R8sbRO9Sv6GtU7VGejNL
gsDEan/pDPR5c/q8g3/j4BNeXdGan5OYOPvWu4SmivmhVrXrL1UY88OpnB+gwMmU
hbq6Lwbnji1yaK7SXQWRiwcHAfYxiCCt4iJKt/8I4CYaUEH6Vmg/B8GW6GAPmPSK
zqSmdL+9FzrDRFDNRPgzz2mYkWXLJKN3PAI9l26ymEE8WpraOsbTRdB++kMTvfM4
avAf9zuTz0a0kxXZEqAfmUWp9qizjhZLXxskoXzWWrLf56iyyz6DzYooWL1VRIn+
jP1ufGunO6J7o4gtSZN58dUPA2dzhm8gYwMYuPt7f3qa+Wfnai/aKpXlMPHjkiQF
HaGrs2eAuLmzlWfzTked7qIql79NJakq7dTfxxx6l7YIYdUsFokPkEwcj5z0VwCC
6Wsaex+RwC+jCqyDs4+k6stF3C/l46UwjmRW4rnSL74sBGPtGkE3jFnJkmWSjRlt
kD5gkB+sf0FlgN8s8VA0uP5MF4aVCfT0oSk21SCpAs3CczX67RLLUM6mq47B6nVb
pRC22ER23mvkVMZ8raRyxxJQrzfACnpOO2OYDN2EGijM8sFZmkoEMQfTIxnIC4ws
bvMZotK9E3b+InobL947TBTJErKatkvJXfq3zOaydGsW8gnNrfb38brwLfvRLtFS
sayAGOljphUEVn8+KmUEERdrHEmTYVTFSkBEF03eUyV8hIKWglrJG+3SdRxjrSfF
L9RcG3WyJBm351++xHfdBE2tJWSGqzFgOQ9PWu2WMgpMoi/Agg2F46Gvd5jWMrTy
iM5xLvxG7JALIf0swuMZb7bmasEbDLkyGSHmulxYRSyM8xPb7/NF6RffMb9E8S4M
5Fn+PLbaRsCvqkp7AqwCMYLtj9+FKdg40b+7Id4vbnbNCr1mvY6U+WBvcWgfFG4r
GVev1yzMv6z5HobnPmRLAKubsug5yuHlEhRMxxDB3OLE9DbJ1/aPylXanL/YXnec
O6+oRg280UKu8+naSe+CugmJqTH4KZvEAz6l8bqZAIpAW5urhZe2BwPva0infPpO
Yz5ERfQ2PdLjWAjoqucI7uTdE2M+Hy9mdtGIpeFEh3K8vpImbmoYt5jQ+XuQbj50
71NhsfXoU0mNJlEUIW84Y5IAZJ3w45UjkU7AudF40vG8uYVQB2JTxwKzfaynYhMT
9VT+l+g/8Qha49VaXPdi6umLwbxL99kf3KDi48aZ+DWJBjwiQgfalFNq1cmsHOzs
N4bFNPLCklYTgE47pp1Kh3an7toIoGJd5t8nIkPhT1katOTDzR6Mi6HprLLBxJvW
+OcpWrecJhsqqml3hN5/QJHmvWGrWqk/S1VaQCF1vTkpOoxY7eyWu6xMD9+GMXnv
sgQ6530nXVcjU1fDVFGfNiIkzqKdj6oI1H73j5pW/aAcSXhlSx4HmqHWx/ojBWwM
YXsRclMIoXcwIypAzHsS80jfLTEiVgABKr2Tw9gJCxw3YLHfO7dTe0RaQnyiuTHr
/m3J92vt/qwPhnzoawBCq2iraAOg51phDDoGfA1kTI0VSKo5Huoxvd/ShKqiTnY0
R4BhmmMojAPkNR99tqJ52GnBxR3hB00+wCJwukWEV4V/i5imuw7HaHQMazaVhekr
Ty1J54DOlqmDSKdBM8ay8GAWI5NGrE3SpyxAU+FAwcGGpzuv9c24SLAgXWxzlvIT
6Y+YEAdWqiltP2NaE9997MGrrmjKXkGyPV2AN0qrdWssGRQgLmKF0pC88Io4mFYo
bWX4KIs8ToR14ybo+8ILYn5n9Z+IlxHd1DFkhAHg7koJCDG/a2mL+gFaOc5Swnhw
e4Dp6uJvRG8YS+l43HyrrPEbD6o73C9m2rO67Q061UWSCzzougt6YxkAEa+y9/lF
+qkl1MlmpFsSVdjsRdtP9LeOMOp9hkgB2ObJ3cf0eBHOiipkTqOILBb99Kt+/Gwv
bARAYI44MJkl9K6xKKUsvNg5PZs8T9/643ktvARZZHrRUPD3I0dwmDVTD28UKbYa
+XiRP8RJYNsX9UU6+rmd/VbNFeQaAhm/CwzqOoOzsXWY5LTdVcJm2toNmFyF/+AC
DtVSfRI5IvRxYbZHKsbov6xv2WNs69Zk7V7teaps4SWc0w8GhvlXkHqaRZbWQZ9L
+gQr9CmDlZfdLk43KcxEnUHdx83SbC4XupCZ+jFHVQmrVJL/m92HsefltV/frLJ2
lysCRauKW0B8BgYHWxfMO9s9YL6uO72+kHVCrPG2CLtTGEeuI6xXFvceJtO1Pk0C
XO8dUx5TGFD9Aq37PGYeN6LjijjQKIxDzldmaNa7Ek6CMMcC+xI79OrB7Tv3E8qJ
NbHI39Cx8/ysWLqAP2OZ4an/lWfBc97zA/zbO0ow0d16ODbq7ndSlyTRPZKgao8V
yVk4seHKw5/hU23NNFGa93+FFwG74hrLlPSOc2Kn4IYqEDr4G1DziiD9EYjOQa5Z
21927KrbpGNkW0E88vk5JC+TcN8Nbw28C63fEBZrm1d5IUwcrJWrWYZIHaHZOyW0
bKZ92xuJ5YbKVon9WTgUl2eX5118y7y6uo3W2l4O0fEQQItg7OwAcvxzreFqNQH2
nEdNouORGrBs+L04qCINC2gHG9UpMAS2EoIU15/2aOhMol4jxCZFZw+bpWMxZXlP
xXg/iabA5HGQsb+mBUYO3q2BBOuWUV5REtV+tRsY1PsvStTXlAe8x18Dp0s9K9qn
Tgz+Do4kaPDUhANloFmZ0PWfRdLOY6qDFPsh1UXjKGXLQbNWlR6u5aqjFrDlZVvf
y4Du+Rp5gnWqcBD/FC+Vi0wwz/AJEipk8IDspMU/1dWAJ/O93ZuojyUgXMftekTt
BtYxXRrIzYPZIC8LAquc9Y/chnzokB6bJRq/EbSWWaQVklFkjsgAUb7zKKSX238b
LJKRXISLqpY3KrF5xQwC2Xzv6l517L0tEcqOQXHL865KBok8ecrFGlRBABU89uF2
I1CQyNjmoN9QGG75qD/grfCniMtG7EX2IK8doVkBEk1fOMqtWVikOuzVfmPJ4Pek
F4oJFGJZgRl/dWA8fP6uMhdPTAgpDggtRtVRDco7SP1n4EOJDQRszmnP3xaNLqXZ
1PwzGArf7TySXvOzOuXlRj14imjfrEH8HMUj0o8hdbnkJ1Sp9YYGghN+H0br5SDe
eU/5nTWAhUtZOn9LEArEmc98m+GaVv4MxR0pitIelBOe9ruNWQs51q7XJ8zqSBLu
4gh4l67kzKJ+XLEWLwoElQJVrCKZhHz/IqqIDhY5hRt51jjreUtCY/0nwGc9Ovcc
EoyK0kSLC22RIA5z2QBr7dSlaxWeDX1ckdqKUziwdInZjaQfmf2/G7abGUnSEnf+
L8Rzu5XU/GZqKHA6na6Jd67ax6829+JptnfuSnbdft1081IncIAUSVTYGE0WMOg2
7zM5Taa8TMUrP42xexGHjsFJFXF1VKCnsnxrMD2Wso+Wfr2igVfTmbftX/MAaKXd
sG1Cfu4jDhI3gnPwJ2OgE07Rm9nDliluS5fcVVklHwsaHP4lzet3T9Dfli6QQ4t0
RnJ4ImTMPqHhf1kNrrE33DLlT4PiURRro3GJa7mpixJ0Lzk7IZZScoNtWNQrJj9l
Mb9wbZovXR0r05ykg4ErE1loCFjQ19V/0Vx8O5wkTozNAFq/7WC87g+/8i+d1IeN
yMpCNJvELlaw2Ys+3MBQHWijvzYvoE1nBV2ZXYtUWGDy5TgwNuJkzLYUt2S9NCXm
9U3iADet7n9oCz5cXON1Z0HSoP98FNjfpEDL3f81dCVW+Be2MtCyZOIfYZidpLiB
kxkPphCIqSkDODRqaTN/peCUptB/527tQwRBY7V1n0Q5XR2b0mcfCcoxpSiGaubb
RZnWDpFu9En7Zx1+wItK4w5kne5tfaDlcV7iyzlS2OYvXTpcYUO6STmNesDUyVSc
wreQxaJZMO/2scSZSPkgwOeFvb5tfQqoPCy/kUrb5Mf1PJ+2kjjE9RxYXccVGMfc
Ud6rljK1c9CamxHgY9glj1ebLtf+jL1908aNYyXvkhz+f7zzQpWHEpzq1vPRmciO
SX6ZeEQZEBmMXOstd7TCE+xqNuup39ebwEel0ir4zlb1WKbh82n2CaQjDmOP/w62
EQqcwTUEDgCUy1VzJbHNf8AosXWLUKuKVEaMj05CLGiNiSevzxGuA4DE2biGAAbO
5QWcbYNY/C+B0MhH9IoOhmaLuqciCbB/DE/pLRk1o50qf373hrn8hGqAIC6mlSKf
6W0PKI/RkgK6Z/+3gtqAsn5I7WOikxSkl213gVdIgKPoQBgMtPbHXJVDcSVX3rfa
8F0FFJJs6zpU606d6ccGHgZxRcSj2sm1wC6WKiCsspS8bKQHt4GnukxrBfRBC9Ex
z9aEoRtSIYRASWhIelYqOlxeoX4V8K4Zc/hx98f1QpsIiGDAUNXY5RcEOAluWrdT
a1vxEm3pu+KScqS86otuDEI6VyRQGXKVxD7XRKXGQRjrLEJswAhuqWqPS7TKZLDH
Azso57+yjE3iD/gubYbrWA3CXWkNIO71spq0wx9ISFfBYU1MEBjv4BrQNIrgSzMA
KhzOwvg/EaEgZYpv9TYzNz0EPMeSHXdurHfNvVZXWao2GwCqb0QoquDEvjhv3M3x
obzor5MNMbpdgk2a0sib0GaCCoSMBD+uqRaqbtLIvLex4gBsnw65rklloek8D4Ho
k4hwdLQLL0HUS/cjkRZvZ/GQM3Wd2RnKTJWrBrV4UPmUSztPua8xsKbDnujihKQC
Y57Tih+iq1l9nhL9CvHX/bpPQE6GsAX2nB7PppLqvwvvpTSqnF5cf8ElXvDFoR5P
jicieQu7PQLEpqfBLdh2zLF+OPsctBb75jL59utkNhRWrhINPbAiQMupr+VFL76Y
te4GgWEYzfOkIcXP5qqLYksl9wNShK5Sk06NXX5y1xtZF2ZMxAqWq/fD0PyvMLiE
1WKqlG2oHn0pWHUCHVqeYyGDyaax5rDDYF2HpY4HiF04UEV61rB6zKHI2PuP3+z+
2g0G58iRG3RZKfeyILhJW6WX83a3l+Nbk4y0w5oFpNZs394HefuIbOkvOaDe6uQh
P2BpSD5gvQ2mLWqDKDmO7Q/VUQfvfvYbm32I2kFeDXOV7lkypcuqHLWmVZ7RwwBT
rBPYoe/C05f78aEzCAGFO4cwBvXFL7ybKcDokjEFkSuEZY0z+VPAg2IU9gMqfh++
CaTkve4dny7H9c+DwTomzeY32Qf1XQ4Eo2bfUm3wFq3cZ4FhLB8o9rTxIdrm0PPP
VRoKqK/CvWo9UHU9GBe44iTHVREILJlgEvagAjOevh8wp0JJ9QiJxz4RYs6+4Q/O
4W4eniUQk3315kL6FBk/WHFD1e75jbWmx+BeyGaVZiCbmFtVksUZh8uh583i93TQ
zkUbm47E2sueS5ym3I5WUzL+s96tmwNPictJJRqopgaIxupEAcc2wruZAA2/scij
Hylp5qfi2nXwX2gFLcPcgL+ReBm4lXLRHhpVz/xG1ioy3yDzYrfL/OQ98ZK0gvPW
0sYYdWtiTStHUh6DvFmbarbEDBwDVMGbixUu9hcD7Vr9maDF9Hmlj/BZ+a6TZBcb
IkpJX3E2uTQizxgcIkmuGJJYFVWhdGmdgqTR23X6uKuztogCyjjOK4+jD3WkqdxS
it+6Kpsl2CBrKKb3qfWbd3P8E0ML/xjQ7don6RVdpBolxZ+lOcktK+kTYM8kZfUi
Gf6iOxoH8xAIgEzk4/0Zf6bZNRyen5NaQZuCWxcRatA4Wl6wojge/VJqrn9eIX6/
7Cw5Z2O+JgLa0LqArVc5ENTw4sfN4LHNXXNZ56gUvNKtiHuOchW3O2dLpkEusQRM
mZbBHrcdj4soeuiIGDyZIF4rxTeAnYVCsA5J/znJJJd5rXPXF9YpTvfp9NrPHZO+
/Ogri6ZsByx3+t2HaW8GQs0FCJFsnCyFaNqcys03EjBQpCZb3bOcIAclEe1HfASs
UBQpElWrM0a70Bq/nbGa9y3GvKo3XX6DbbyXShbWGODCEXtx6ix4CRIsCibBG/T4
arqEaHFpUUt9CqIzqeee0OhFm0M42ft/OcW+RKpBO0jizSuTutXFSuEPTOmJskgO
EwwDBYp6kXqXG7+N40vZOaGvA7eSJXB2D5xOHVmGaOGIgCiLBu+mViAOm5N47TxA
9O70g1v02CCdET2g2nx2uDU6E1UFMgF+k0ChB3Uyq4dfrXh/0cyjyVbjOZeruNpg
kB/FFey2dslArHvO2fDz5dDCMbnp63Xe/oVbK7ftbNHeFGQdmLvdx4pcJFGXTME7
mYKHSf3SZOo/ZiPZ9grZq8KCK9Yu/tCLK9GWlIgcq0bbSg7xxIVuSAB5tB1cLO0n
MYLXna6HR6L1GMaDd6Y6tR5D/G9T09OBwmttj53VK5DqGHaQGZVLB+ZD+ritQper
zLs641c+27U5/fvUgTAhW2dGzLwDW1mW8N6joIkE3TCZ0UmN7oCSdPb7E7va1bFl
1eaZSwQflj9B6D5Q4xfYeV2pn/i9w7qEpu3s43LWCwTPKsOUfF0b2HKYd8zYjVxu
QpfOXewswAg2CTMi8yA14XWOo7vPWHfxRfB+P75f2JvS+mM1qKoRnMeRpFrfs+tR
S9gzDzJdIIYwvDLFPVy4hUvzuDkiSY6FLb5R0Hey1RDTydlJbNnNggsm7+Dtb+dx
0CcMC6CTD0Tyqj99qTeLn+Gq3fgyk40evHMlpYqIvuT2Ra91OPxe1tiDNmDgVOtj
kF3JTu8E9a+vF5nCcZIQwdD4ZAFwEckV7t8kh/Sd/jlo/MCr1Sj95Zlr57Zn9Sul
xb15X990tNNb25ggu/k1iFfKJRfmwp835LQ0yoSppTBspXRx4pP88oET4aMe8l+R
eqPH7ITnmoEYd6uzuv4IOLNDk1lzryEeaZGrdCTywWeOUMzj0sg3JbwhPAwBfebc
tQJxG9EZIM7MMi3F3jK2KMJLZRc5pEPFpa3c0evdgGVOXzjSMjcmE3CAo21KLpH1
Q3aYC8bPw3cSW4zzLfu+ZeocYk+woZVb1Vjpi9Mr2Ukf35Ul2S2chvmCOsyQBPSW
BzA8BdAEchzUOMlt5sKV4r3CSXOnBBSYQ6CP/6LoOolPgDKt8o/EYy29aIfJI4cW
ZiI5ox+zokttunMWiP+aeAmPOjckD+CinrYXg+7jWuP3iSXwtNSQSD0eAICUOad/
eJEM3urdlIrPXmV4n95Gzvrrc/3eyalXBn/BnPLS923kfFUPrmDb+Zxsd40oag/7
u2PmuwnHUBWih+kUokVK/KvaMH8hw/D3Gt2AJYgNNhsXCdZBkSZi3EI7nYzIabYn
HBZ1WXZFYjmoi0b18tZcyg++kcsCTsi6N/DlHOHtZ9YU+cToAA607rtCNF6DlAnM
RQxmBZ+zkW7hYAwYTAatSrl6eAsXlnuAEU4umOKdy6oJfi0fpkYMHskrY8rYFGFf
hLj/xkJp++2LSqfwg31luGMRmlbaMPUKdz4ZtdHWugTtQrleLhGp0xlrFA6ygPW6
F4WNNIz9DzeFJUgHbczCbC0Q2ugQOnfQKhQEi7ULLQvyyoSNyLVMSK31MzvhUwEZ
d9s/HVxmtzCnydScqP7Qove33wZzjPm3is2JwE5MxyHjYq6fI0mNBhSPAzeS3K1t
CytkSeVudUxf3nhk9w3FClmmXCUvyT7OYh1vYolMzV6LpZElv1yup2/OD3gWPERH
vHXwlcrjJp1eFfXPWgpOVyjBXe5RbzStsr1UXU7Pp7M2Cyu0zVj3HHsL0Q6Q/hmn
iH6Sd8NXHB3+BD/B9L1B5c7nuVv7JdBvQg0o1x2eNEgV4ccp1rY+dPFcrSpuK2re
hcv4w8TsDB0yililsGfJMTVfOJ2dsBNvMntUTCyFfskv28Vlhr3q5M4ilKtvEXCx
z6hbaILQd6UvKU0hOLi9v9dTsZdgn/1UucF+t1rojlrWiX4CwJknxNNLpSzQ0csg
Y2QPCKJ3qkloWhFejYlkvarmtpZWIM4D94oKjYV7aom6sd2eAZ689bNK2KtyL3/h
7gswLxsfi+hK6F4ifYAiaVp6n6dZE+LJoBxQqNwEt3NP4PkHDUE+f2oc17d3f+1R
XTAaeSXNiiqnfuZ//BkMJJUotd0Sn8zHr20co/+dsIdxtRfaZZKoJvqwcnXY4uLP
otRufGXSUEnTOxr92rwqgA1GVyVVbfdM4nT6WfaV06odYfqs2IR8pQ/4a8g6Dqsj
QH1YN40UfgbFNRDpUYxLCQMoLNjXjtZeA2kvFZZAXtRDp0cemNY9VyCdTiBSppfL
NSzzF18wFcgbPYJZYRtst3pbzcfrVOKeioznQ4isenWfTDcPqjF5dmc+O8Y+nCYn
Vnm53x2IPexXmxnSKO2U2g==
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:21 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o68Kttsm08/d4lL+e/lzCKEZR0TVlpr3qhoUhaOpf7nQ+m5dn/F6bOzKIg4K8E6g
lwpYIFM00ox5T8IXmzTXEHiqaJb1BVZh43nPz6AQ7qiFEpTObG+ZU6lt+O7152Y2
6dEoEajB03hEhSQ72G+GE3JTeKpovTPE8URVXfw8LTE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 59184)
V5+53TarFn+CKfPDbn5YUuS4HsS9spqAOvoWQg1eY1AdsAJZTteUtPw4zknIC7lx
oEWEWNO1vWWe7lRZMRclXEPP5b/1PGY/n4eZI+eynJf7JT/ELxOm/2Qz62X6iQOE
uou7LWAHShgEMw7izuZoYKy3GPPGvT4DHgqpH3Eo/gCPiF4O1tIiHo942XTQblOv
39NfIcLxvFy2WC4GXVZoa32W9f4GbjtVRAQ05h4J7SEG05xktO7fmndtIDEiSwfC
ocPT5Z3Bn/ejHUVIFugD6R1kRVzxnSbQyjgaPy6dxKe8cUy/8LyPeeWl89hbJ0wU
Rn35xrtxKEB0M4W9SnKlO+/r/4x/goTmjJR5JP6nNfQsNiCXdF9Nc0E8P8PGfI1N
RnUQK7YYGkSBWwluhMrc7xTVvOpX6VEvUiXUTq0j/INSQx+V/BE4SM16HBvXtAga
/ioYu/uOfXXc8zXXRArc3Lz+v617fSiRn5BDDiI2YjpONcNqMmE3Q2IwM/NDR5TG
qZ0my7ZQecOcBvk8kC90hf1p4IGJrBYXv59jA60ROnEFuSnz45ja6JNxM64+SB55
m0MHoT7H1p/X+EDHTY8r5f0a0UOwjTKC2LlEFpG6yXAQwpwwExacjRrk8nl6RlSo
V+f/pRDynlRrWVozkyP+UtRe6oUZEN0MEY5Agart4MBgaVv025omsdN4e12HfvmJ
2OS35SyvRuxBuYqheUu+sbU+9+WwsQgQMyw4LqJQVzjwxu+/OjX3+s/6ysQOQ5Sc
0DC4pYb59qga6lUwciprFrmMhGGGa+8Wiy2wZ7vdReUBcyQNxzR9tDAkZEKBgegv
gkAJw/ZpyVI4azlmhBA6ztYNEVtGMSz38zOOVn+L2SLwRym9C3pMuXPZPh0WWiSa
3ine3S0wx1O+yeLoc2GOHE4USIyveQojaPd+vwKjLa6Zb8AVAdEMYo4V3PEpZ/rr
CFhCmmNxeInvtv9b63UfYzdzZVbuaQgr1yR5Mqsk3ioWxVyupB8qUF67IOuFyilr
KQaKJcfmjlhLlXwIIUQN6I6rCairc6Q3cv3maYEgUI0aKSroDRbfO07n0Q2HYjcC
LwzmjC/1pjFWWEeZ+MBPS23An/gs0bOSwbLxKBTUVSnG7qc+Wg5pCj9q1uWIav6k
5NzUv1afE+2wK9R4M62yWvrtFW7MO9Mz7njzi+jIudcrdBEXjgBkWNaRJsc9fxBl
T7cybCOBeKI1HQbNBPTb7v3TB2m4uzNAMhOy2RUaqPlQ0Ot8R1/NxlxRL6l0bxmU
Wpjp/1Y8DiLrBeX7IhlhqxG7ZXIFCdbcQGBlX9uV3GmjetjCV0nKOjCo26EMl2rX
wkSIL7rvKQVv7MB+OuRrJzM0oE8mO2UOOJIHSJ2RR3Y68xQ3XoSXG6+d3WWItard
BbGfjOLSertKTQDgmVT6IZtu6XNVjGnyUDbDSnSeWC6j7KRg/rbe8fdIoUgrgl1T
wR96BJd0G8Z0im/3Fr6WJjPqXq/IrR3MdK92MqWUW965iFF7d8P7U/9dnlEmCKg9
0+IUsntrJIv6JJyLbEmrOiBT4Nk4D6Xf4gGnsQktFyHoDQXUurgpSpMtxo8437se
V2k3YpIYo75uU+EHaRd13mjfVyuIYMBAXWWgNJAikG9oaC3uQ6iXTgHAdRKMmD+V
RsoMtrk1LUZfswGSeyVFlvFFdhHeWN39Tu/rClHAW3ur0Tl5w2khfDoXlMnbvqMl
0djmbrOKEf7rpVwyeYFlhc/5IKUXlHEV4f+241VNe5m5znTnrX37GoE3GSlxpbnp
8vTdMCBanLiBfLm0RhyDHwjU4cZYUvSn1oyTt2AdVdn0GvDslUh6Q10zolfCYgra
Qoo9xEJJZLeL9LZb6zrGgoTZFZTMqvjcNNmnYsIsB5N5dGvRmMGYIkinOWE/MMfj
lS9U8pVOqF0JsypRk8PGuOslI8+2X5XqRzL4DQe1mNE22mlPtjcpbXJBlcev+Ui/
khUe+9X1yGVaTkyVJA9UUlBw+l7B8+/q1iUIsH+zmOpDSlbnUVlBzROAWyAhwEgO
/NKgIXR5tgs9gAjtaeXXkQL7O56A/oYLdwZPnKyMEUIj0KlCgcQuEtbZ/HaL+wlH
PfiAwQ66OzOh4iOLXzM9B1f3hHVjJCTCmOmv0EqCf24TsNexfUltVrOoc3UDcrFt
LGfL/I/EfdDiPauKy0mgjLMTyVJxBVUxwNclqX7O4OCuzWb3bpfJYFdLN0JzUDFN
3zo0UWKXDWUINRT3TOJGFxFKLDz7aEoVdcaM1OXqeZIhEK3URRabYiF7H8HCQ49o
RYlciFgHoHwA7r6li07v76l+TpP8xsnn7iac2SWD/pumFmK9i7xVdtlJMCZ39Qfa
C9jAiOuQUnCtW6JHc2oFjdPOG168/Rcgq/7p2cyvc9Qogmc2rEnyBpiOghbvgl31
TPROCkX9D+IlMI0jKB/FMuyQF3W17W+rX4S7blNtHQfSkR4W+Xd4KTdAwWsxnBFO
CffpE4zSY/O7XKExKSSNFSzB3sVGTwfhbWPPd0JRB4XJdmYWolgIsZizPlBW6vyZ
k1YlmK9Hhxs8rXffWY7a5euhrIWof9eoS51+9f4C3mIR6mHHTAZwIvb42GEafbwf
PzB4fq+yz0eK1kqyiLEZUGk3BGHTrpVDTKtWdvg7Io30d5vLoWekxgwRnZPDZVyP
1jTWLPPRC3oH23f0SQUQ5fJtfkbaZpphhh25JGQWaxQB4CaAL7LW9jFwAAJiwhTA
pMldTE+wiVybbzxxWQyXAPgzLE6ntpNO8m1yhWeyFG6nBayHghaURv6oXysew0sQ
hEdlkh3wh4X6SjpSDpuyjsp/TxhOR5LqztlAy1wahlzDvJoY6Nw/9dLF+KJF7J8J
MKumo4nB86IUwuypk4054PWqe46vzoOkvJJLou3zhVH2oGz9xNSWuljcrGzLCK5J
FE1PgsG6HbEbCuA8StFBUpuVGyPYnsWJyxEbFbXfXtlzn/jSJqcI0JIFWjjt4rrS
Ntfc+ND67iQQ6abfTVOAuJfKgKVV7dpdT+FgPZ8i5NraPYtsp8UWAMnb1RqvVDp7
9OqjzDJ5moG+3CSLKjerjlvMXVW618WYOW7JfGyqpSoaeLjcPXFGi6sg6lzq9Bpk
3iia13Bes//Jwmk2GN4yB5uIkAFOj6FUhVYahD6/e5aCZRjlO96DAEhGdtuETqqi
rjiArRcxzTFDQTHLU/7YsswOZ6L5VmLQPHMGysVF5uy/K4tgmlRMlXmEzrlvyLA3
hg22JX2Cq40YPugkU2XrCYVA8zyhXgNF0NxUZ0SF/ZmtqC//O1owd3eJMmgOUFdc
auiLADMPAPjKoEFPrEslb9SnIVwkVO//mWeHj9rMSgunk94rFReB+DGR24no07iJ
tx+LvL/TMexPgUUSf7umqPofJ6cTRy0KwOUVnGS4GkrstSwO/XNcjT0E5Nj1rTac
rQnQOh7fMko56m724AsewGtbQJxH19U1Bs4fvF4qdmxEXPozyWeqEMHXkSQtKLLi
Jul5q3DEZ3IplosrPXTwpfJyauprGsf3rTntJU+hXvO9UI3WjPKzpvwTAHve3Nnr
Bk/NJMSPBNIZo6qiYWIMw93bxxY0raWSeuMeP+JN3/bOjE6XXXTWgbXS6RyhgI2E
WrmligCMyVs73YBJ+8oZeCEQ5Fas0tiDpiqA5a59vsCPWE0FobnzvuI29hINoEao
aTb4YbWhu0I346TV+IvihXEoefA9S4MSTshpQ02zh6vODQb/oX0/myYsWJSZ0Aau
WTLIxiB9U+DIlxvev3LO/Jn1BSDcHLmDnpxbkF0lzk8euBN+QG0FHDpkNFW9YwgN
7TbawGk9u3bl4aiYL3uLBCubvNjdJc/tfFjXjEW8ylVv9A05ocjjF+Jjepw7NcVT
Mm4lbowTanCsKAlibKrXSGaVTZs67SeXqoIxCOMHF5OepBxmRGttCb34xj2jf4/F
GvKl331zvWRDE/e37pHlQvWNEagRmdNcKcIASE+Dm6hCRdWE3wtBggepquX/Bdn0
9LHTA2J1mS+XATQmxYp/LALUOwJNG+6tQp8gYBvc6egBhXKgboxphl1XsTofk9Nw
GqHH7jgUCvvnHkZS4mQA5TxeukSMSjeCZsOR0RKv6HBDu/XHRmlkYLTM72gdTBTj
uTysQVzv6AE4XdUO7C7bl5PeFD0QBh1pqUWjbpXpwQ5rthXronGTi+m5pKFyJWlO
Lf2cl19OVw0QbntTIchkXy6yeD3SwopyAOjZeVvZjXtoFnoPhJm5fVPRJOBvqxe5
LK3aFRKMVaOej0hfspzI9tmU5NaSwAQt5QVeQmAfERc2vxZh4CiLj7P0W99wzZDC
GdAG9svQxx1pFP8X7q6QrRRh101fy1BXhRtLGD97drqyaOpi+1991c5vx5pALt0r
+IC5CVqx6hlq/SsKkymIhArGt8gDb9UjFehuD32zdlLhF+/EREM58bwFhpHIS4YH
pJwDuljz0GWEk1Q3hKZUXBow4XBkV/pWDim2u3LwBDnh/ievn+lAy1IqR0Q6INNQ
YSP5Gtm6trjyLxjE/P+r1TIs6ABwrwPcAppYlHH0pXNGLlkYuhbpYet3d7njWgsa
cs+XkAmqr6qwBcZq9/fOq1TPpf+92mNnEXwHlZY/kNWutNzdlSYuQ9AdPrkVZcEa
OHf00/ulz8+eAR4SWrZfVWO9ToC/+mvJWXKtH4MYYXwZG/mw9O1pgVI94D/aez3W
PHCOHFvzGn+Ja4DZ3KaOR852nTL6BdeVivbOXEL0GpT6ebQo62Ej1x++q3fruTeE
U95eVozO3S1AUHK03zPgZILbARRGBZRqB/dgmEaA8cPH59H/S1NHgyWGY9jUEnN5
OwPsIKqdIzt+aXHwo80sdYfdxO/JzbNVSyfoFIyupZpcjBtbvSkc4eJpO2rzp5La
pOtKZOuRM7sR706Fj2qfnZ2n/OfRJ3ya76aBX+pSiMnwTyFach/MkU8et/eD6mKN
L75atrjAiv2xe8YqR8+X9ZHZc2yCZvv4DgrXEK61tlTxGq5UPvbFrRTtdzjw8kDQ
Va7nM4eR6+GMrt8b+lR+SjWGhFR0Tu1qJlzRJKz90O532rwlhgz5Qdb3OcLIvZPH
VZV64U+gCUM3y/b6n8JUFlFp5umtfh7qUeeGKJAgMpc814Mk38t1Bie6MSB65fTA
OEfTUv50WdZvZr6BrpfaT/JCH9apVeCXBTVG9IDWzmIbuqXPFO5wNL3gPUQR2AXt
fpuaZNDtccWbRzOsv3vY37xHI+MLXFP4Tj4YEL97gp0nz7870vgDkYILECVG88EQ
oSjm4ATIns99kjJVuazUDZ+cG/NQCDoyuDvqRyejZoIDNbHGMbaQ2bmou0WVE56/
u3hdUU8q9MRpBLtERLPR/W7b9Zxbzr/wLirXkfsOZypJe6r7nfoH4LIwjzg4cU4X
MsLJBcBxBvBvpxt4aYoVoTuzAu1t7P5ONZFg6e+PkQw7UcNRppOe9rG+1oy4+Hsn
DlkHLb493VRNXnckkorWzPkGtDZSYHpaokDTJN76OfsaJBdVigj1jq4OC1VZR0w9
HBq1Z/KbDNE5l0g4qX5beLyYc7M9pK9Yj//TkPZ11jL4eqB74VLD4VXLMt17qbkk
zC+bii3yV0HtNgvGEx39carYe6KXnR0k4wXZnkmhwJ8BBJgPUUw71lzv2umvNdo0
dUTIQqs9xWlMAo/ETh7WmchNs7MxY76/f8dZP6jVXC1S0YpyWgBVtnjnEewfXZGq
4BCogwcYty4UJh8OU8JOiXsZKUCExqor1/rv2QfmK7gexhNj7lrMDQxALGnw9cEG
5MGTCQsearthNApPTAZ9qSFP4+zMAxNXJs2Ir3OYc1TYB365jOIfxXjwNdSPSYns
Ebkk8vJi12ermx9Tn+sJ8OX+ZNXpClKFufpPa5PX4pbUNAmBjL6LWRJDTZAt8a2o
dCmQSdbkU5KB1+9LXv4DZsIrvLyV5IYqyDIYfeLug8t8Hs7YvRWdzB7ExzAJ1+V+
nu03c67yy/l/ONpBzI1nGUBCrBIoD35W2c053EnsoFLrzpBfIfjVX/hR/rJm9CXQ
OWucsioy4E0Z9bx+qv7yGHZ+z8HHbGf+t1LD3GEjHwFbXh3hqK2J6JALSYiKcLLa
tDsxP90cs5HWGrLIXiMQ/M029dYsRahRht+WwdFlHICX3dJopBswTsNd0ZltXWk6
FdEE+a0r8nWkqAJ5PI0Otijp96ISdPIExHGCTejOAepMJ+bC8msEPIdrIXH0P3pv
OwXSaY5zJBLh7jEBNdkA+WlAX0xW0W6rPPH9d+tbAZlPjzIVfMIuh4ljSWI9RyMi
CxBEl4gVnEsSThGQBCP5sjIipBnLorPwVt5mETu76/liIS54mrZevO8jSJEivdxF
qZLcOZtBXZxPg7As8ctOrmAgi5NP03ImLg5GmN7NZ/UiVp/8fDqJKqVl/hdRnOJw
GQYRCi9wGp+heQm8QfzvYEKMxFvTUranWQS6HkUwa66WW6zLGuf9ukb92nKUkmHJ
tGqheLcEmaKEFUDyp2DePUG7lQ5Czow6NtluvkAK2cP+jLROO4IqUoDPHGNaw8mh
ImHgyscEtFVXsV5czV3UT3wJhgtgoL5D7EbxGypZ+b/5hYsptGt9bVrJ1kA8mply
JZR2nzKu5AIYIpZdnpMxbWCC5gBnxMniHKL7c4dMjYg7YlgPufGpHjT8IzQ6x/cR
YwgmzT5nOVNY/+n+L2LERYnlAC3WIiYv21CPpHGZ4k0WlGjOfhEAivTX2EPc0vLH
TmHbQ9I+rMJ8otXBN1HgPSyIVooQFRQj06ba1fTTmc2nWsVw72u0nWaP6gHpDHZ6
FKEi8DJmsVUwyZzqOxFWeCjKNzx2aI0YKnc5IKOenyKuml0s3FhZxrEO7xNBamce
vpacc+28GhbaurBZI9y4+jUjAHBosXsb7S194oryxuGEAN++/qeLccJj9i5HAMm4
ZhEN80oh9lZ8jkDSl5VGqdaAGt8+tSFAVi8mRYxt3zuFDTXdNSOI8q2jxQYoi+5k
p9TmUbw4qe6ZNvHVWjN/ALAKGhSpRALZuCgzJ6EB5vv8mxQHUXnLMifW64ficYpK
NpJdaGnXuv5Dq4WHMIlNVqvf2r3AVs/sk1wGtfF3tb6AGgzkl1rpg9t6FlwCGsAe
xKqkXdN0CorMs1nM0zxwjzYVc/0/0ACKY1FPIJaK9rYjqv5NZiNRPqYsxt/N581O
mfGEfeaGAFtkBKCoWkr+C9CSO006/ovle5b/KssYCR0I8TPZ4NfMXBFAjyS3mDaQ
5vbtkvDkIOAetV7uQ3FAX6Ja2GOLTXA2ni/u5p2kqKQEXvKQ1xq8rzQP+sKQg0yn
ucskBzIFbdD4mkxn+kFx0a6gntnRhmHraTrKcKeEhzhOVSWXEC5wlWxpAo9dSIeo
Th6lX0wQyAocZfQ//MiQIBRiI7u8dr9vDx6BYT3Adh387ncLP8S1d2fATrC0ycvw
cnZCAqeTfwgasJ65nGLiu4UbL+2Ug3QsRSsdB3roD6j8Dzsdcr2SFKbXCZ3++YzW
uUgWlf6PexMj4mraaI5CdFeVNZ+8EvnQC6VhELC0JpyweL01LZnePNubGDoYhXx5
mdM168MPe/7Ty/ZFewFkdEqC9RcP1YEF4UZNYxFlwZMoN3QsmJ/UnlrpNznw1omk
ref+ULqhdIQgRY8VO6JX8SDN6GGN59EVuPLyCb+y5/upORAsZZHfp09Dm27Zqn69
N4n17zbAiQhsMPiV7JCDkOTr9ChxDBNBRDCIT+3oMntHP2hUcn0Ek7p+LVjawvoK
ozUskzbOF1FLMNTShvVkkWOYiW/MSJf7kUF26C5du7oNFErSpLh+MRWsYi4GgGuC
IbMYdL38orl/gzInxMILYrVee992c2qQlZ2kO98sY82OUrp2pG/jlvT0lGFtO5Id
Nb4xTjjubiUlXBqIdygknnE8zp5oJ6nrcs3vMy2OwiXSFHjHcLBCvKMjQRyOAoxV
3miVUuMKPgRcyuZ/5iZh3eY/1NlJlxFODu0yqZuQu7qwapL9PmOZlXPuRdfMjRT4
/TZXX6skYWDOg9uHdyQo3eHK1RvS7JuQ7QKhIxZZhYpmov2db0VliGWBU4FjJUg+
9CgLr5xZ2O21EMt3WvN72/P1vawaYRj4qYXJ/X+t068bES7bYii5/aEpaGAPNWgx
4UHksNMUO+0yNhr3/twbfJ1B7vCftBLVS7ypyD5+7+cQuGh5cSy0PEX9EqYiL9h4
f1iYcMcYgnVmcZj3P1R46nGI6/MIxJUWQZS64s0ZMGe7wEFF0qyWGmlxjIMsKvx5
HyL48ZB2TdyG7/3scR3pmu6MEuBHcgkWVCmWGDYEMZNUn79Sl0xfGWd+S4dXnWUm
FgoQQy4Iwl4by1xk1MhMa88iaxLeSW5QS6ffdt/V6K2lCB1vpRWIgOG4ciRJpija
JJxUPnkM/pfl1KL2JgGMxFMtfx/wRrKmUUEgXfJcuG0SSRz3mlCWsnLr6t6PrbeY
teYYHpP8mh4IdMkTHXFOWle8LBVRcfz85v39lEeVGyMtUfNhtt56bm2Dtwf40J/L
c+ql/hBD6TlRSy1/oSJ5JnNC+1gPQ+Aro3QqJ+GocyuYGFZk9YHUBsYrapLtJwjN
6cMBSHNXf52QN0bsvi74vC/7ENdzwRyL359LoVxBrvyWp4TUi0gzV0kJD9XKyglF
Fhe+6gCmI5gwiW/3A5gSMJMFX8HhQHk5bHxFi2AWHX82uuJuxetKvFFsWNyHGVZK
P6+Qgf6KnEdFfqfLM6exKAJdmIhGfnwWOcrRiy00cTe2HbSenov9Qz5qafUMjLsF
3+BA3D5U+AKjHQpYFSmeotXijVtOZabWAdNrdez3J4duDbn0Pddzi+X0OQ87AaWJ
t3EQkNgJ0a5Lu4k7lUNJTIFSXkSGE02pesd/hTAsAfWQz2/EFNgkUuK/jKyXuZe4
fvPiFQatDCQUVdVK0aNfsyW945lKvhltvUb/SD89c7uqvOWg8GKQ8xKnFIWagPDM
ZlmrtLTD6cO6IrbDcDPxKDYdoRCjBi7l2GDU0NJAAlqH8mRYYlNfgj8kkW6B1Je+
fiOtYBol4lXlf7bAClxksZ2L151m5lVeIZsmJK4Bp0rk6b/oSk88/WetePbFNwDV
9IyNJRjJsxMXQZV1OBwVA1lvfzDHjAWu/V0OUTV1K3rVBR/HeV3p6A+G1c5Pdqmk
SFPiBFZKKHToCCaekgtiGK0QwH8arLyp2SSNLQ+D04qkbfPxsJl8aOuiyUwROs8c
jU8d3VKu+RRlvCsNQUlHR/bFL0AzmcDRFbDpx8OLbM6vMqT97aDjBm9MhkD1YmFm
qOZ0KOzsx9XNyzql7GiTFs/eD2oRzTgoQRkD5kqKae7jdGliYgUKZU2i8ZALCXre
upG/HLn6A0U7N4qU8RiF0H4LrQWODvsHsaBIks/akpR+VGkm50aYpcBVAiUYeYav
3QWc9ugmYwbhFZ5vb6bEJKJHJ77GGShstRhwONwPptZH3umvKBtB0tATRAfyLMXo
WH/Zss2aeZ9HGDX8V4KzA9rGhvbMi1bYfIOWD7ZA7gOu8tDSx0PU6o1B+2oKf/AZ
XpNlobLsN32rNFTjayo1BtfOtB4ukSh0hXSLT/49m7fTdjl9affSN2TpTCvu+28w
I6gZIQXirZv9Oh+Cw6POA+A242HZjD3+83+heQ4c17FTApyagWzbSiDBunuNyOGa
vLmYKCPLlhS1keIOfZ+0M2pw3DfqBCllJJhacZDm9WpnwW6IltxDoDg5r1NPCUwl
ACZKsZNpFOwZMkwW7PuJTBNLf/Jzxh+WRBd8rivBJK8INzHx+cQ+kfh5btMhZMQh
1Xy3j0dlAnqCbp7chAprZiKzmgpobYAdZQmo+IXqhWHdzEb43NTzc37dkYv/6Rwd
fx8yDZwOQg32BCztm9geK7CnI6nBDYVg2jIwJ+OUQkA4W4MqZoAML1VbaRh9Q6lr
YogSlPUDC+XMZqo/xJvvg5AkBm16/BeeonRTWnIRn4wxLGeDyaBnYTCP2Ik/h+qu
wZz0+UrQQa6nMmX/F9M6pSRw+Rb0LntDQsruD92+5Br7C2luOLOoXtL41EVThlP2
dAMSDWdRaVghyz88KV4WuU087eQY/wxGWKqQihanYy2QjA+O0g9lngv6wjE3wOLx
wpyloffvgPZkSlMcD4UtQtkYvqxqNfTi+6tCXxWy571XAAIIuF3DSGBng97EhHts
rHluy9Qu6Y4EcHffr56lnMCp5yK7AxEv2F264/OnLjNryKf1raA3P/Mby4zTINYY
aGb2YLNxZAyRjc+1u4uondgJq1mfQ0aeNMBrqph4IixegEfvlnoZqGXOXysJS+vq
adyUak6+4OiA6dVQPS0Zj2UPpAEaAGdc85SheRKTv+OsOnFK4Y8cQA+nJJOSLCQg
1aNd0pWUvgha2DVf/qH6zK37McPGOaURtONplSLml9+grPM7DmTP4xBxf5IgddJt
8GExDIGiNsqwrPJwjhiX33s2kIOfZoWPIWQeBm2rGVnVGZ0ND/8gJEpaiJkQU9E3
h3r8d/r25RHjsGo81aVUF/TWFYlVzemzTn/gxazI3wkQBRrdSa+evyLfffiKSUT8
vuc23oUuWrKhPyDAJej2gskOMuUTNbPIc/iE+9I/geNXLM60ZhseQIZMyItW/lLY
8PzV36KnoTpoEmhiAa1OiV82SrVPkXAcJyTNUr/+2v9nnPXJqVGjUxw5vbpHjyR/
rZ3GweeyXHahv5xnKAHzJSiMmCBOiDtNPGOGyejvlr8MaoiI75E7YyUKbwB18JhV
esBtaBuE0E0nNsLhBbWPlYnLDK9DsEEP45/C+eaf1qHwiqO1R7249pWWVQzREmX0
8DK7XwYeOmUpR/y9WNsX3pAm1/aTavkD8pznyLHKelijCvhNlEvHWsbRvaHQ1Fkv
G4poQDhPPbiov8pM44Z31w22dnNL1Tx+e2QPfSp+FYiPDYXSln8LcTxkD2pVCuKm
mLtLiIaNuDIi5xRou4IaickH1SgU8F58aflimGRdIYCP2dOGwxtXPvZgLPSvQHDx
5Nk8Ujo6ljuJe0CuputNOJ7uDeqfYjlY9mEwB/phJRnhKOr24t7G3yWpYuRByH9v
z8+16gB9rXXt9/9HcGHv2ynCRo/Xsfc8k1WFPjNMVwcK7MHLH3MiMcGEFXg6K6Dp
oz0wS0bZt2Wb90Aq7xwGOiQtrRSioTkauWJvr2ItnC77uwq3nEyiBnwCC2JdcJO5
EGVV4x/sOpVEF9N4nIr8Tj1iKiu86tcXyoeCFCcPUgj5hC3+6t01Nl32EZ50R/hh
pwEmH4MXtpclMLiQNxOv0iE3ququig0eea/15QZx2OsiWbiEHVgEqpz+gJXdi93V
VVr5P+Xvf3eTRbz1+1NzQDnSX5PU4rhN/vzSe44/Boih1i9P9nisfuiGGaGNCx4N
RKlKCnLJWy7nVjr2b3plY+by2yWy7EYUEFx1KhBsL7xRQEOA9SmVKmZ/3jihjCQz
YFZzyvqrTSy2uTBKBOAxwJXKSDLXbN+Ga+G4jGgpPM340B9T7kaoP6xa7CTo1qSh
tr9Ynrebubnq1zD1uvlHoIKtbQI2QVLpcIWjHjk6YwYwmWYCuM9fQ6H/u0OjQFuP
zMnNTHlmb4Km7NgR6z/JeUKxOp3P2V95wN/Co409FdyXvwHxnKYAOSzua9WoAzO2
o8zVvkIoOfb6RIGKjANdrW4AFuiuD6H7OPxocJrKF61Vb06WVTKjFhygOgBbXTcO
DExGcmwGLqlj6jmsWYPeTF4Mc86PCCwhaGIXR+j229CB7q1MdEVGXKLwMq2m1h2s
sLqyMbhmdv0ry6E+PPK0wZziy+1Ezi4fqzTAlYOBbfkyJ++myRUjN0yZTTgOQp6a
KQ+hHWahOOChPQkUR5CKCnRq6hys+mKBzXrBQiIdmxm2uV4ogBUlOYBR14SxP1fP
dKN6bpaoYfcYNfHtad1Id90xlhrA+IDhFBhRgihAvL7eQekLZ+hZtS2j8CNPWDo1
h9EWafzETQnwQ4XdXi9GOvmcHTEO3gf2mLERFRC4KwwbxuGth8bNwmfWgTo639nc
wDBtPXvz/oJBVc9J7yONZYxGrllcHPKd9xDXot7C54Iq2Xwkimr8nnM/E2E9sEP1
78JoSoC75sNQ22ZYtyGJ46S4RLrts/5tMGN1ohnAIyL+7+VqXYibmQVFci27Rv4O
RMS2ub3O9SIWhq5rbIPYB26AMCP5f1pojOZ0Pwc1g65mafi06iL2c0Mgoepdzjku
swTOL+v2U7OEAB3CrQ/uljiBPVcHY+vjMOjtthdvPlhNf798AGOJQMZht2aSsNjX
/MwtUP7UqwG8jNIDeqm4H1dLRKUFURJdAjtLExHSTgDTUcCQ3EHc6KtPxQNEkitJ
p0u8g0BNTRXtgN1SEiK0HKtYxCeR/YTlXn4GVo6n59DlLDwNY1eNAc8v9WiUPuXM
QDyAq++c2lWeRVwtU3zgeQwTpo6j7O43F4cfixHs5o05wQyEQr2JHLrSTeKxPSy1
xr6zM8w96dmWriJxvAFi7rKCAVvrDHfssTf/b5lm/mvDI58Jtc64HpZTei4TDi03
V4nkzUfY5LKz/+DpjhSLGcCUcsHpkQzUzTij6nGOhGd2tAvW6IDTln2v71/hZb8w
FnQfn40KdjUZ1Se/EUdtaI0WKg3DrKJWimNA2XlJv+W3MvmhrIx/rzK6VKHR3rEw
R1h4m3NMeULF24kgOmcyuQ2oT4Kj9KGgFuuJVQbhxJoQr/s2Q+QFPT80fJDJ3y8X
IJGEArWeW+4H+uJwuCpDIIw7VLIhRlvghpg7fl8zhaeW8GyDcy4tFamjztIvlsNm
FyR/zaB7bvrfdB55+rt1FR11+o5h8at/4ylrtiYw/lB1899qhSPQrJqSVf5v09c2
tNB0GWOIxKXN3S2HM+P6J7i7+vYOUynQZqdv+RM6sx2dxKMmyH1x2VG6d1qBkFq9
Gdov6dYbGJ8TJ/0Pg5dGcIAVplTlJXWegLaR1z8DYhG+n0RX65HspI2+BgDfJd6h
78fEKcEvBIjjhndxzY1epbDbxcDCPgRkIJtnVzt444r6w/jQVifrM5loI93tNyA0
z+9rFbrWU4Ml4t6PLLdFTZumTJUxqYVh+BFBYie6A0SVwrZLiHocITAKgACLbM84
Wai505OWU4rdDf1NZzZaW/TSWPOegIIE/vAAVWt7Rt5XeRu2rH4e140WCyG3b/pO
DVMuO2sZEioRKFJFMRxIWDHTR+XwE7PJ8UiQnxLUUZUpk7KKu0ybCgfIK78UkvFH
n2oyzGqtfAXUN1APIJ3VuL7ZgYZUnCq78qV9Jzt2XC+28fMkqS+Tzlaar0Mp86aj
nw4bGrkQ9FDtZHA2xPvCfKdH9oH8jW1Vcvd9WyiU5Cp7MQTNHEk3w5owYJcMsDuM
r0b4oz2AXpFJTnJ+gvUeVTRbPVbr5wjMqpdEgt+JFk8xXoOQG7fEsF5BEvOD8ut7
lJh+5J10Gv8H1bCDt2sZBzP7zqbetBGbuviMJ245ZLy0v4H45vmi9zd9ycxURz1h
WQQMNCVEB07NaQWE/frFrL8Z2cNygbLJq3UeXI6FkNSaqhgy7Os5IvM3wlPNFXkl
j5lqDz3B7PipOxty+HtlM3iOxvlOK1mFDO+45Buo9qH1Je8FpTfIO1mAOpomXPmg
hTcWrjLmiDdYk5YhwlA6klOrMOcxIO+alXBM6AbbM6r5IIYMblrP1M3MD3O0DlAL
dQETXQxJTMug2fvVCkC34BXgW35QSAcDkziCocoUQcy2JPqIZgE012Hm08l181BH
Rz5scOiwzZSGPUI2m879VEKOfSXEixizfrGowIHAnEJBctgs6UCZ/E4v5zHuwN2N
NHdULZSK/IA5eNgxorfcW+8VRsY4K92XYwpGLnPY58xXQu/mN/3PaWBhfHyQE13x
GCT8EippCHUBGrXlcsHw71sRLWhnwjElMhBB27a8N7sP/IoO1vMTgeglbzateI98
pGIUVPnck3u0wIO7R8jDZT7bA7Y6UIWp+2Vjgd8kQeyvVuJyFKKTz3CkUYAsQTOx
zGVYWS8Ehx9AmJOcO7DC1XvoznGinIpIObH5Zx5YAf90nGMdVDAnFgfUvF1tA7Xd
6lQ3Qqjc1wq0GhcKVwE3wjlYB0Mb1keOEqWH7lQmNEic1ChujtHvwxdwN9/n59DZ
h2yA/cGp1h3jbP8LTz5qPmnAu9WU30iqfJsubcgD/+3pPLT4OZv8pa2iMps1PYoK
wSlp6/QOAvyhD6T0dOauTS96dYfLW2m/DzeiWfyVREeVK+KU01kKQbsPFlPFi0nl
D/AXXQ6g2BCKDTDqMbWSXTVSV0nSSm2WOpiqyo1Kh29kFMbDu/GgIYS/LSaZQ3OA
jQT3aZWQ2tpZFKjl8JbPCN14QPtSUEtTcY5U8u+vWA+6p+2JY/eVmFTErVMAgMtq
y3MWFj7ZGB/FBUs4h/75uJ/ohibBXgrsrLaotp2Nopl6UjMZER86MH1mV/BKswAp
oGiAzyO9zCKjHFCVtrJjvsmI+6tIJUafIVf8mIUKA6e2+6yd7C2d508PSK/oSyTv
r009KsGU8VSiVJaapG8l/hQU2VR5rglGvyRj6N0buffToRWuw3lL+HKpNTCxVF5z
VZA6q51JLZjDir1pCv+9tAPtwBPNK4uaQwB6K9EJQZVBAggrWCasVWuJnyExC4E4
wwV9cGYMiEFgcDu9N/16NuE0MkGX2ah4Acd3q6jf/hd2JFU3gzJvtMkFgCHE7gTw
vS2r8SeNfHUECydAswt18lrHVrmdWgR2g6VaUNZM7j/VCH73F57UdF1riEx9zJ2n
9TOr7iPvPArnvFWwGjsYAezntf9Z0crbTfWLjZXfbei4P6U0Is42Wx2h7uhTQjNb
w7T+zYklrdvwKjNPMYYOTuLBDOG+vjZM+q8HW3ZF82W/pT/OZBOcd7UkcVn0hGdb
3+E0zzj/PmP1hJvfbAyHHSSxAoQ4vhaxAQrUPZMXxwJNyk7YU/atYm/fsBKSy+XZ
wKVhDu7Z/9hm6Kk8OW1I1BnqqJWAG4z4OZmERMJieFJqL4nsD95kekhSzltqxR+e
r7IjqAEVDzhgCBHz7i1vNjhvI0fJAJ9/syPIYqS8Pj9CnM67KRY6TT1C/PMgpzX3
vqnx9H3VcPMPjtvaibY9/6NVkmMuWe4y0b5nwKmT0pAp3pgedKAbC7YE99uR2mHO
y+mHusc4vJhK0+lCpDY3zEUwdRX3acBtGE6QNOLxIWXRSOA7l5+jJHnv6esQAjc+
C5v7pz9ARomBVmyU7V/XtTYHDfrQaKdM6s0+VBEMCzb3eSUsk8zEZlTI1F+fDAFB
dTJ2+Y8OYT1xz5aGuB7oDD8WZaNbLZb7uJDrG85Wx5Tti3/FmlJwnYqYWKwqowqE
RqLm9Jzuuca5MvDupUtUGO2pG93lkTkUdvykaAMS3LYVCZ5NCnm6p9FS0DZa/HFa
lUg9wJNeZI7+Zs7XzeezXA2Jw6vQyBS8HWx78Cb6ZGD+0b4GWGogApbsXn+pGt2S
ah1kYO2sBp6QHpiWgofiL951KHnIsKJ6rAy93r/glSBhLCzI8swYEBrYPncaSBKT
jFZygfS6FuZYHhgtc4nduLxXvtqUtDQBIULOppMbYDifahj7/A+lq8A2oMxziCDw
6S0JXqiHgdK/80YBDeNxWzw2zxNCe3k0doemzEGgAzw7KqIPfRTVD0tpzrzkmGSB
nkBtgEP8LL0SQES+o3VExN580b6Tj4Azx+FpZ1YV5xqAidoyDSDnifNaHaxpZwuF
S/g/xMUIW0L5v+6H8SKskyuT8QacuwMeDMHJ/Am1bVPtb3S86aRtwaJ3jNZCG70y
vPOeoOFFHtpywzVEwDlqSnetm+VYbE1QF2Y0PxzEdFs2ITK7VvfpPY2lwxZeenR2
4uq2A0uZ9dCfPrez4Q35k60gNfTZiTmF3yH7c+GeMxq4zZbQECQV36L8v4swntn4
KkPRo0E/6kA08hndYtDCdxjrODPlq6m7X3vJg3MXBAR8tPx+RIG2yUHCMhgiFNtW
N1YyS1XTYK5oCme47kWLc7EvFTSEEMUxfu4ZRAnETebQISvqwG0vBlLLBFambVdo
lKzJk+vYmwW1LjHnbS9arJEWQE+xARQqGrbSeN+bGGXHeRentqQJfJelMJv5Fmxb
YGYnlkosOqiFqeEMtQnpoi7ivucG+5h7yu7ydsQGQyaTkkQXaRDE6QESVn6umU+i
tl5FZqVdbLOYslx/bkbUm0KOK1XnphcKgRIWLWD3KgDRb5dEOoFbzCqprg2owUiw
Q0YR5C2s2+Q6XgxE5rtoHnIgEKolaSjp4BFpiLijN93E+AcXtj3PPI5KjwiSSZgE
9D1DKrbXVX5RhFdYYbAmkByZ34jEYKFbOmC1hNzxhC38gN1rW/Cltz9mCnpwshlG
6g6XrWWoUyTaMHXfCKzJvIXLM90L19VSRCgRqznV+JUfLEVOL1CqJu3f9kToCm38
KrsLgruwEFtyhhh7Oxds/h+macAixvL5QTBx5jOQilJx8PgTj+RqCI2qxsBBzuaY
OZaQ9f7D5GLQQwcSdBB0PUHAvTmpuSGMufLL5ytidZpBwIZvztVNPrXPQseseRwa
uBBndA6BFum/zBkvLkDdkjHJyvW5+3d0dubhm2s89yzy6A3yHRm72q+s07IFYRWC
2KmKT2rcwXQcYB3jvofTA2w1qEhCt8gq/HeUbamZYi/EC2VlGPLs9sOAGMMr+P+r
TwV/An4worLcoVbWm2sGfGXOMhQzuBaq1tl4ejAjCwaNJjBzPs9/xbF/Rc8l0Dyn
AdNqLTsZ22U3o1xDHDxIM8SEUPMZd5qlKVUI+/6mgT/a+/ykQVMXGb1hnCwSZjIB
PwN65hSm8qaJYpHfvJddA5tZoyavZd7AktnXN00lv/hfyVgSR1SXdNyaG1cUjfz+
WqAEHARij5geM7UJTyJRJKykRJ21RhkqXy3mO2BTua8wYeFR0hJnfX6UJua27xi/
laOxqBXybuP5PbWDoUxcICddNl4OwTUNbe4cGfE6oVEgaex5qz+t2TmabaeKv5qq
zFOiPtE1UhtwqwFrFktt7DAXxeegRTwRIHiftblYAeL4q7c6Ua2BxoWk3dEGBtQR
rPh73cxw9puqNsFWkvC5NWsAdQ1mX6J4bO8gkTMoiHXXVGkO8iTZas8nkPV5aJPJ
pbDS1eYSD/Is7plrj97HaWxLNJvoadt0wj6PN72zc1zP07Z42FThVrCELUOUENc4
9aMYPLrKRiVdO9KEjz8Ty8T0rYaOhioo3Po3eRjjG8S+3AeXJu5O6PKvKVwtis1G
7QLwIyVAEDZRFrxCpm34BuOGDbg8oXY/q4kXfyeK/JOGNYpzg07FuLgznAqKSKei
ghToMH+9GWypKvWCQqipcZJrDLeu+M6ca5HY5/a0cC85vwKG5sixYCbBb5UXO9pn
pRqdeOhwJPrz2uxTmy6JQzptND2cqoZCoDHTkSmxt9rWi2KE3SN0AMw7aLq8egon
S/VkvqV2M8Jf1VBx/BWOYWtdXzV2Xl2bRBLgf91uyGAqYRbHeAPPCCFqZ+ni2pUm
nOa1Dt6TIFnPIYDHigvG6oTFcbsvd5MVxIdNea+oXZdG8B0SIHTVeVQt6X0iZRLd
SZETLQ8G+5tXKmGY6og65Jj2/3ZlrO71tjFVUsm6x3pyLWLA1Fs1kJuXGcOk+VgQ
lVbwjm0TIe5h5yLy28PFuLs+jH8CKn45CQbXb+RSWvyTqCD/wgTfvQIml3kNZfiA
X2EI967qJ8geCxi3nqxPpFENszm+mBsIkR1h+lUHS3ueMOz378kWLs8OmQC9Vy69
rmufYEZLIOOlTU0RMShbR0WLJAQONTd+sC5eODZmrCR9tFFefi1d8AOtQG6HiyAu
iMQ/pZ8/IV2Lp7XQ4MzE0vl+/nGQq8Fq6LqLpVabjU77dkdDldHBiHiQIAZ3X8UD
S/IQjhzG8RJIHgQPj0+tTTg5rB3XyKSbQJ4mGlgVZ7DjeH3LFCL+IC/aXkrvhYrR
qHBxdMOKG1UxYPBYcIru5nttS9Ev5uco9IBGEBiVI3A4ab3a6G1nyOPU7lzMn7hu
i58jclcKCVV0kpXZmLDV7Nh+qzo1RcGD50TlUInKZ0h1Rsh0JsvMDCgxnIpgNge/
fB/tN0rxt5AL5kZNn4hn285k4MYDO9/9POM2x3Cs/F96TIGL7bSUULKl53iJLeEy
pEPecyvU7GamvakgV31Z89/7bOmADcpq8HmTfgTkmpEUGW06kpG70XlnfNAn6gcZ
BHhcyOcnDAqVCbX2XK1VbH3G5yM40BgfGr9AkpCjtTfb2h8dq8izwULQE/NCB1MX
N4iAc/m9ei4c1GW361RL8F3rJ+9onlN50vcZ2XoyOdW6hH1uQtMCVRDdh+Dcix3B
Lf3GMvvCz36hu9frABeY3NZ9Dd2q++j0t7kRTZ90dzDBTNZfq6IkDQ4v3k0kF4Zj
20TUZ4UYSJyI2ZuD87g1qOejW0nuYKPVPR9q8HDN2BuOe/0vdkppnHm/6wdy577o
pvWTy2soHJ93Kj5CB8HL/3RJjc1dxS0iIsy9+KOK/Tzh1wUV7CSHZ6rTtOvpfhol
lzJhK33HBmtYKlIDXaA7H7QcZQdDiOZ2IqJIdgO/BE+UGEDQvcGd4tZGVEehFc1J
4SRfRFUJ2FJyI8Au7bI5uXK2/zmuYPA9PGvRjZxC7HrZtmrPlEnrLh+HfCv7jBTO
KnFwVXpWGU8gDwb5H5YszdMHrp2yo5kgj+ftHP7jVtl0+L7Iu++52E7IM8IoC+zj
Q6hfgTQPDgM7URvRBvJh9XZobW9FXG278ryeslSgtz4heTG6fAAJ6Ib9J/RbY/jA
rrFLnLzt7x2e9BEPrgqNqznl7WRiROlpTjmPBcRVCT8Xcvd47QsrMKEaH4ijYIue
wigpf7IAUXHWa02c1BWG/Jn8o8BHKMD9cbxLFkgv+iJQgH7XdutZkLxLPr5J3hju
wyFmeD/iAm4hkL5k8tD8lqj9KT0PyaEFdr+3T/O80TkJUPHbmKB+ECTZGRwZnBxo
keJLFOczhh3szI9brCvMvZE5b8ZLTQ5eRrSIkfLy9LSZcDhUaOUmM7UfJksfJA3C
bXK3GRWcHlYmecRKOmwC2oH86FM2rA7m0H2dtr6v62xFJW25L40gEH9nCeAlj8j7
n6F1G5B7OOEqahjP7fxfuqW/vuDjrr2bfNbGHqHCroqnUwF6L7nyDT+PL6ck/Cz8
bngUhbMlgzm6EDRD3W7Wm6YRORsp+DzslK4NnpKkqh/YkZ69qpyIjHmItaL6i8ql
HGRFB9W8UFVU4SmjulJ1mPEu+p2II0i37KVLZUtE/6dogLtesWdqWHla7hj4iO+2
tERyjl44P+ACoGaKS/FiaZaKl8pOTKw1MxBo+E9V6DC2iDTwgO5RxYv2c0n55W17
xb4GPcUk3DFQT9qOQOn4Vhcyd7jBtMqLBQGrp7y9IaVuBjoJeQEglwKY7QmYTr1y
92clzCKOuRB7R/AQ2gj11ZOMnDM5yOCYccDyct8+k3gEfh9InChX0Ta0gQdS7Lls
zX5p4a8ThY9ApN2H5EXOW6EYmAwlsNguWAwugh+0msFsCuSDQDBj18RsAbb37PdO
PkHU3yStCPQD/B1sLHCofTECUAKA+4/AYzwBKSwzsIDqcnY+sTVs+Q/eedTz4kT9
PQXFffhSU49U+kBgwZW4IDj3mlK+hnm2xYQVBTymZqY0NbHXYW6qL5cypQI6S82+
f9/xf8h1ThbZh8uwPqQv94h8mYrCieVeaTQ6jRfiGO2jHUrnc+Qz1a+fWTEVIdNZ
/5azEufBnLPyrPv8cXUgCFbmPJni05eZIxwpnr8VtAv9skJocAxIs+fTdiUzPSW3
N3WN0zn4epoQMvC8iDMi1i/1wEDt9gt+dTtYdt0cxfyOf/+Q2JVdABQ33NMbq61Z
JS3he3GflLAUB62QPzJLPkph1t+zExWBsC6fzDhGireO31pox+dpEGly0Qb2iWZW
ZZ3spXUr7aJjNBwZtyI3h3lVAdZf8o7DywqSFuKc66JCQhrA2gDLg5rIQ9Aspmjd
a5cymgQOvA7yGwpefWILrfmR04RZtAHf0bayT0hYB2lHV7+mawHhzuFGtx1Q7ajb
Ulh3raLrLXbKtSwh6rgzbJDQ5ChDLnOSxab85rkPutz2DsPy89mtvQ9iP354F7Rh
QDHY1i9GEqeI9fwe8OgePNfIVZ83KB3TmdO5ysEG8ioRDft3QcOWiFLJ0AV2UBdo
gPVSyEZkUbWZwExJtYjf7S2I9IJ+KZFh7xJFSwZ8z2QnoeOkyfHYLMjiYIp1naBs
48xB9JAw64/yxb+HOylAe7UfM6ikIoiP3oRlrGl9WsiX4kY8n81l+Vdik+vZuRn7
woqw3V5e8eq4EUHq4RhXQMbluhhie6FNrCe7APBzlHe5OuX0JqLzTwCu72GOpSwd
2VjG9TkVTxktvd7vyYigiSWn5YlcV3iC8aBLZiRUc0Z2F8DdQjfWnt+8s/lTi/oH
V73z51SS1HbmUsJOarLYmi+W+kqfd5JauXcpG237dvIGm1LXifSowI/xukLK1rXN
OhnDA4R5ggt6Mo4G7Xos1VqUPJq+RpJK0DBnhViGDHD6vUL0WfW5ep/+F9NEPt1Q
SvoywJX8gTMhYEvXZgGWpJd6rue4u78gHXoRQgWCntM3ZrMizMen+VA1Z1Gb9sFX
E9QSy+jcig5aGFDscuT2MXqsY6POiu6RWr57bvxJKBLEzUnW0wsRtrJJR8Zb0MWR
bw/dHegjGpGmzXU7VHLlrY21ZBChJNMKgt+SG21N8ROCapzhL4yhrYELEG8iaibY
gNC9a389pOK9i2gdb7kH0H/UANKjdd78qc+ueQtVFN6vbkfwulcnNmEk3bHs6o2L
B8N8rgDquqmQUw4u5tUlOumWrC87bmnkJKCWPwopliiezBWNEVJW1bLO9f/vaSRs
inliuN5ExQwTyEgJP1vAdfjq0gOpJ5fgVScZLGC0ZnxrKIxXQd3OxWnsLxqwroIq
fyKXuj3Ml+ex/LxX1e4DmjZw1SVBxX6NbkixQwP32Ej+/nOS7o8n69X9gHxZ+mG+
cTwMc9nVaS2jlfGD8djdGGJemFKeCkgJVwXqVsdHvqIu9lgySh2rdpMitAWbeTzf
Bf1bsojAygvzcz25HvzEU4El4n3PDE3oLEJVuYnewyh1vL0w9dtmi9btkIB8NJkq
DAA7a7I9oiPIknllevHQ6heB+UIbZ8DP57LCj8vXEyrGEfSe5n8WptPtuq4ur3QS
EtsDBBW6wLN9+DCbW64V88/A/cgdJV/iEnQnJtfqCTsqv7Id9v4z+zYmA2OCEnUx
6RqVGoM0YjL4kkvO3lL2i8mZ+9bdunNVLCEd0RNgzAuoa2Ekn5B7gB/xzm/CI9Mq
WaQ2GoZZ9xAtWwyFb0Y6s8jvJRSi6L7mYcY7HC6GfOOzRuVc7aGXYqV7DgFEixYl
KfchyP67/5/AUE9hN9LvGHDZVjIdGCUgtxCnc0u6LgzVEqkd9Ng3djdfhilnxIbg
hDLGce5c6Adxg6jlJM469eTAV1Ku3Dm22F0p76DEeeEm+dJ5sD945U5auNejMkkG
ibLRzmCCJbDR5rdzLMAaJnsLOXluH57BptEFblHn/gowOrohcrPmJVzNHKLxO7Hh
XlcFwcyZfXi0CUTtvAP869LyurGJM88gpyw0RLb+CrOhyd0ugWzh7IuJ3evBDJlS
KFTiG0nKjI9N+UT5OmJaGOj8NIAAWktzARdLTHuTCndpRvJebfsS1Hq9BDFsz0fg
o6xeucCsC0taEA+Cn4AX45Ql6NntYGjoY+ICzcO5oMtfAon26rVrLNJwd6uaj6HI
rqEqlLhqrr49Jwd3ecBT4MXMpVCxiYz3aqCGJoInA9CnTRsXVKUwEaUGZTUndCHU
t/eh9afqIqhJgS5u2rczv9OHgaBg0/CM8BE2XAiEKZClw3DQbOfDIkSgcTHXBYAd
I57CLs08MzfMYNgAPxaHoDSFvIl9+pA+BOA68o8WV1fsclt38YTuil0fok+q4MZU
txLpJ+AnORaTwSnBERo4+QO5zSET5XazpM3yuPeP9ET2jXlFwKnqn9ILbV33AMcv
SFZQZsZDsYY93vPssOzRWTeDwmPRSMMEVHPBNvCx/SdVPZ5MDjLKHRPSaz8kZh6h
wE4iaf5/Xu1oZemj6YfWopsvErBzqcGRrnyJ/iplaUSoXvqKZD8FwqTY2eW6EIpb
ntFVQIpiaBUS0WrEd4nQbrTvlr6zrK3oQ6pA4h3mNAz+KOtyQP+rChkRSHIM3GrG
Q5Dx+uz6IX79Mx2lfU7rTrgr+ATUQrhNixSPMj5ZBdt8dlgd5lnuQsXM728twbLy
ZBzMI2xunVcHh+JyCWeWG6kfQdBg5hY3tPxOIutg9jR4GDb7g0CIhGv9vG9I8Xjg
J0N0BKuSigQ3EAkqvNmppnvWbZxcJGjYMOF4rGvWfIsk4SkiUwq1nnmpoIIWTmD+
6xGMGvbi0chi94sbOt9PS9tBsbWt6jVmPAKWoMIsn+HAhtWoy0HqKKlC9ShjRAvW
1h95mksZn4BCo4daaqW4gDdp1bzpge574CAlpCjfeLNznaZndLNUZa/hT4KbKGXp
KbgoRPS7azywmowDP2hYIBOoSb/9/0DoxHoB9u+vaNwYT5ScNhsAbjVoIWatvVjx
dPDMg1ANZzVKmrfyFAHctye2VqOz4ddH8rq/I5fOUFniAK8rSoLlvOZ8T2WfnbLM
tU3Y71y9Bv8aBr1rjEM3X5uNd+y6biyWDQCb9UNtqGmymXOYgFTNvuO1LMv0l6ez
s5jt2YKD/5uirN+1vPTWNJroDWeHPsCx/JtLqm1ozE1O8hfJCY65d/q+7NeZrVrw
Lojq5Hly/rjvrvk9rCOWrZFWRXHm6B2b/lM+2k24K6NLZsPAI0HS2khQmSjk8F3y
7X7vIyu9uuQ994jj7i+lRo0RX6mDQ6v6jtZ2xTO7s6KKK7UIeLi9JlFRp8/oMLC6
/WUvf3a/+IYTMipMvI0AIT1YkxHVJJ3bXERMPIS28cjLY/Mkuya37fKJNlPZKTB8
dL5VfMDh+EWPEI7mNahqS3iUNHnkF1xwPGFfGAZO0TUFWCe9g1w2IfxyprIKHtGQ
3q18vB50pe52T5WEBunyfnzy3ELRmK/pu/Y6fRh5UqqV7p78BpY6fVrCHqXc2h3H
gY4l1iMtWFkGJ+06eQ1nY7gJk7W6hO4Ph7VCNcCo+jPliJ7/emQsRBhU3PDPXLsf
2g3A48X5eJzzcv4sf4PkKpz2JtdujdrOXZKvb7UP/0huRUCixDPfkUex+5FdmuYS
9N5erSd9YCIjVdgsRr8OZft3itmMqMy1LkWASyORoDk6UYRJB/S47f6LskaCdg2X
C6Him/zGsynqAGHwfZwpCbRuEOt550sMC7Pas8xeUCwJ3klJ97hNvH8stlaYLwuR
Av3B6T4cQCnPPdFk3OMmEDg0PXOz+QXTUWwu3L7myFdlhJ9kI41g2v+puy/73pLA
w+sLkAKENzb+6Qbi8CWI7z/d1a1HggLkN+ye5q/w7r11NkF3JMgMPg7tcfD/reOF
H6hSFZ6Ar4JhMLu7X38D10KYvd5S2W7LtBSuoJp9zdTT3OPywMge1RULCP9YrVp2
p/FCKA2PuWcreNFW0ACDyw8v89YXBS7sWHnFwc3JXuenhUVHywG9Ug9GXyjBDvFV
RHVlpP02dh76OEQbZFNvvyktKCbaQpp1YQL0GvjR4XUJ8dgbibzlcRrarOlEwVxW
dHK9IEXA5Ua8Io1JT27PiwoKDTepbbr3UQs/iGTdbtTZ6kcXf/cNjly+3RGZaYRv
Rs4N67v1qdjCNOGEZoTJn9rsqFUSUltnhknDx84Sb9xhpu8xo9DunLLRZyDnVjJo
lyYlkaNu96iR6UMcai8NkaS+4hnWKaEFASUt76fQMOrkDr0P9E1ZFPn89MPxDkOH
EtGmXoVOyg+q2/vlLMyCc/BFxOUZPHz1pv+ekZXNzeBRmET2x8QG+rzW1H+RUhwH
jDflhDKFdwp8FdzUnoMHMiVPqdYby7mJ3sY5Fj+j/Mrt8ssROWKJvLhl/Mdxxhn4
cuwYigzBxf19f6bRoHD9IAlMn0bfwbfksIo7M016QiF3bSQdBskmxFG4hMthNVCK
d09sSGh4u8aaQnikDNA7MS+f+c5zRy+8UKDqg2T8ZFhyblJ9r4D/uN+LeMptCfQy
AYSv9bSMNCWzHRI4/0ANAG5nNn3pDKCtTVmZ4wT1RhRGLTSb43UylyFNGuzpkUu5
CNZz4upOBJ43uvrsUobB1rrNSDWikRcQHphn+BCMWvxv2VxGeMVDxX9jBnbGkFC0
PH40vL5xTMuIRkeep0a4LvfcU3BaWnh25cy8VoG4qsF+iGKyuyPLRpBMB1+YRFKX
srXKdA9fyYBdspNFih0lRkurZj2kOg/VN58D/3UOc1wQz2KENSSZhVRtCh27fbiH
PDjLyn9VuXlHLo4D55epvhq9AYr0jQn1LLvO5PVpGN+xy0sJEoVkd4qYf/+DA6gb
1sZ2d/zx6BkX4SD6l9/t8YuXV1cTkBJZy40dXRnsa22AAqewlGUzryN49cNisG5t
IhUz8evMkJRX99m1bGMGMO2FAlH6snw/HB0i41dsoo+Q5e/FivhiV8X9sg3LkG2+
Kc8oLYEoAib/MLTpYs0Pf/KSTdIrU5XOIuDlsUNOAPTdFfcY5PFE/ax3lDiHuF7Q
UauOZeky5sOccEPMV2yEmI9AhVOjhSfYApqrIKfBuzJe9nBWjFcb12nYOv7JhQNF
vz07LGsvn1JcZFq+fQzwDoBMF+ra5nPtr69oYOLb+oW5uNVKhFGP+GW0rlEj32iU
kcVoRAZ6uXNY/BSVtFwk4QQvDkYJLzLAAHDTDLcaC8NOk7vGLYuMlHIgb93J73pX
cSoNzAwu/tVHIssAJShSPxfHsWr4q5uGz5TQpQdHgPMTurCX9v0gSSrkCBN+ofyf
pBMRiz93HktjS9pTrkQ4vTLUhQK5NgZVhmDA/AarICWfx+dZYNsqZB3qE1/jNcJq
uhREH1zr2MPg2jT8N19W9VUenfyw3uLTnjVwCmKdUVXLZ7+Ml8w18NQ4w2G6/fmg
cGwC3zP/iz/SV0tuZpp0as3gWhUKMRd2pKWxthnZ/BgIBoA75YbPoysQcnKvMelh
Gz/625yQAr4WnbA9d+U/76iVWdRW09NYIBvtqkgvDqLqDXWvm9gSS7SrO90UAV8N
LPDn8f5CtQjne1xNwz/bHUjYvd6yEJDjjmshqgCy7QWeW4j43lLCiwG2JagEuuDj
7s6qkHFOx8iEL4N6D6Wnk7jHfA3mqRiv4uXHHL4oBPWUb5OLr3X+M9hqFe9aysQ6
Cs3WTgjc9qBohR8Y3F3yAi5IWclKqsQa1xpXnuinw7/uLNJnyo5GJgk8hk9snQ3o
eQXoPXnGh0AL+6fbgjj0Xltcp74Diu7NvkCIzJY7D0kwPTEGLUue1/qSmbP20KfJ
07WZRX0cMX7mWhJY3yxg0pb8fOpdPluO1fTevVgx/0/L2aYWx0fUx7DEH/M84LsS
975pdyZopO0hurUwEcZqoI/nfsTZDO+hE3FdTEfIastpd4iNmldJnsmjCwKYIz+q
FuYK/83BYdBREtAtcI/SWqsLHR2/jDLVjghiMPjhF5AtanVaI+wiIe6IjUUmg/eF
BgykMNT4EmZfakGH1KvwyBsy/rniNlBozwAT3xw/su1EJG4FgrV9mGRQ5UyE1fkS
3PLL98T35LJeAi1HSLYs3otrAscL2q0nzeYvwEZNqdiAc2TOkAuAfRG32ffxde8A
wLMCxdIi9oZqoT6exBNy5jmBLubRA+s1Tx+B5rtWBad3R1JfxXY2dT2FSR6YbBI2
ETxyzfYl9E5A4nS75PWKyxERAsIFW/+OiNUNt0uJpaKz92kX3qkaF5XQDl+vgLzx
96alLmYU0FbFAgjOBnMaJhmUN8/KMLpgpQeUmy0jGvl9TXWwg2I/171feAKeCY3h
sCqsxs4lrSwTOwFu1BMXxWK7/irRdEUT/uwlDYFkOFck/R13DNbRd1mSWZuH+fCH
PP+FujuV6uUOga5QZ3BzqmmWIjWKHBRJ+kZwXg4aVywmob7O4ttzvg7vh61w3XV1
Ak7NO7ZjEKsccysHEbY6oLNPhpjNwGvSVuVlrIjQQ3JhvTzG19QXjEVURkfieNr+
jnhQyKAVwOMG/zBWPuoHEZVaZCgUmYITtP5nAeAG/jSaV16H9XhvIfuXhR5V1Ass
sr/aOnwXGaq0O7LKxyQKdzgQ1ldiApa6nTxVi6NX5Z0ZDtEgVbnPd5dX48wcJ0Br
tPXtZiOCOXOHtxVSN08QAoSGHerTtFGKtGT1REjpbLYN2McPPpD6fpBY4Q9YWYhP
IrgDjl3MXgv/15tp46oFXGfgqMU+YJ7HdQGN+nGbcjcLmheh2CgPnDUpcjZmOCIc
KwMZl50OqthTvz9Wa9rot8RDLWqkWygc0/k8r4k/0zKyU2k2eDvlHedP9qjbH6OX
vUPMka0pkq9bdQKTrZS0T2yW3frC3P7QYsolb6S8FX3bW+8Ghcg2Nb79wckVSL2z
JzW0ivcje84PeKJOtNYIMvZnUKlDduGlFRdCW4NnAknfgVmssd0DVy0vkK7GXILW
+23hmJDPXlELas5i1YsS/l8uQZsTMD5VgnSoZpprLFA81FwqgiRNzNwp11uGcPjB
P7Fd4YlLwIyy2zVMRATE5IH7pf6UDbVki++LwE1nW7KYZszwsepb6HrjXtZdaEmb
xG0L5Tirz1EGXee+ll2iVzr5nsi8NLrRS3TrUOU0QZbU4w7vaNSjr+7dWQMz0w8o
2hscqKLkgueo5fumbozd87IBdwgxG0ZLU/itApoyZ1pBWHNSqyQKsYzAdjXnqOKQ
XVuXAXCl/H8mne6Ec/stfKyNR/Km7LEwxbpR6nnml7t4W9wvO4oSX/HkrjgGLZAc
AAD931JS8uk/u9TUCIkvIoFcQa5ATdIuyvGg/uwUUl4BxiQtEuCZ2CiKu3n3FJhx
8aF+hAFp5ooMMqGm5oX0JJI8I02Bbbd2WpMd/7vwBfde+9e40SjN0EuNSiYs9wxw
7KDJWSro8iWZeXAeY+uQQZqqz2Ivt1wMUq8gCVMHfxYx0kripBH7ECZUCfteHoX8
EZXsFO/Hsc4DG5j2AfrKmEah9J9eAUsCewIwvTyqv7jo+rmvKiW4lFpbYqZ07i1z
qoccpQqcVe+mgmPHpzNkQJ5qIo9u9a5QEmEl72+fGID0FcL661GpdrS2I5QfeAR5
8EsU3FqiBjuPrhGD83MVAv7vLkrCAcqMCFRSudcQ6/CJr1h0kDpYvjl7IdMkGLWJ
4ghFQPDya8Q+korZV0vRegklshGGgumFMpy8ZIRnLt6aw2aGn4+u71QXdMd0Dtjz
Y7FgdY87pHWgyHAC/wj7qIe+UXS0/tKoCUfvvNzhx+BX1gVetRFC/yQTzu5f8+b6
1Oo9q3pMalT8wNXCaxUGaj7jcD3f0SrR1WpbrTIcGFXFlW4ZCxviYtzO3SU66iqN
zU/PD31aZ7NoG2zXMJ0G8nZZ7r2zFgigEvUr8C1fOtj2J4l43f45+eA4LzZyw4Yk
wo1beFASgF5PtSedfRq0cYy9jUOanLBNZKkV48Vpax9fs0o8WVZzhfbWp86Ayqw8
YM4IVZr6pNU2n0GfnHBXI8jBdyeT0gJKNil5DPY+zsm6HkGIdd0X/s4Bpn2eg45q
0zra/TIxo/L059hrWvFdts+xfu8nG7VZMVzzpRUd/QZqO2vBl6kTr1wsPbg4xOfO
8PWpAa4BkDJzlDlpAgqVKVDL0ZUTivKspujLfzIk5jXkqWJ5OmLOig/6HLTedBvZ
5VGRKd8VzVVyxsL01kz0dV1nCax7vROlxc/ycafEdbyzkBFFWkMDR7gu2kAcoDI/
jXNTdgZ1XcnfAAq044vXcVO1NejsjyqS0rbAPMnzEssszoQnWg4dfXXa/CgSbYtP
aHJmdbPpYcaDM1v8DovDhULbgYgtu5VE03hMvwj3OJZm5uJE+18trjawuY5W6iXu
91EvQUv2MiZ6WEpJxE5ucV3dC8mEdsEOpqkRJkRjYna2yo4CkAJWP2sC40r/thSK
3REdOI42S/DVfOuOxfPvN0S6Rh2EspAEo+GPYTeKkLOFLQRe+SvlmHh4kbCMplQI
qwCj0Kyti0v2F2S2n7Hau6L4S3KtMJIBdqSxDxy8L+clKYyOVRdD8zmAnLPJZ6nr
c1WhvGJLoci7JLsF/mZeJVEciPhquxeInLpTVWxzoa4BmdxgoPYfVnv+pp3a9ukR
42tSTGsVXu2ctfR80Q98Z8MCAHDwHOrPxFRGqBTKznNMH8M9azOjfefgkzIUTpTy
yBGjhkVCr3j8F9fEwl1d6BNN9YBYbt3mGTXtJbcN7RMGg/ib27E4dCqBbNelQAAI
vB1xMscLRP7DYnCzRRW2J0ujKClfxU3X6LkIJQbvUVfWsNeX8L5rjCwrW59K+epD
+HUtMc6KydPEvQLEkzfDn7+9iQFUSOY4c7GFJo2VrsQ/jBkch5xiZtoLkEnyeVoV
N0fW7gzZnK7S00jUwseM+nm7PAFAzLevTL0X98t7ItpZsZ0UNZbtJg0EzB9wqIY8
ti6u4TJCdvITxMqtzGMl9nVPXbOk7DPJdti07VpsbvKBOczkTDr94MuCf56BXuoT
unCIKgxxyCRp6xhja2//JIOX+B4GpQNJfvGjyOU2+TvvBvOEMosEO259dYoyYS9+
7tMfN27jxb1UGXbbZu+X4x/1rPd7ErF2lIQXFZ3+G/hYD+3g/u3/wK5dhomblcV5
hrx4+1bU6sEB5pRxUqStECN2DcTXCQmHLVXjzCaeAaUKjUWIwBdUxXPO0mktCWz2
VutJRgjefmpjlbRdFue2EzaP/5B2at/Ge1J0CrOFd64FD08HqeqFRbCriG+1UuCU
8J7M5WqoADPMsDXdVZWJ2bBjW8w1ac4kCKAfpqO6t8wqqApp6LmR0C+oh7Fr1KB4
UT1Iiwg2iDMxcncnlweM9M6MnlYIxIP4XrfhaXbpzLXsB3myJp4wmiRBT7LIyPwc
JxZQJnDzENL1vRcr1wF+OgThza5GvD4pfUWW6g/eBgBE+bG7fUGwWdjZaAe1ZoH2
42pWHQQt3POVOkC+WjaLiYng6QPF3aiZTxF+gUeqD7Sv85QdAN4oz/uo+7TbvSKU
ug/+4yodP6Pj6EvP+1IN/krRxbwhP+4gHMeSnFxirm51aBFiRB+IRvjf+yeFwT1n
BhApaYBP80TMKWzMTSfFjITYhWKvdcLbrBparskcA0kLXo1VpheipRNYv5AnWNT/
0AI/1ZHLAaIJPTDqnbEvBKy+8BtB1a3fhht/TNh8RejwFwxeYg+FlDm53Sa0dZrA
9Q6FhFsQLgCHI642nTBLbfozKYhZvwUCy2gl1EGasrH5Yl7RhJL8dpbV8XsqhXZd
YNH+hCudqL5SGJfZfTkMaj27LqmkYAEXZpto8g3GrgGxfgGSWVJqfro+HGFGmFEd
Dl/r3Ib0io/W8ZBE6wXWZIsXgSt8zRcQZJRHkNKufZlNcdY7fZbRO7LUB/rfYu7x
2VXGwrRQfjeKM6CI41lO+K9fzsAL2ngRIwKkwF4WWeWYcp9TRc2ktluuYNYNPn65
b334R7k8OQbW2BpAZ1OwpdcAAeJ9mdBqFtz5Zi0KyJc3TE0Sg9/IFWu7u6izXgvA
ix/ESsbfx3ntb1K+XfugPDg2SgLMn+VwJtdYywMTXhnHAodaqLVrLOsS6u4oURT7
rLS9Nfk3oBDPMo0pNRuCrsbHfYu9gn4FW7J+esPGMHcphrnDHJy2JyhKjsi8tEac
JjHvfCsSWhWQprSsl/+5LWtoBBeg6t2jObOxVATUbOHXAQO5b7TROLkK/o5H/w+H
ycHr9x1YogX5l8Y3CKDZWAjHrLVUzFv5L0PM43ZetzExQvJLMAyjURgebijFPc6V
Epo+kvKTDaxhWWLJDXuEEu9qCRUFDWo2GVv6H/SL5AELBgA5ztQt4yFMnc40z9+e
gMuPyziZOMAStK0m4196WgUFAhKRxoFz9K8JEGRPnGgGOLYb1tBOawx8fB9F/aTX
sHtQclIjoDobFVF5z5UuCh8e31Yk2RwH8LTHFDxOjPSk6GgVH4iWUkgX7uWPzfWS
O7h746J3QFiOQqMqOdrkKc9cxIPyKbdhCBDbEllnmZ5mR+77Qeq/kPMMfFSzmH94
Aeah3Wunz40O++00KX0KHVrInZmPd4mR4703uE2nXcc/Ld5o7dcSKE7ZPi7zM6Ot
UzfDriOwR+QyMGQ9+MepLC7yCuE3x651ZfCwpp0rOdYYywbrk7KvAKRAW6VsOsUx
0qStshkhP/KpJxQKnhoMgo6380V/3d27oQTAscCMzFqytvodvBY/oiaqarn55gyM
vSoZl1InGDfTjNJm5T+Iyvqv3zelIrYGYx6/tIunmVX2QFleVCHC21QPUU225C73
MbiF8TdgellGc3u8QAVep16BnDj0limdGWaU4bdoGg7yI2tjX4ZXNMrk9qpYKtVE
pxJLUVgrP8G1BA3a1RDMXATnes064xJHUNYUSw+R/UJt8J9F2FT20kuoDuvzM7Jf
smcV3O+pfDJPJ5nV0Biz0LOwrH2WY0atxfDymvjlXLvw6s7WdnJZH0chzS6k1t9W
AgVMTPo2pRPcPzjspCJ620ecWn+8SndHeRrmKR51fYQn6bxaGPtRgI+crGNoJF4R
SDFzRsVt1Ety+f5FpesFamI6UXd43q1cZ0PJ36GZgeziN2qzyq41aaUN+UibC1q+
EJ3RLJei+pZq+RZTtj+pL14YuxIwJpb467uo2QOi97vZ4IsDVZXahRC+qFvcQHrn
2Q5mm9dCKo/PlRkLcmtO2CgTzpied79FE/E/ErGnGFXxVt5Tuktv0iz44DO/7GSq
kc9ESG/cAjTWwZm3EkDt0stXBhTeC0Yr/OamI8q7qrSDHWXPlP34qNe/AN3pku/c
1tojgfxEW9zXoU/d5VkpCFE+HVsYfC8pdnjDLM4ETyjTuETDX4sElOJ1QueWIu/T
IKtee2WqnHVzNpKf1zzAeZL7YCdNwUf6Y+tE/YQyJSKjZgKL6DMsPe9RhiBf8sIL
Aiwh01lFPLK32UfT/zmOsq3nzqeMLyrbHZedo9SDeyXGpAwhOCk4+5xT9mFF8I6O
fTsIXRCWH/ygUPHjmk3yahvDh1P+Sc2+dOgymsAPYVskXnId9ZjbhtNvS4qID0ea
HSHAd9caL0xuq2cou9Z6zKKNvqtl8GjmzkOiDK22W06gGkrN+OpVhWvOJjq5/2FU
9mo/QHiE59hDZNSg/8eLKmIcp6BrDqPbsSN/ncb54SESEIgDhpJjE9Wz6P5vYzQp
1yrrFyJIjtOtwWVHdMIuW1z9VBW45WIdbFqt9h3USiHu8L7EHb3Kr37zSw3BGPNT
zWzYrgeYX9NeypJZXIlP+kW2UjiJPcgzRQT86u0P6EFjZh44qPHKhBno2Q1OAynR
kOpBLhwx06xpHyWBwdxnibeub3Aa6pxBhaLu+WoaFX8PnwEp1GnuWefZTcmMGbhG
knGGAruGPltXSqShj3UWOuvrIeNyyaVuNKIGd+BimWA06mDP2ZRAlcgtAKel4b+l
AvFUSMepqs8nW1uauKx8eWeo7t2nQONBwaZuI3n+U9qCXREVGeDyWH6ZZ8Bwa7Uy
S3b6Vej+sK106ux/Tmi+tGcJOageB/0+QUGwUgfuf/6vLVoMwWjLPVmgDjF5fEk+
qTQ1R6hewft7is5gqF/cFwtssbkR4Sfp/LKR4zzBqVJFK3nJbT/NuEAG/wz3N+YX
3gfWgRM4O5rKqivOtSvPxybf7L1KZRRqrt7waFE469kSfkN09RXmXHP0zwPRgnJk
nv+EqUAdRi2+BqPcnmhwl2qRk/RG3awHWuDThqY62h1WsX7L9Ynstedd+Db3hzLr
qu4BjaJflU63Q1qfWh40c/0KvCAmf8rc7gJIZzguuZ2wbhoGkgzNudGhCInsSo+L
gJzeIBe8gSAR7xmxO5ob23xx4rIlC+JFptVZ9yZSU8myHx2XU3a+aM/Zzr0EPp/m
neuTjWOTTMgB/hnC1FGQkFvEJVpnElY+41Ne6132BhIcMY0BOTgLo0Te/xcE3yxD
dytyXAnH9hhmLEqSDV65/Ft2ApZXwQr5BAXeRHrxd9kApB/0ctJBMfPNx1xT7ABD
u02xTSWOXortob3XVl5sc8vH9YzJF3kDn7dIytdJouwHIf8MvN1Ndnc5HWoYk0zz
+LpL0w86X2g8/kyF+uvrg5okst1SJ6JxnTnFb76/TSIPbWesdg12OPUByjYW+h0G
VmWiGBpo49zfbO3KeCIBbEUQuc75ZFXEfD9ONSnFK9baKTYVX4yWQgu2heE8FmkH
GzWxuY5yO2uqNQeNuzrEuDSjqQjms7HA76aX9yEERqH8uRtTadJBWZ69CwFe6ycU
oVVoJDnDmBZIvsbMgLebrsv3NPVytJV4QIKCNjTzMkbSMD1FAGRGjAxBKT9HQ8VN
unDdjjSROcylMVbh8NeL3ywNbg+RrhCbNQ9oUY6DhMk7UlMJkHl9rJf7ngrMvuYJ
equmF7DrCR12aCc+5tOtQp2nQbF/QYQbOUmhwcLoT8VptDnLzjcYSkgQR2hmvPuT
TZ3ag3tUXFgnu9uxzL8tPMss3rBA9Gj+ovKhTRHkEKbftxCaRMKJv2UIk+gzvJBQ
MUqXCj4ADeus27m265VxTrtbDsoz9bLOBfMHeKJHvNnFLyW9gJFu8CI4Z446utkV
kD7KhS3xzB3oBU51YuGhhJWPswV3Gfgc0+AcBnOfQ4EfzYLHUcYofaXY8+mS/iTM
KEqsGrDR7ZSQNtapko7TLDvclGa8uCOF0sCrhY4gLGytvU/f8GHSI2AGEjEj8WQk
uRfOgPLHXBUAU+93GcaPEFvEey/zsuX/DPTlTdjYkQP+pc7QeaCahB2CFwHJ7cup
Xl/wndwoNp9h31J1Zlgfd21t0JWWayPP2Pf61cEjeAsSwawH7Lw8vR2lGoyTVdao
gg1t2j6KAgQ4W0hGjqROKMQniKrvrtKJ5uakJmlSkxfqoYz+UFcZZPALv6fdKmCD
nDCtVjszeRWGeVxkXnM8VMJjOGDCSsZjLtyWbStNqPD16rUF29F7CIkm51c823Ut
cyZcngtI0Frdm3hRDUZP7td3auj7INg7VVNaG7NlzfIAEuSu968ZtTK4QCRS11XP
mbN/L8toMoshb+PYKWPsCELk+vSKRX1WgH4t5GOwJFmrWWDOy7CzcYS2d/LK7pfq
QQZrEKviw4FRHOruxmVRPCj12BJq2r89vF7xgyEnntWczHlnEoPJiyZO8ta1qRol
fBnq+tsylIUVMVMOSLH5loq6dBMaQ01JlhLGlcyfBzBXNq/LFmICgcu2jtEQAiqO
Se5fX+m2AxbCyeYt1bqH6dtFYBk9bSicOqKL2werY21wcIewhXbX5S2A/PbZDBAm
wtfJCau0xgQHOlJPZBdyoO5H2irZ7HLgjbdVWVhH9ulODvlfOToO6OXAvZYGfzrO
JdJjXgAAxlNodeHiwYYnBv38Y+JZJkRhQ3LNzmict3oT0rucqun4Bz6pi9mm/rtq
r6iJZgzcFZCMj+ylUKaMsdbb061QbsNbFI62n1JL9D/OT6VTLsyvXXjIG+FTVF2s
w50IO0TQ+9YZHncFlqDK75h+HmGh1IjdZ1RIjgK9W5AlY8qgy4jgSoBpMhJC4Wmy
Pxk20G84rKuA6ruxcw0LAhu92v0oZtzURQfcldpCcrF+LEhvZEdcmge1mvk0+zWt
PltDFgp/mkYG31kUoAYlHeIi2D2K9/Pk/U1fxULw/0wFHQBBH1tStS+jHDzSVYVL
4xRpLThDPz3T+kAQFbMi9h0CiQ8O0m36Yy1zfbJNhWEZqLSEM8SWCKBFrrwh7FZ+
MADv2uZehGeWMFny3oh4Hs+HLIIf+l5n4guB1ikCp7GxGApNzIlW0R8FfdSnjaVk
PS9xj0ozudljF1dUPyYA2b7ZuGoL1cXdNquaefmUN4yCFyVwKRIWqXiCgJCnD9vm
1nBMoHzxKlvGTR1kW5H8sTZ8MFOF10uwQ3psRzkKMQ8lZcwqk2w+aWXWSHcvQu+G
HmXFSKZ10p4HPm40E8H0BoUibFL2bFEVaQWAa6P4swStKVp3kq6tinwsRgyW1oea
M/Bu2VdcyBOKCzs8ctqEkTtk2bo8X5WYLrmK6eecxfs11fzXJWK9D3eDqEYFY5Up
s8c0THYMIVx7HmLRlVsn4K22BKMfnw/eV5FgnzjcHkXN+LhDCps2hs9J7+1UsNdF
tHfVsXqyLLOYePnLJoUfgeyvFOcS9YGKu5P1hCuNjqleTplMC7j8F1gl0lOounEd
QOQeMKciaSRsvjNT+I6tq9nGZJNzAhNTMIeR6NEFmLosXM2xWpo5tcKv+Nu9ht/r
MKqgLFwqirq/5M2+uC2Ioj9LyCeXpoZDD8VbPtmsFL+fJTIhBtRyZJvbWILHplKY
DVHmQMfhxA7/59e4abC0JBWmGhSK6nbtsUb8tTGuvBYVznM69Pg8JwKfCU5K5X83
HEQ3Rkze7ND062z8zwoGuivgIZ+4gyoFaw9hvWY+Gu/Q4vhUVjO1p6zoQ4K2KVdJ
3vqAkHzupRV5opaBR5qDLeklRQJ/UbSTZ5ikogoIDBUad0oY9vmo8My4eeui0qD8
y/NpW5JW20G1ug/1GZ7AHCk1tcdJSgEVxO8j3ykbSHgOu8RSM+kL85N8vxJnr6BY
aCFjKgpTMDms87BB1kVfXzFU2NQ/gUlG19QIPXQ7YCsLHAaBmg42yoZc14uMgAHw
Q0iHPpGFEeynwR7zuYxMceRNAxTPgrTYAUZ/pKJ7LLEL8+c7/vZ/qub3LfgHV3K3
ews/NIr0lr+J634+zpAq7Apq/Qt5RvDUrpwAaxdShx+cwaleUv2sgffaALkfxfg6
lwFRCuZiRFb8FlCoB1V46YDVFOtYf4Yzy8ez1XYMognVD8BE5vu4UnQSPIK5Dtay
YWiyZ5HHo4vsvbs1ie5MPf1BPWj3gu26LFIWTb4JnGCKJOtezok78hR25Hp6VH+j
T9+U5TKbEFglUoP6U3sYHDpEK0C8ANz3781oulxf7swE+ROZEx7t6xzRrlL2tpkc
OcPKr3LM+3KzMoDq2z1MrNRMuWcYuERCU5PsTUWvW1Lp59+s9R3Ll5GNl6K9APJu
nQVRGi/m/uYbfe4sdUGD187sTS0pxPXggKtJFVaZn40QDH8OWV8oPXuvZitBZhxr
rFUGWMqnnXZNJULcEEpoiMWZK0uhzRbkvcEhB2XFFHS0zaYnQYfZWbv8RoCikddk
tqPuW1WwhvK/NZHdHorLGli9Wa6gIfMDBkL2paQvs6uTmtIT5ntEnqzSyWPVEtXh
WkuypqCuSBxC3EC9fVPbH1Fwk7AYn/3KAtGXcpKfqEeAvw0lXrGYUcIYnkw1+N2E
SgipS6EjAHDay4ajuQZgz97aQHmmpTx4hNuzW6LYm2qtiSYHlGO+gIPpFa+l/3fQ
BetR8Lj4heJLK5wKqIf6GWrf3e7a3DcsloIJXFecEtZMhcwkzMgW71R+zrnLbLy/
zrqxqzRsCWjAzWfI+ec00czXw9/OcegqbNktJ+9Hx9az/gtRguUL1Co/XEK6KCfZ
T7xhXeIRgPNWvwnVlGoOCuhn0clZL+QC/D/cBQV9DXEadXUGYbhYEQgdyHDtikam
a9/8FwbbyYYLg6XfLVEdclDzC6EBU6eGGlDnwg7iOs5X9HFHKBJJk3eAeh2md4bm
caEGhvDJZmYMivgp6cbG/H5KWGDImQ08Z7rXHcPSGYpi+vx1dpwTVm0lA2FxYBru
49QX5rob1gv0h1q83ngL34mhCvvn1Szuw52f1LRrj3gLQ72dJ1VsjGewr+qoLJdK
Slt7OJKGCabAmaVBgBQHEeDUVQDuHLkfIWE8hEstsucqcNGKNYAINcKt1sFcfxze
30hDj1YNdvceJmKEIbxynC1R/SPbSjCy0BDyvg3cNJvR++mhK1yK5tPJ6gX0Wj5K
016Dz+lRl7GsYX9j8nofLSzo2JkEpqE6dNeazTZs3iSvJusq6g6aVqMb2tdfq6Cy
LqoQ9bzOMqlI4qHZSQDwLudTwWwfhgSoMuJThkWphwJ/zXPZ+UBGVkDZbZVRe7/F
ljTHXAnzGMhhmqzx3QuE5pYCL7GAclasPZ7WhSc0Gcmv/Hxt9H+VdtMjooI8Pu4H
dJWz8zRiUer+R0GEHelP9387W7KXxELMRtoghkZurp7IUXoQpY+7HyQFgE4r612b
huYXTplC25nAs2hQlQdjnasd45FtmHvUHIhfU4zhWcXX7UBoXkVhrE/wgTKjTRlu
92XodG7vghwIAcDcp4rXefpwuSIYkjW1Y5XNX/zuXniCWFeyFKwekOKDOFHfW3SA
OIKXzTducUVyTB04RMAib3UFdodwDSOHBHeamZ13ERFmz/pGlpzpISL2QUHi5hVz
XrQl3k7gT4wTtvakWPsJilAnJv5iu0/3DzsXKKVuWZNtRw5XyIq8M+tXGmXvQ+Uw
KnVwt6eRHiQR4+TNOlRWQqmNeVonAJi1CF6I4whE1g2YWFafMYV78K9JbBWwkU5q
8DzTjOHzkPAXR4w9HScSMWLraTbvkLJCxzXPmNcdYPT14l0zKCmq+BKi6ND/Oe/8
qeTuoxQC41IFzbhTvOOxRV/PbRV5vSwWAE4Vf354yGZxGjR5D+u0SvApn3aUaISZ
a2bFoXRxXcav6LtV2Vqv9l1Z5ISf2cdpzyfnEkw7WT6lyYQMcv0lTtk3kIFDAbNQ
4o5tAMzbsop1ikKGJRZzcu+o/Gh8pib0JRyjq0VCE2JKtTtyHVQhw5k5I5dVrfgU
BobLbgvd1uzMYpDjz97owWTKmz5iC+WaKfRyDc5z8g9UdVpyj53u8og4O/eCiFU0
3uLM6kLBqn9apSv+vOToBE+5A6Uo2+Qrnzq8fAvFU+5OgmA8WbV3Yyl8/pLBRL5h
T4Q5PLqejVyv4bYSSuxX6yaDc2qjBH+VgwtAgHGc2zl9qlxV6ywFJOUE1eSBNRoM
ke0hrzZFfWJv16zN0f/2WHvBysI0DCZJVCRp4W+2LyjsA6GFaqKTjMzsVHMUBlw5
8mMixPrN6H0QB8AXp3A4RtVMvRakrfdezXIkjTtss4yx+fn9+N5+k08zdh9HxeCP
LsV2HBCqXoGn02arrL+kB0sOACv4tEKpazKlCxf7lSreEybIItpPF4K3d8s+JSnJ
k58g8v9ohcXy7tGGOzhC1+EieV1xe0wnHX5e2a39m8HXpIQNoFwxeL5nxvV85kqM
/DxRdQQeiECNgic8mZqEFDlv6FN+43Qxk+yeRCcVFgt6neBlE6l7p7+tieyiYZp9
KHQJYQZGe8EbBniePJZ0p4GQweMvetN/kaaOmne4RbO9atyoqT/ZhGeNrp6y5dul
xQ7m78QlwCPQ/xMqyKuD2gkkt8g0Snp4XHqD9kbDJjPKhteXZv9ssKBTt4Su2Rl3
n3tn0GCpHEUeaFXtQaCwSJ51iUBVNcEPWMX2Rz56rJOYgI7lnrPAi97E+FXoY1s/
p8SdwYgKTWUYw4bXE5V/Ns1R5WUtJJyW75tCTBfJzMHPYmlT7ssu2F3j0+FmeJbd
z+qswf+XyCxoOI667fieAQ1U5Ud08PueSmiXZODhqge3IeJ0MlK5VR2PHcIubERT
AFdunERmv2tstDZy0gsSFw0HOV2uFlSWUGYhIcLRzcTuzU1vLg9edzkf5wnbzm5M
cSKq7jY9ZKecG1Fe7wzv53Ub9Qqvm0V/Ldwd21WtW+va95UpRa6XGA6DzYyWAX6R
0idc0jgJs7JlzHBg3n6kYfkWCfCN5eBXRkkts52ooV4Al6PKEL5yCyGa3NUWovwn
3DD2f5sSJ4ff3h+pz8+9Owmmy1GUtnX8S29I9y2UPYkj5smvoDRk22TdokE1vWpa
xXZnbAnteILiamC5jWkDseYssrG3QCT3+VcjRlq1Z2RzJpScyEg8sxo/AmzZ1AFk
dcfSYtFyh2ohdiFwXXYA00lDrXaIgT9GFLiAVgWJhu1+CXzHoegAFQ6A7nK+Hhxj
WmPXhomKOtk1ZjJm4yl50mIQvGDnTdYyEpw2/OtTt79csT/9NU8RmIK3jcUKFfnh
UpbZSAcnrZWxOwUbpR6l/bf2FywxDnbRINZPCljxwDkQ/nHkmJU+SmCldpiucXh9
+wMC8USgZL6AJ0T4s9crhRJ/2SJzE4JOSAlJfOWxL8iW7ri/DUFbmPt/hYga29XN
mGNZ85MNfbrJWJTegsD49j9/CQqcj08QLw/O3DLJ6bD+RnvzRB9Bh2luKlMnFM8H
PLZJismItfecx5MzVwXfqOpKP+iyBXxuPVW1bUiPyFTaY2nwyem9NNIfJNjTNhB9
BobFD6sG1GdPhfIj2Lg/5pQxR9z+TK6n8CfUoAUlmYODU6bOjnrflA4s6THTB4+l
9/5D/95fIhemHH7gvfsj+cEbsIzY0ymmqDYHCgcq3irGoHju9YiT/MU2LhKGDiJe
8rIBVeQP5FNMKFcgadE9XJc0KpSSg32SZJCL5yq+1sv5IOGf2NUKlA/sNVp0D2kX
8wQHOfme0f0qTmNRvT3u/Ef5b31lxlnzMWsw66lewq/Nj64EjFSz5cU2t9+RSED5
SfnQDItNz1OmL2Zkxr+nszFZ7CPDj2NhkpZlLN8zN7nu4emWgo9RQQ7VOQ9ZlbDO
13DiHevIV+VcvMTB2p/Ys3Fq7ZNIimgSMF4rykEJdbInuDtmU8ergZgGgknxEFrq
iA47rdHzMBjKjWIR59mBZA+AmwyoostSfe+tSC/fgjSNy88DsJ7u9PIfyrCmAhBY
i+DaijdgDZVoNpoLJ/sxv3aQWkHM97cnHehFHsYbh7X8iWBzWmXKfo4AJShwZ3Ys
8PutNUzdxOJOy1Zwpa9EIgYC7Uv2kR1Oki5NgvG6HXyMZpDKFBEuD5CZQ5AoE87L
mI+wGONjcjgiAddZjU/ftrPmadA2qm/i6QBlNie5sa1DDroPnGA5BjRW9DQ3g7pv
FgX4oE4WSEIbVo1njPhZO1+52Pl/LkWHQSSb6+NyMw7ez0mMo88VPv6hwOA50KYE
ko1jaIqznQkr0zjwIC3DR66GXwR3mHHFVj28FGs1ovFZb0viR4nqTiprdbvi2toq
EPkMqt34xeGpCio1kUC6mj+1HTS1S6/OXiSam09QWjxcgzKTZpYm2d36tg0KuSAt
knFSrIdhcQ3dWq2m5vB7gZtqeTpH0zxZ7euPx7qsGVv7bPcxcr/ajNkgGAyyUD3/
C8yRnwfSC4C8VW1r8Kqr/DmKb6nbKubIxFVt/L/O1gIVd34fr/bzAnI6mE0oY36A
v8lJgbVmVq1dFGaM99WdJ3+QeBRCWJF04TsK/HNYtYJYVrgLCXQ1barb83+5T4qo
uy7GYFzVJxaaX/afjc7iE9XACSdcWwICV1ZypTP4FZVBkL8USEbr6NvSS3vBFxjV
KK+dQzspY3XIesU2Hdwntibn5cpLH/hXIu9QIPm0khN+hzte6jDXb3bjELZyy/y3
NiBCJSJZNWQerxfHh5yaNn93R04HPAVWU/2626j6tb8E4SMOrK4GMEDkAAhqkrhg
bQehbfXgbkuEEaudy567zJ/k6P2Nc+4VZkWzX0QEPA3eDwOhZdBVOi3/eXj8Tcbw
7QTW8DmNX49nvn5oi3zHWK6pPL6rsoCJEjeegZRhLKfBKtq/RvoN/NpjFhn8zIMD
BTqXK02bDuAczg0MLbJrEhfEzukteIJe0Tno/7lk47AnKBH1FCNjHjOn7a6gDSuG
eVDFdxZBPvqiFcURg7QvcvAw/GsF7QKNdMdL01+itQOSuK32sGYZv8tE4zl7xyWt
ujbaVzE63dXM26S8cvIQ7SaJYDwboO5JcHLebimM5aMjWyPAvuxjEhuoW41f2PRL
czH/UCZ1N2+cmZVdGYwIeik7wWIaRievJFRKfa+7gjvD/G1iBSionTwaawvd6P4L
rgvx2jEaPOHsEa1+WeKq5y75Zb4oeP6ZA/qcje9rMN19ZE7dpzDI0qmxmMrkaEeL
YYcg1RXQ+emlOBnAUWwRkch52xQG/6YuEnnVKgQf5P5/HkPa27mXHuUDBWsrN5uY
OfE3jIgudGC4zfe820BWUb0Yc4sQpInYIqWDlfB8JWHXafJF55ECYnxDDj9ixZ5r
szU4Ne80DTdtK/9VmrkKGhJcn8U+oknfUfaQzaDR/V7zrbY5SX2PnjGedRpCnP1G
B6mNOuAbLApPYQmTV2BBIuHm0HmzvTQnCpsANckqvTAezclCK3K+4lL/fiEi8FN2
iZ8sH4uLUEuyQAwKqx8ydTJghtDcrG9OkJMh1L58gaAUpUXG1d/csVKWWUa58YKj
6gUkiMaR16kQtvuyitwYG1KIK5iQUFceon27i5XyOLsRQ78jeqZB6P3090QpsgmY
RoliMxm86UGcxe7QOZ2m1qZcCBvPHaBNOO09L/X1Msh6zhjRuUqkrNkPAEgcnbhi
SVaj0vYvHAX6vCnS5z03P/Aoe7Ub/8UUkoQO8QJPZBFGFRuE7RkE1yntUbcQGFwH
e4IVKAuqAn+znUH8BdCf4Uv1rsqHZNWF+yWrfQhQzAVOTSlF9O0v8zQMSqCnXnVE
NhziobwY59d1bDPCp5dOTwFRVH77VQahfOv6XcTHOXYB8BviqHCZiTFGBHSj9Oyq
1CzAJyhUlzeeRe1OZsB64Y5XF0bO2XuB2vYiFAM/oT3AwaxhQx8llVM3RDddD5L3
3+y9aFzFEnTT9KgHlYjSsM2QQl3xoevzDLYGHijjhYv1YF1zUgpyfMxUbnV63aIV
7E7onFtuGdsPID5YWjxTN7hADXSrn1jImOtrkmvUj3Z6OWHD2ljX333KjksCRYBl
i74W4JN1xezsJaFnBqZwPC+TDRPc5AiJkIWmUWibyaa7CGyS8QYz9GKaO4/Irdrw
3AxxcPfgLF+tZ9ySQY57mWEgIEnCbhHklLxSYbHMSa6r2Fck1nM3EAdKpegMoOh+
160WS0tqmdW5Z6SwzVSND0bXVyNOPTzi+P0geeG0KdXAIi7QiNSgMRGJvw0Bjoum
bLKAwMXGHaSCxr66ja29n1MLcRBOVvnUeBSQt9c4Qv2JFy4Dsoykz13CNCnFkcDM
2I7ybTNFmQPMlsD7D0v4siTPMwPFtym052kB9bYutJpiXHMe7dTeqe59BubgN4V8
BZMlJRafyelERd5MQDvxqc7mXNbmI5QQURVHWqzegZnA330zWLhnbIwU8waCn42B
XGLyws1HreJdDk8MshTfoeIEX9y0ThIIqtqEWKob3AY3r02bRyinjiEjXzvTZmhQ
8DEjnI5IQbwf2oM+hmAeycMrfLMYXPn536cp4Oot8QUrK4l7UGNarjrzoLiNPPTh
QAi4GhiFgCZLCbOVqPzLjAJearpMTHFiY4dzUs1gdqXuaFG2VYAx+7CsHkZed7+r
CEeHEQtx7L0pjZpgMoPV1Kc+wn3Nd0+nlfts45Vy7c4VQniJKZHgBEawLKw1KhGz
4k5ZHz0QpMbIvFh+kW2eGQ+EnorejukXCrOdrO0w7pPZXI9D5NF2ksSKKbeuS0zf
3FbmM0q6hq3Cs7P4Oe2dUWRrmgi2ZoZSMPsLb4IukkwrbSbZong6mi7JM+4ufpSu
fa0TN/zaLrZv3Aelb66zfmYUQKuLu9OxZr4dR1qrWbIHTLSecz46txEwn9bzHp/W
01psq2c3HCcKfCk+80900z9kZTlKm49KTsTxAr9O6MbOltUnrg2AKOT/Q4q0qcWl
/bS7TkYC1rib2TL/xAVEZsIeqZQ9DyL7vQjINIVGwLku8FLByogetcQZJNaXXhK7
Zfo20lgYgluF86GnFxl8kHV6jzXgsZgGvh1SQhHWnvLVpCBl7fOT8OrZnLjR+Ery
73Artz5b1sEQ+mtu/XpArKi1dQL0V2YmB+bJ46i3HMf7M5V8flToDCQNj9QYsgdq
N1qgGXNPsTTkraBcWenA+rkY+NCAd+xI29M4yHjESWPJYB7WjqSQEQOySePUTR/j
na5m59M+6oNM5m4EChsIGrUfMKCpsS/iicdsfEsPw7y+1uyidAyJ3v2+heIdn7Mn
Lt5QpyUjUSFgdsDaVH1xTMR4+Gygk4ICMWG0vpHIDZvu858AqZFdq6pVvtxb6aDU
1pXBXmICfah7dJ2AmHLxAyMtP8Abp2/njGsjP6axUdsxytzqx3lEopKUW2D1lxp3
J9+5B45xbdTI4408QMCQnwhQCPA0/BkTnQq7p1p0idWX0grjAG5m6/PseGRwBVQV
zvQ+h2Yuy+4cIiTXx9q9H/nA1tP55k9ztejaA8OvLgU5yEYJq9u9cvy6Mt/sjjE6
mAPlvAVGhrDQMDVddvMDvRZoGNLhrymMlW47k7c1XGGneGX1S9NrW3Va8L5hIGtP
dnybQYz0yvHqNgJur6vAYjspjT3eigCyWvfc+9sEbX8/bRZzSlQVpm43vRnY57UE
Pg472WolhlvnGPVYbLsVQ7a6BnNunH/C1wJwZQkoOBbc8wHBL+EUA+Wj76F5O11M
AXsFbmOk3bjPyGkOh0Mja9Jyn0LVCnW2pPOZK+txhGNcgi7ZNw/c2vrUHOH1ltaS
fzkyKorulCERhH9vAd5pRLliqAalXwzbv+xDZFDxE3nkDWpx6mo7hMjwltzP9tu9
6lduyLCL6spIH/NWeiMSAx5DkqEXntxlBiXjIXTY6pJMYnPjjgTE4azWgXqooRt/
4u989NuA1338I8xtKtrO1gICTFByPE8foqwHUDj1sCAmjeA4XCPb5w62jr3xawCr
0YXjiA/IXEtafufXi+dplcP99eiN/UVucERwF1pJLiwcdwCQEiUkm/L5Ef8QMv0u
GoVMi/wyTqVs00XFtVAlcFyZxC5KWeFFtY+5gxBQZmB5jLl4qvoBtQUI2RPSias8
gw0safzO2EY87JzVxAqmpzMpdwekKvj/FZUxy3tYaz0B1zvckNVlMVwF95hNmGUv
slvo0Iu2RyZsqEWVg58fyp3k4xNCLVlYnnmAPTcSaBya1r1BSvcdNQyvTBt5R0Ru
mukYHKUxylA75aHcTOTh0ULV1b2EQ74pO9j49IK7B0SVglMth02QpqdznZygIoXx
sZtdVlDpHuRGUFYrX5UJIEWuvqLG0+PF85fTORBJlPkkEsbrCGKd1OryH0WVJjy+
bWND7PPiHZDnTdNRaPjG/ec4JQpRdMMCxABqD8QU1mVclodFBPcGlR65EK7bJ2f0
Puha6GF2q0pSA+jXFKQPFQvEAYWNcYforfxT4jUhYpdLbKch3uZgtlSQoh9AJ+76
uWNO7WrsIoGa9kHGr17t4YlxjSV27dRxDOM4+HdQpV0d/Ji4l61V+cy58GtVnp6v
5kwwvIRTT8EE3Bu1lVBish9P8k9XvxchHEwNzMac5OoywglD6ehge1divp8gtkV+
iSsC+G1+l6zCqWeroK3An4Ebk2HdJfsfsz1Ws5FsEg5iSIRGdPipf18kEcdx2e9N
tm5Fd28JlUM0NBO5m7E+EbWN7c3qqjYNsSzdvNII+9RrZC/vvOMKQv9M5dO7dAe/
t9XHNl+2d0a7gV0pSMHmYZzlO9tfXW6WCr5TuolbtDh8NbvWnD6zaJkXjd4q/g0B
KabiFR5GDrdvqUJUfuUoK+t/wUPSZk7dj2th3d/U4Gbzx/qZOS2LiLtfkdqzCdW3
x9agsogfiMlBNy9hRs+v0iI/J5tYGaBmtYpvkkmdSG9Pms4NSy6dh8bSY3PQoeO1
W3QLUdmHumE20B47t8O20am8XU4maNpGjn9JEqL8gEjjEGN2+QmPzxDozCaWDeeE
O2QRSi56uVWtMMhmYHQb+xMt2z8Fd5XwSYZvKo46sS9HluaIdHcnkWU5EinXRXjn
Cb+9yG9XlwQWsOyziFO+6p0oTbTLmtw5iN1re+ubLh4ib+Eu7HYPuL5n0vPJR748
rtv4ajTf9Ou6OIIiLGUbttc9r/oepgp5j683K83wsQKnW4HVdiqD18rEcgFh3UH2
4InUVozxhjB2rI+rRj2CrGpF4MukbjpCbVH2SMc6xnqLEtWiKkKDwBqe9zLipdpA
XAYLNlwBED/7pHS3tKSiKj2b4PbpcqJtmdnJBpUjO/zbsrNTJyMtGIWu1khT51kS
ugxE3Q/u05DetXBroe5YA7HwDU5fxOOs9c5GrAeykf349MvWsW5G/D012XcE2nXU
zK5tiHnF64ouxLRcQYA5j57T3BhhtaWbcGMOr9PV8hDcPqK/qJpk0HmwChS2fVTc
jbq/zFYhc2kWICXqCmynn2PTPtcoZ+o3ZOVBXEhS2PyUBylqAvlRmt/qj2/I5AlW
Ka1oZldA49XzF3vkMAyofE9lohfcG3gI1OyarWua7g6Ny6gqhN8SndRCCVTpCB5U
uuaQMDdiHhQHPLN7ban//VetNSDZBCDRVNRZFJfpXJEe1YhdZiFqBPQACSDuDu2l
XlSJEmX/DPzDIukj9i3bapc9ElckLxAYpGejxtZv+pV9zd/MZX/V9ZJJQJVLrgtr
aFgdg5ljd389uzX7DOEUf7NwKsPb0+cQ7tzgxDz3LYk/RRVVfFKR0Xi2gh7liH0F
88iXlAIK7ynhKSFth+eiD8ooYROPVD/MvJTCnnWOoNVIs84ngks7e3d62m/mlJCy
vtfgweRXCu0flrT0lmMoJwAjydfB0ex1jPNWlgrQx7mtbbYAlO9uUPbpItoTUIqa
g3v/6WIDNlpN6LNw/65imQGAYpjV7t9H2kmug6o0U3oKAodnH+hTeR52tJ7M1Whi
KGd91T7Y6ZvVjW6uAibOd3X9iHejP//ZXOGwvEIrRJgL9Bz/WXMU//lAHRBxtURE
N8XKZ2XV8ab13xirpqZJ8q1p8Hv3U+supMfbyMzQ7ufJy1lKdVlCAqpFdBJGVqy6
eAOLgGxxuhLrXVa8hfn4biPTlMWoH++4FjuBKLLetedCP1d20UEqgwpWJZjgaFPG
STAHaYMrH532PZ6Qe+7YyrC7wP2w0eB4egc3aCKbzqZJ9ZIoL1zQzyrBUavqcAVv
jWJFbL/K6Ap3oLAslYrNkSkuszltAFltV/Hf1gZmgniQWG/yrULquKT2BWfjKoNT
1TsVw37B0y1Qe6kM7ocpwaggpWsbPPWtqrfVnvO4Ie4mvSChygGL5N7guWC8lxw7
+jUIV1fNPRD6Mn9mNXoCzM7nPowWD11/AyFzjv7BDi6g0GbJYwwxgmb34Sg1lH4D
FwfCk+IgfWQcCvQ6ESpISfoNJqn0sLxxRLp+++dZLbeJVb1afEwPPvJiMfprbp0h
oj10bQ0TZArVFWdk7lEz8OS4OS73R+WkclSgb0qSRcLpTTwhONPXLfHFWIiZccNq
Nn360FwZbWIpQfo6NppZWml3D24IJFLK0aAe79oXyB/8pLVFgfE/r8+Aqfwe12CA
wyurY49LXliTpvCz3R0rAqHBmj+uVlwRbMZOT7bOrmQ0qhltUZlGssbLe00Hh0Bb
vpDlJS/0kbH1IssC0cWkXfYHh5C02bFeaHqojdA9cNiemiPIjrDrvD40YTte7OrU
YRM2nGY7alrjNjRIsQ2o6TvNgv4W4fFHBk8A66Ks5YfNGS6BV9Gy1o0zLk9lKPLS
pjVlvzERpiwpW3iwFWUxQpcOkzsTwHXFkaNT9netF0V1czf5ZCXVOyuu0ok+mcqg
hfheSEWSyHuq/WCwt7EDj2y1xHwfAfClAHI9mBzMzIxd+uZ4/VlbkasxWtb3+Wyx
biCh/wFG+1hTpM2A8H/lRHDaJGkUrERh7F3OKR8WxTf227WCS+/XQCkG0Bmz5t/f
if4ZpGWexWZB93ZoQ2Ay8KmbBccTkrK7XDay3bNMcMcIDUhux+fJ7MV3NmLhosxf
MRx9iBK7U8+X3AoCR3V1ipQaNJNaoMkbmQIcJGzCz5ez4M+aEBCdZgR0azF3/+WY
R7yioOxBFNjOFkK5oGMSejNkCcdwcCEzyuVqF7kjUe2zBxlOxIEzFy4zxDZRw/US
UaFwjsTUbUA9JOzM2lRu+BlEHW+FVOZc6XWVBE+77McX01CYvhKw9YZkOS212AhP
pkaQY8YwA/fdGZOY9e9oP/KV+zUxD1+q3TM26XrX222+ojiDpSBsL+ZXoxtLSlYT
47bqmb1vwRSTUAuI/nn7CS1zlnVvlJbOajdl0sDId7np/6aL3ed59IIK+M6JTf9i
Mpn1PCihDWr+v6y7yhshWP4fGerkUXkkj2ESRWrpndKoz3015+oI/JJWQQvWfE6J
tQW2t+CcFo3p7m1zyNhfs++SLXqNj+bKvdUCJzMwy0c7bS/jI9iqKN/u5+QaR13w
sKB1rVs+Fb1Q7mLuidYe2hyKbIpO4hWmQ1ZjJlxxjg25hd/gXTNsxGLdBZKGEHgF
8YINxMKK5r8IfB+G6UrlETwBwt6LfKm/he2DRD6uTRQjEqWJwXzhL6LUGEyywFq3
Z6DP1LWBfjhPoIpkM4lP3AaMP3o5Tnyomp61Bx1wWhF1LOPsPS8Qs7pEZSZWjwOP
uchhRD4s1yapLJ5TYZaRpgh11v5M4nyvwT9FbdenvjGBFwbompwsmGE4P6tR0/gx
h+PqCnzPSD1XbVkpPoZmWioOsUT2jqumwcBZhQBfXv6rjlwUg6dOR7As+l7vhont
17t35COPUxM5qld7v/fhzVz8ZBfDshQMVT6wZIPK6UwIuczS8gIWNR63TOXfTx3v
d3+QJHr1jw4OcvbJvO8yKziOTfs5dUK9JroTZC9EyVgw+rtTzRfs12M7wp63g+ea
kAb5csSZMGnhAY13IVz/ZrC5AbWrWJvS1cFK7QgyiDrmFDyQP4AX0QtAih65Kk1y
5U2Xq3F/VG0uBoVD8X0nJtOv24VPXxNCUQlyYEdW4ntTcDnZ2ruQtN05lswhJv4o
T1F9jVFViEFyfoHcn1yuwyOHShPDREp0O2CQDURM0YriknfgHAqzuJw+r5yXTXHy
4AS6y4kZ5GYIWAwk5GajUfr0c+s68bl6XX0TtfOyPwqniwmfisZZdxY4Sc58KrL7
d1XaurgPdPhISSZ/gu9Tm+BrOmHEw/nehH4OhoIT0l4egT/q8HBCuMkgm4+8m1ut
fODxO/bVOWg/XMgqHN8DAgZren+h5UcOJSWClRZ7GHGltufybBLi59KhZxZdolWf
D33/FS422ouVRbf6p5nMqYFxWlQlrBpai3PQMo6SD3cxR6YU/hlfhrv6L7zSlaQZ
IEL05uh7Hfs7nNi1tLHJiF14wiaID8yzk4C4yslaHTVqyHQhbR1IlLfdL1qAtiBJ
9CAwJ7P8whqfOOHcpIn/8PyKIQHd/Mlsh3QKvH+MMK6uGS0bAQM6y8UeJdZeQ2cf
jwmJsty1GlfDDrjsRz26ZdvuIjtZON8wqHb8ct1XwtwWFkjJ325LYbATsKKzseqB
y4Lb7fJrgKpPviigG6SmYpHi5qfD/QveywTzY7UQbLYQ+83AXMzzcN+zw1p/sY06
7UwtK5g0cyYsTIfDNVv9VI8MX8+YlhmupaRMQXhR+wJale8cZmz1Xkio8bWT0C+A
bIH3IQCdGQKT1R8LLX+pEqjRgdb/sHdSUBPsIEj48uDKimqJx9GVB8eBx5VxRme+
Uxj8bYnixbERTpkMFRhn0xdZ6RDyF6SvRA5XmRsf0R6pmsJnDQM3ItoIF4duUaqg
PKDavZsLtuJPP7FZSVoS9w2YtrYZuxTeyYo8jtNnN5p9bs/LKz5zhxn+bmu3hlN+
zKu4zhoXgx+li26mBKACy7LXW2NlwHdKB7tumapFEfNC7yebGrVCC2IfTmUfKL64
YfgNn4USjWu05DOoUWVhXy/EpEsJTiokZcnKDqI133xden3MzZqZAsrQxPMCeVhV
3fAVCJiEkrsSRXy5EXVsK9j8WVOs3SR+IcIeNohCsDU6LNCJrPt7ncMiPrEfHSJQ
mapVst11WoV6eycyxPiVLkOjwtpnf+pS+SL5tozXEhkYL20UDpmIWGo1iTHgBbx8
bOEzcZmZ400owtB7KhQg1pMCPfEGd7dOI9KbVFlaXyyGUj+woo2OcZ6UDVwCL7C+
301/vrD+uLc96qHdEf/t9pU6QYRwf6poPJ4NK653fwZXx5m5bRmkbl6vdE11uyyJ
l7ncuNONIIGa4BXWoPVBh8RamfZONjWh1sO9XRHfuY8vlcgVdqez2lrnMIrW5Ahy
zg7g+iYEoHsJMZWHjgBoFpJwNSdyvgvh8JZocVI0Ca/RkH5bESwvfVF5ID9236Sr
SFtfcpl/W4AYnA+mofCYjile46lnuTsYBaEalfZdFcdagcupBbWWl/yGbYRM3ZmV
NkqfBv1x9PvJA/KaUnw1ivq6sPcWWWZNMSdACriUhRtOVhWVrKBT/7DpUWwAXIZF
MAq8S/6VsnOW+AIN9DhSDEVn8DZCVx9AEvOLgH6ayKURQ3Zw4XEPNlSnJl6x2HA4
+mvtcAE5DPr8kSORPemLiTsmQBJDvGVkXQMvPtC6XKy8fk0k5uoSDR75p/Sv5C1f
Q/N0is/pcpozTwA61ftQQ3eB8RXvMrzNXfokouqgspjd5Ib2ZJxVWhXeKkVlyD+j
TWc3tV8ROfo4pVRXup+KrK5zJJONMA9sVr48UQ0lfZRph2e4jwN8YJxSKxkvwYaT
XW43WSNvCKmIXl4O0lQhHzChJoxjXhnX/7NV60a2RmdrSMyTmk292pmmVGEyrWgn
bLmucv3B3MvOoyShmIM9tgu+HOc7Fq4rtGodwkKCo6Ir9W6sS8Aa7tENgi91LFW+
epGQhYn4X3syFqkYROgRZHn39KzH77BfBuhGD/97Lg7UgTz6P0HUQ2cVoNvzeiGd
sX6sSPOslExTDm2+LPWPlyuRRt5d0YI2/e0dsBq/Ba9B03KvCecLlJbJvlStv7Br
6WHGAi6VW+e5MNb6GjvBPJouYmFhmd3pOue7sKH3HvGFfGYEvb3UoWdugfBiUnNm
q62XPN9p9qT/mbpYYYI7K9zCM5GguxqeCAIVGY7qd4LJFKKpkf8jUlJA03a1Onhv
FcG1ec0GEGn7c6a3NiTWeKSA9RlKwcCVyUYxUBoAION0eMieD5a0TMIIn6TbPrFD
ZrwjviIbM4md9NwvqjYp7nq6lOgm95+UxsM50wOer2gVDa5R0Jkcdjmdg7TxNDsW
DN0t9g8o8bQxj8TJXQnTsjDkmk6IUjGDajUhnU+alGdGPysdVOewNqSYJocGOhCt
mUHqUGc0mO7ox1j7qQHPuNKLfqMOBxrNp5pkOdX85udfodngwGm5ZZPlIxxNoH7f
cgTfckOFZbeWngOAjsapycjMX+RRIgy2ID5rK0wjkK1eQfuQB9MY89G2oqfCBsuX
ZJoE5OU0ZB4jJqABxF8bh+Y0ENs4jUGW4G9u1uixz6dmDXsAnulu5s1OcZxXb9yM
c1WwH0CsfzmhdWcrTIyEz/nBViK6dYX60jOfPFwe5JKyN5QU4LUAXplK1iJHskvQ
ZZod6BbI/2Tw8IhfVf3+U6hzBgLEgKpOliotveBfeBmZHmWRiGZa21bIvQFSAHad
K9394I2RguMO5K6TQp52Co5eswwpEAO3PRP9iPAVWtftbDmXm/7wGgiKcbez5Y8E
UsCcFLykSBYroEV0su2NEo8evCDYFvpR0coQE2REczgi1kVUAl5zfSeaHco2fh+z
r4UIlIn/PGiOryIpBFw+RKLsvKe3XkfxQFZ3qazJU1P4W105CVZNYLgXCVN0NJMd
PA4xAzu6b6kFeUJnX8N7xZVUMY/KPZt7PA31k4IyB1GPFXA1JGJvKvMAlMA24t0s
1suQegQ3+KkASEpEIQ7dwS5ngCiaTrD7Qd1j/DFq8H1lNI3FWuyMz0OY9YhBSq6e
JdTDf3b3CLLxKtFAd9cq9XhqlCMW5vq/brZJmZlJes+/2ZS2l4pLof0aCUhJ2Iba
mcAgj6V7IojZYC0kvCRtNLH7EtYog/h1xzGNQZwleFjCCBAl7EKMwbZ7tFNL+zMi
FWWvrNQdz55jl3oRkTOq2L3hJAf6ehPK4fS4dXP17QxwPbHV6o5zsjg1iGdEPd5w
5AEkw2PH9FinXB7vVubTKqQCen0i7+F/y+73wddIIaR6iGd8Q41a5EIkUU3M5fxq
mXpmnJWnSTHzsjgPwypO8k2M01DGmCiUOqdfKQgOEnDAA7sfukqlmBSd0USV7C0x
2dcnmFxTmQFZqcFmgFJIIQwem7M7gAGTA3JKSMeLTmXwAnPN82gHXlbqbizdcjfx
QOZ+bUqMHDb+14zO3CgT3Yk3m+TG9vugfpibLxFwSWgHt0hmQNCkaxVCuvBoTsdb
ZVfIirF/XftPxR3AuyYHWsepWruEzBS7gWPCLQ33GYv9q2K81iHXqZ/8IqMQCkbg
xEmgfesJRoISuaVQ824E5/0kM8DrdFMlJ6PyJu8aIs1pLy1DvdNpzuK1HbMYljPB
EFLdXqhnVARcw007aNBz27c+GPZVsBdN0FLSPNTB70vAKVgIslDN5DPdJmupg1Az
WvpXsA78jNvYOxx8OvUkIhDOKL6RACbIORtVxF42X2zGMtgmg0WUoqLM3l9fIaln
ntmtCUX6vNqs2p9KKmVSe+z+np7nALVdlsKTRdlE5Z+MuohWWZTx2V7WcL2U6bFm
wwBAz5ToIzOCGixbH9cYoDSvjw6ZCHpIW2ztX+PAKMb46gNLdtcJ/fhFt1vcKee6
gzKgSL7yVj+GtX1rQV0McGwUvZQts9uen9V0UubMdDqykwxRoFOHN/nnfFKDWg1S
reaxNRd2Atv50JKibMgofrs8a1C135erExTpTY0Jvl2XKo/4LbHWCYb0b3dvNFC6
izaEG8iZiYIVCZpp8DLvQ0UtMW+JFRNmHcrcH7AL6mbxkasHB8p/jLD/X0qAxROJ
mhFM/3XuQJP6pdrS6CPFy6AWeWzjL1xq/M6RE+gLXPPW3Wa2kTckdiRoC6/ziWeL
ESuon78Y/tue8jZi5Ik1DqFnSJ57d+LPB6rBAHemyZXB5n6zellLlcHOiZIZGL6N
ul/IGwVhyPS8656Lk+rL4S/GnUHRhHWLo1o4LOvH/SpJH21UXToYQ2BHudKuPUwx
3lCkbWA5cKQq8EI7MX1e7ikhIyNi/bWAslb0zLfUVTp+9VMPfRiMpzqOS3mqtrs4
mBzF4IpxcwuT+IsNqDY4sZv9Fd3CWAjyqiMkaVzfnGP9tuha9oEw3ivwzUg9nZKa
h9uFyCaz+iZ88eF9j3Mak0EKdVQVg6IMnAZi30v3nDMTCSlCo8/lv8Z3RXbrKgCE
aXKg71jWf5iaFC/7jaWR7saIJPunI9B6jA0zarDZ1zOEJT7HKBH1hmo60aUvGA/n
5Tskm6Nn5AU8Bmk+jg4NbagepBctqpFFOR/Ftkv0exJUX1CSTlIck1FjzP2EkTsp
YcnK5F8ZBkjpKzUbeSAYDlPxBc7kf5d91XAgsd1D+waRGOH2hBDU8STxuxrEqSN+
4qGc7La0IjSOFP0N/t3EDXCVAno3iIqv+cyvkHSxklbfn8JbNabjVz6DTyiNX3tg
ekx9EEklcAWv8qILeoqf2ethJ7wenhmf0AWfc3Hz64nqHOs13qrjiAGjFdAlKUzq
CkNgQFKvSeI51anO1wyjPfGz2wkUx9LTLntTUCkxPX9BfRaevQ6b7IhRMb2fY1KH
MS0tlOgb8wsVEJzrlLqYL67GGBJx8MdDwtIJgZkzcefCRdwJG08nCkyA+bGzBcY5
VM/2mtgBiKG2CqcryvtCTS3+QaQlBuZtREExXZJWDgErtGk/vlnSOY61hSiRKUYK
scq8yWlUZrsD9z3UZS2M4SvyTGW5D6dGcqp3zeJFhLOWVTXuvnChSBWnD9N2SiAS
Nn0Pz96rAfbLLpZq49wnFcaXmjGJKvDBAu7NH/JMeXcRltVFjC68ha8ro6BX5XcK
AnIQYkizWcgUpJZHD45XRvhUnGOXFhuq4/CVZPsjAu2miD+VoMKkXUl7UyLkcv9l
gQeCad7jjy7kFiG2Cg0UEdSMp/1Re4z+MnB0Rd8IREHBm/a0txkCyYwhIkycNpLP
jqmCDXj6vEurf3mg/pariXyv1cRtSA1jvLGJK9KWfwhrdZPpQEbAjYo0xaNG+1su
4NZIlk8gvsOrLkb21Itjxme8EPjLIpxURHB8O1QPwN3zhsARgqVHJwGWeubQ1sp2
ZXYH+my5ysin0BJDvVkzCgRkv7JMPbwKx1PsRfQwxQ2hTOvAkwN+JusDtSzmkQW9
Hy3YqIiRHX/VV+uDeLWdIvRt6ipTTIm8IXTdDith0tkw7O2Cx/Db4k52J4EzLFMC
hQZmKn9ME6rF0akedcjAdXtsk4hOx7vYtOGc4UlvH+ObzmWjcNVE/Xm9R2PTVbGV
uTNtWu0Fu36bXIdMV0FrxeGgsh9MrlV1g94yfeiFaOAB72AXD8jY9OT0a4ZUZi2b
0RC7QBuCdaFF7y9d9udyQ4Xx+7RkGr60d0/7g4NjGFZyfAm825e811WZrLHCKY9T
ydXIoZpco02zr1R1PiT0bNgSwVqWvgYvfrt/iFECi3jWEdt0a/wPMEYmB6zKn9Xr
f1WFF65pO1wlDJFiKeeeEGsARLcGoLrnv/n3tSB/jyv/kEG/w5rtEzRUuGbjE6xF
DZ9UzkzSxHwsLTH5F9fct1SxjQANe6EXAZ46dDPXadVBuRYWxDLihT70Ux8cM4D9
cLWSyYploMPp/w3VgPwr0lkHfVbTOiptFXF83RpkZjK7V+hKBO4IzoL9QFLahTNS
Dm8nZllr9E7HEEBRyu9zcsf0BlJaO0PmusuR94rI6lQdabI7Be5CMXOqatsZPaCd
kEpa96LQ8BbaLe0XIfhOk7BRh9CiR9rqPD2oNUm8VA3BMW4DMghyglk9BWpOfO+M
gV4nnXhm++7xKqCsN/Havgvc4KpKqd6GhdqXT2HavATTnffcQfOAXVOQCD1HKznO
Y9wlHHIR/fahU1pHcZZBOFAG4Awyh50xdKivaTPHUT8qYV3E85NvxOgh9QM4EuFl
tdwLrN3f2aq9iyDbURKDPB3zZP2yMTd/fPnAc0w+1EFe4VKiB/CHeDw8DUdoCWxP
sbamNo3v5egFW2WANadjHYdu6yklaS+uoumDBKaUCSocTBbKSzvB2u9fFTcScQgO
pwt6TAbeA2Ak2rC3ns0cYEz419pm+LQfTKJdHQ2L8XK2qdons80mSmJ9eITcJFjg
MEmiCzYt7rwm3ka3OgGUMXA47EF5MZSR0KkyYfdIa0WeVQTwZ4Qmbbvf+BnKIDNx
/ye/ISZW+VnhsChfksQdgkLM071/HohPhRs+oN8JhyZOvabdNtrD/nDfPWukLuYi
UzxZ4RFGec1KTRPws+poqO4ss/cMGK3McZeHf7/KD/ErieOt4GBzW1vkn/gDAg4B
LgWuXR7lPG0B7bsBU2/ieJxNo0wphg8oi2/DpN9AiMF+Ja5XsXTp6Illa+sd8EfS
GfJLMYy8LV88B13/PodVZYNRlROgwDFIl5DnatGS+VGfNmTjkGj7uzdOTZZ+TvUV
ExfPxGwz49sNcv3tdGp5VpFsdAomqNKqmqiFYK5zpJfEw8WmAFZfWuu5Oy8hewzq
y++P9YidKCI037mFQ8BhxfSNj6Q11x9ueZJPsuIbbxVksA0uGh1RvpBDS3UQ2E3b
N+0TYupobmVSuH2Tp0H7gisaf+MhdhhEKtQjq4aslLXTbMmjGMob54LBvTvo1bVG
hRYMeXUVncWk2ZzPaaStgXjaDkKlSglLSGrpHvkV+1EkMIy6hP77WgWggc3NWSWL
kuZ/W3vTPAI+J3Muxc2/fTMNIbFZMUSHPJN7Lt57M/qNbW0HkSg3/172owsAifPf
bBxtitV4U1xFGIGZWy8wFAE231rlId6NPmDZ59WUInu2i2DvK4tdoYchkl8nIBGC
Wz/mcYux9WbweHRGYLqD+RfIXoQl4kiu+1c9qmznr/MVZzqZ5bLt/tSZNTOgRn5U
ulh1tlDiOifIzJ6D1CeBqJutlYVGlKOzxnaP/NDuFup23oIQhYRpOzleFDjkfbZM
EMU5C6GO0nTtSdJw38quXtpwSoNpnUiy1K91IEs9v2/DJMFBFwqY6UQRa/nZ6JZ6
UwzxCmbA47GFDhYWfwnW+JoMHiul5rllm6Tw8gnIklF8Yn/LD8aIHJmtj4vj4fB5
r8koxb31KwbHdq8mzOBZzs96/Y8k88Be3o+MHV6XjZ9JSBy1W2aLm1GE+himJ2n8
NJU4MXavDhORKeQK5dEzFmLOOlJ6dH60zWpWpCIwltfmIWaFEfbBjPNvTP5LUyC7
drbcGOSD1Ug2AZeCkaOGP5VHYNUExgDuXkXILXkzOeVrvNGIhlNedaM+Z+OWzd4J
BSONkJUadBRmcRRTB24EDHJO5h5mlKPxClcUa23MgMe5V3oZkROFbn6cybzySRct
sfJ6ikFxYcDBog4wlSfuJNao+Jn6XnsrAqKo0pEH+A+L0pyWIYUNRdq1h5p672Ed
2RQMWmh9kWZb4Jc6wu/RJgdJ4H0IzRDKRfJ4ypnfMTwECFnV3H0WLn8Y6tsV0Ll5
ZkINanK8LR/sZLT8ZvTijdgktjMywmWeO/IaCY6oyw4bz3FZ8NBEuM2XAX/jA3st
JDwXP0B8ZUsuZG/c9yivPGn7iNucmLur33n/sb0YCF34RnkR1nUpBZpGyUOAEu9f
DeQ5A2qbNhvQNyPzDuc+Z5RaShnPhXgk7SJTNGZja5ubt5bywgx07JZIql+m+F48
yJ+RlAp0HA0a0JeVFqYTm/GtvqjQosqUe2fWnc7Ux0BzKD7E3IvG2V03u8GZ78gV
AVuihL8G+x5/t2ni8R6DRAJiYRfxkb4lJw5MfZxd9VBbcQGtoRzFFzDdm2h/pNAm
3a+yf5Oh+KuM/jx6nQchqsiYDJEGtwhyS76Vi7XRBmYR4FQcWboSLdAaXun/M8a1
+Eo5XcgygbVCDkJDN7GyNTDg282/n9pqwixwNFmdDEFCyBQXtPb7uWjGE/rKsZuy
z/Qnnf8fjJYWo6HpM2mPQK6OZmF7oxDo7unbYTS/wkJZ702DaNrNri3uMjIcaZC9
8075IhOpwSPDAMIZzB4dplZUagc5fZJcZHB3BEhNAOoyhkF7qs2BtEFc/ANiwPcd
74BU96F3TFdFvCpKGgBL6QPsuVgpj+ybGyGhVp5xQVhR4GHkcmTi5AjhPrCb6UA9
wkaZlPHFtpmH/BcMs4oK+oMXQEEM5D4hqPRUDYwZZXkfKORnwPJ/DUoxkmCjzT+W
iWdaOmxkA/MYrz8Ok4QBXYKyX17HBB1N1fEE5vz0Fcudwk/kUbNscJTRgMafVY4G
BAHeL/OpWZxd1LCsU5RcefMpBz00F39blpChsYFp7AJBndEejpdg3bZRQD3EkMjx
62iFf7nyZGYdvu9IdfcyfQaHYYUltXIcJx4e67z0seaIjOvjc+WbgoqZktNyUs3W
O2sUuzLBihbnw1XKkHRSW8Cf41mHlluyEV5QhyYOItz02HuhwabRlhuxVMSy13D7
M3qSfmjvXvPM5RD1bT5G3o5kgLSdq1WcZbtJUl17FNksDeveevyE6vidLknLYWZc
RPsYVI+KP8IJ0g94GPGQXkcWIw7V78A7PMCFfKYkknCm5BDLuJ0zWznMI2OPXJgC
RHHEqiUGFNWSvaedmVPVJTUxrCclbk1347nOw7cZ1Mry4rivxtIHWrwQMPn+qquI
uyQ7G1LNmloPhDAyOXBOE1vRPWiei9qmPnOV1Plk06FsFFqH6rY6k3hGk3phruOC
MhbZjUPksT71LFKHZGBJZHZ77Jyqkk4u7wFaKGQZj8OtQxcVKf1auc/py8Z+L0PL
Vh/5aosuli0EyTKKmlI1HD7yEAAoFwWLEcGQXGN3Vj7uDA6BpO77cqv63R8PrX4i
LDEfL2NCxoVumxA78rqaeby/O7sOk27ATprBCNoLVdVYIPmTcgYWlcaxm2g1pTdb
15OEiVVOxsmJygR4u83hP98H5vMBU5atsD8j1GG/q0Kd9ONGamxyMe0nKRSaW68Y
Ac2jBEnftp5bFn2TiJ4+mHm7uUXchnhYjs731PiqusMGAGQmPwgxFDu2nGVEvxiA
DERqLSSfnM77xPCMHghSITQMEM6D0vxygrTGoffbsCm6x+Ay0c3uHEBvq87RQOch
9GqkLBa3RAQurtHVlq/+H23tWG2TzuT1FAnMcGClmfeYGO4DPaOy+teXy3Fz7cPa
RYD4KybCNgCI8xR3xY5zTAm9XmWlQaST0vioppMW7LSeuzpnnaNM8zIgt3IjFsk4
UjoBcyjVRbn88JS/UHXIGEheAA3qBtxmGh251ajEtY3swMpLvtNRP4g7b8hjOyJw
Zt1Z5rMlD190tB9qe+YjXn4U/IVChJAGWwEPTYBiXhoG8z1pziZNndYnN8IXgBW2
nkW0mTTPNxC/mzdgbP2mkZKUnCEAwMFyNIVerNQR+GfhKylZm+e+AxkziAcactZg
raOkgrQzzN0FjDa0DpRdvKD0P1Kw+Drut8iBh0XsnGdYSfpD2kEGbLj/rIXnh3/E
LZRonrOWQU0dtAQLrqcm3pZ0u3vgtc1aOPY76bDdmXibMZaDhtjrxFYabt61JqIH
bKHEePVd7Ref9bG6F6AzXLM+L10PegO2mGDw9IG/1ngDjeOkZmIWYq61eMpQ/VjZ
cSkouo4HLrA5I9ml3omEGiHQShtCtPm97DHA2OXMXkaPCDGHZEXsXot9PRkpqHJZ
8RCe4LZkUU5Ay57KSFM1SOcJq+itArlQl0uKyfRAYl2NQFX25mV8y87tA9yDBPd+
fPPwd3eqnEh4mJZCyQ+mx7RK58ehFeIjOKg+Yb6jgoE89tCYgXDaE1wmUoEIgImt
alxSRjXW2xG6+YhukSLPuSKhx65g3vLPKoJHNDQ7h2fqkxum6TSvfczNluc58FaK
MkqOm2uk5680W5iXfnsX/kNEb8yqaE8dQp6cdltxU2eub08MfNqDzFYwpNnzvRTe
J4+4Ovivx1Un41WRWRQpLp/E91EvRPffZGusl5J9AQ2DEcDEVUpCa07b99p9kot8
H8g08yT7+q3L/DWaQB+blSJoq33jA3mZrCnvLCGdwJy/IawKZPFFOADoJ3Hfw/JE
nUQQJYurvEIZqJAGtUx/eSGIXQGOFRlaaZuMJVZzfgI02ZFZvprGK6b3lTaelnEo
uaSnTrJY4yd83TFI0We71EndwPYPXzDCgCzgHQAiaSJNt89kFuEFy4Ylwm6eh1al
TgoP0NlrUUs7fmStGKYYzneyiB6ow6HkcR9E6dqAgcNqcq1605XA4TZ4V78SG3Zi
lWyOptwBY9+beOXcFPKLGhgEE65QT0twtj33nBtF710dLS8M4VzE5BA4ENvJphB4
UYFHYApZ1o+czt93O+pt+KTC3A2aPVrgPf8T/dD6OEyFmI53sE5CZnEHPz5NUZXI
dBIwth9CdvK6lqk2b0h/fE9HH4AYfEGG+xppyC9+X9k3gdcCp9ffVZ1H1Oinswut
Aa/wEjHAA+eYYAUbi9d1ExN41b01WuIg8P6CT9bJAhMy1LUFfFW9xE1Eo9zSqpd5
8lnoYZll8yXcjwypJIGaeerP/aQkcPNr1r/lmrK1sfUggJDgeKZUW0m5DnEkBA92
+PAuDB8qa+hyM0FHKXNt7uQt6GtuMNqMHzR8bLdK4mmvffCXafxxGwtajszeJjmf
dTDSialVAfxcViQn8oyHVLwfQuy8NYzySrhbZTM0oXbSX0RSGBfie+oLLx+nGadI
Zx1W9DyiT3UBUCdM4sszhYqXQi+uKjbgtrHlPCerhxg9ex9Xs3jrHXd/o+AJikRj
un2tTsHXlMjARzWjN4uDvKxiToE6z1xUcdng5wsh/d81AajDKvIk5bFTt7Ax/Dgs
N15q+DhVRJAzX+fbGG9HFlQ9ap24o3+t0FByyBiajksXc50ZqmCvuaGnuPqvX0uo
ZcmQ/mGkcco6MJn4MLkSF8WkfC9TDy9iZr5vnekyw3Pm9LChzKtQ62+re6v7wtfh
TCG7+Y8gGsRTLqdV/swlprXo+zdiR+jFPKXk0KPn7nv9Cv+RZtMGATRG593/1Uam
VLYDlqmzoQJAzbAmzYoNwTKBcOatR7dvDPf9EXgcTqXdsLrGEZXm4+ohW9h/HZFy
QY4eDksQccWeJoi6vQ/HUV847xPXr7zuS9+v7vgtzzwIM7njasltnyfsQiHYfvOu
gIO5Bb7pjQL+L/F07sr/tqTFZt9GXrWZsJjLABGYXYyYbSlq2pkfsBPYp3T39vDc
nBx/PzkmIln6EuYkID/Du1yHXAXG1HI9KWZ291VR6XGplQ8aTrNLee/JZbWrODqF
s31XM3m6ONOQ0aWgmKVuhvDbSEtsZHP1l5o3pLV3ZD1N2oNRsDLYaR5KFycGenAO
Q8MTObm+HiGcruTKpUmnf7NsmreI0/RlcEdZ6t5OOv9/l60XLlgbzkzEvDcd23JN
C2hw3ccM5LZimIodFuVTxnjE3lF5oX0KrQlD7WXnZGYwZIe2q4TLiJ79xBp/HlhN
rQFp+zsAQocRq4q9J/rkyk0U9OUBh6fd2NOedhdxdMZBNKi8QJq2A/6gIiyBt1ms
6mdZlHtBRuLohalXDCZzRApzv+uMpd1cAI+lVqTeVzng/neTKxWLesCDhQSc8pTo
zyqiw64qvErSagU39jvGJO1dflAp+2hGjXDx/NfCaFgHywlKBOuAKNl2qBtsJRt2
CJnFAQi4xemKmXIIsTGXE/IaUVl/Edg0E9dku9PNNSn23WFXXIIRSfGr0tjsGSlY
ZGUHVqA7V4RH31mkiJArrMDn+37FKRnfq/xgL60M/+6b0dGDGAeGEg1DW8QMEWIa
A3uW7829JVLDKL3fkOTKRM/RHaY8dpUzL8v6a8Oe1brJmetdjvVXoURXpBNakOc2
44FxTK9k4Nl1pqJG0QDQC5gwf2RLhzYCwlAXabsq0amMKoalE/XPf/uMoGoyZyUk
k09L1i0o15cyKPnvA/Wd4NrLQLFJn9UyMkscvXBV1P7UUnTK/ndS5TR5RxPLMN7P
CdVKYhcyqgvreigmXsvfpdQWKufOzQ3t14psSuaroOuLVZew0bacCZ7UukK5PjDe
V8Kqeox8lK3TVntunsJXS6SLRPp88W67mif9hk26z7+d2sDZS0ZOPpwyThv2ysdk
cZp73fahI4SlyvQoeY8au5PSptCZT5oJgKkZUxPyiDxtUroHskrgyZbnBQedALtj
BZBM0Py1dFlbpOK3crxsMY1j6hmuj3/V7Bkioj7jCtiiUHlxmWzYANTZqbyKw8TI
NVC6pilgphi3VwezAjgVg1F7b7sto28hrsudSNLxaGNUlIv7HA947VzVrlteoQhl
16NJMhJUeU+C3zlXDP2W/RWc4hTNrClR8zjQ3V9f05PQfBZ9C0l2cjCubzkkIiXl
Ttit49J10BLE6ABlHqLfc4hpoO4HFUnXP1SreB3r6Lpvq4vxOrBUbLyvsVO2vDwW
PGM/K08OT+L8mty0Jv43rNr99Pz3T0FgHZvm4UdnI6nVlFJlDK06PHl+1ZtXh+kC
xWVQlDf8wArIrbNhJlFXj5t+t5Aw4E16B/Y2Eq5lgpZiEjzUVTVhHsrL3GJLhAyH
U/i2OWUdVCOrC/+DU591joPQJ8iRcBfjDYE/Lqig4GQeLJqjK/5q6Q9OkXyA6rBK
psiN9xCLGyCNWWyu0jCkO60UZT9iZydlaImKF8aBvLUAEjr5gCSxlAZSrGt4eUYh
gaMi9tZ+HlZpD9whPkJnQVvStbC9Pm/4ZFubGV1W7EoxSVCxNBEOl4nJx3aiHY7n
NHGg1rCIsPEpmnK/kQdxW9SdIVi4TkgO6UYNoAKu0o6epp+HICv/aTI6NFFPLz93
I1OxlVyQ0XsuyoMV7ToKLAAje7tokWnCm/rSpvV8kBi0VS5pSQv+a7b8xg/oADg6
RjyJIAjZQ1be+zAGLGyf7NHOhc4jsYyi3WS42Ue6qyh4J7vaq+/Dk2iZy3F83JH6
5GBeOf/MJk58JqFL8RQ4JQIjYm5JbpWtxIIMAN8+PB7wup1I4GLTCV3P2Kn4pRaX
cCt/Ez9/jKF6E1Tu+35XkiaVAIWyNPO37pScmT3mj9bSBGs80I8ZJ/YK+b/KmQBA
YXB/o1Fo7YWZYxq9gV6+d8pZySM3JfqRk4tGreVmofuNK/MLDj5Vv+JgGy252y1D
MJWRa1CBJdc120B2klQHHjNY/ZRqkj8Gd+vZ0y8SpI5V95bo5ixJFq/8Z61go3cy
CabVGA1b02dTDnUQO5bd5int3Kwma66UHctnkeDmDFmPljStF8Z402Il2kD+ptNX
SitgK7dmlzSZKCCVngy3JueQeTgWIWWM/zTdLTMxaLH22+/vfqqjJ+2nuobmjo8G
dzhVvy50dsnxI5Oh9zrfFp+9VXdFYodOIusZTb15WBYcsS1+4o1VDgY40y+CzUYD
4NBCShGpC+WniWWfuL2DLgEl+dkDhRY/KGrMtUt7D1djXxzm6zRCgwLw7NztyZaT
YkSG30y8h4v9+FzCLDVG1xabhaJh1e1Py3iCVt/rXCAgzi1hRDlZ7U3mKDHVdh7I
7yHW/SgKJz96/mfkBJ93U6++tPiM/Y2JOJx1dkgbee0PQ1rEmJUAOLqeON0Z7Buf
iQMKRQffwMMQx0JP6vpoAtUf8/rDv/MF8pQOcAH1pNPqEdtjz31PHDL4kmmD+4xb
HYnkbPs3l8DI0aF8WTics3G8/0e0wSAi5skiSRa1GHxcH/gwXBEPG66zaK2R3zl8
F7VDcXtj6S1e9OJkSsbyWXmcVAF3dVbZJ0iXf1SW0Uw38IePukkXy8cL3oy11J28
bDMtmyV3j97relQ72wGCqTqhW8gCc9D/gq4cQodK6tP5+lpr8MtIzHS2aYvJxk3/
yCmU8koFiZvNBl6k5py93Gl+4gAtn+dLCRRYoClDGFEPk9e4mqQyCcAmmxp+x49Y
rM8/m3Xxm7fLWAUFC2skZnS4spT1jgBrtA4/4aQBJpPdsHZwD3vD27LTuVLNDDR6
hA7V1P5QEv5vOzqePuYagt76lIPr8BQejxladR43xLkiS2k+UC5Q3sFpZEY6rzCG
7yS4HCOL3F++LLrH1UHpkvHgRkQmPunA1/ecftSiFnzjtzeiG8NLmCezrX15IzuX
d6DDTYgefvlRKvcniEjuSKfXMXSKQCUw6zrC37rCFMGdSr32T06eah6PTEu/ivN/
K5cJgopW6xF3JRp96DaGe15rk+ODYlmZjR8mHqIjhg5We8VpWTqujWm2U77Cq9eM
RMnD31PVOgBkVZ+v3Kx9IOLxXfzwgy10nAxLd1Jz+4nkCqlVTX6+mY8jwuVTf3DT
abnD7WmCPp2SnABDXxjjGdX5KTTOTzOGpzdd5X+tcImvMnzbuJdEIEWFoLJrpwzL
ywWFMoHk+ChU57t7gkSb2w+3iJUoLcLfm9J7jonVBEQKvrShP8ciOxsG/qE6SzHV
T2Pk7VDcYToiwfR14qtLkqDrPqnZJtdvdqOWy02HUcbRFp4b0FgTyrQBnUGht4kR
bK9dOAZdE7gEHQR45/xbeFMOm0pcrqCPCnwH+9ZGUNFWiV1MvrkuQcINgTqYpYP+
Ya/O4MlDPFaFXktX7t3eMMVXstST8Q3GT9GFd0iUpkEdLrSDf/7afPHWNdKJitIJ
DQezBEtAQBZ+jgZHDmBu2SbaSnl3pDkt8oha85szINDkEW8IOyO0a5+BVnCk3+DW
oCpWlg0qKSS3ATYo2+ehwvJxm2B4qpkl4tg6XJ7THpLAsAjL7DVZCWLWh+MHF5/Y
15clKTuUHFkHSNwtW78ustLLZkHrAqDED0DBCtC1HXQ2g4N60lH+1ZbEIXT7jSYX
p9qdnpbPHEHJhE/lC3cnBF5vr56u437nt3wzsO4l55YyWLMbE1lggCLFbeqRFALL
e//nA2uhYu45iJdJ+0lUtc5qcDejqT+yDek1RRtcP8YVr8yFMzl22RF7QSvy3VbE
5Bkf1Z4rsQlGByIYCKdWOs9XNw7lPFe2Zj32sKvhi1q1Gsfvt/H3Md/F9zaOQSgz
aWXuZ/UdqBfqF6SbFqs57JweOTbcAhW+c2/6LjH5g2Wzi3dnm09OV9OWJBPz2uch
03n+mB/ZOddHjFCV/dXYnZ1aKAsBaAWFq8O0eMooWARQ8iLM0VulRGfPEw+IxXqE
XEv3uRgzFpvts+tLos93xhGScYuA+gL0nW8iBsaDJUppX2NlWjJ/euCzBPa9TCZh
ztzGZiNlg2Djb72cF7Fzm9ia0wf4y6P7H4ioBQ3Edw2+aWI4JHTEu0PGL59J528L
+6zqrkwJyOdHOGRtZwt5EkGYdSB09i7zz8FNsZHMVrdgc5C38juFhzlzGY+EbW3u
vuzwzmelMizaBHjB+16hr2eIcPkaxxYzYFtuzYeRf5hjOziuTkoNKnaCpLmjlp5e
3veLnQrnmNOz7maK8aUOuYCTt5tva7zWTwTAsKk6nqAS0+kkz8oZLnV4WBn5sXUJ
MmdgRqKI72+YRcK2MueD0D2alyZCx/PsVrmy5rQaEnj/xWQEtG5UwTongIbnnu2K
FeWe6SFsFnonzwJsOd8lZd07jj9wLKY/ZBdwanigXA1DpOatNB1VZI4oY1jXmMPS
zKQ8jNT1wbEWxrROYfxqt7eAbDPCkYzT0a79Rt21DM/oDFclHMNGqMsZwSVyhcm+
QS4Qfz6Grr9aEo4E/fWHr7vNufd/sSQ69YzWSawofGIRY49VmhU/A/n5+OiKi3zX
CEmZOnfP3UehceR+MLdt5/rMPXSDKJBoBbgVP8fVZu0MNbRswJxzyyFnY5xIVbVk
jqRKs2j2WgNjsjdCUrxLQo0sJPItu8LOQBku0076NM4/5X2qzpmeoktOmdb0S7FD
9CC3+hvS1VqwRzY1OnLkIRGzjJWTFG6vg8AUncKJvRYLlgCIN5sdCtxZNxUJIT0I
2fQVh870KY0c92TLGoDPfK7d7dxzpuoH+SuLb2c9atrYfdBrbQxZJZx2R6ibaDGJ
3DwLOd+b9PD0iVfOFB9WyP2SBghoS39idGsiUqmx3/eT8BPTPhyj4tm/NzmgU2T2
8/d8XK15qgIf3OP1ZoHt8QQnzqRL7ZuPCNUkNhxYj7gC7jmKsI/0ng8jm6RiUBFb
3eKIGtTdTaPTZpppxiooiZnwWD/Wo+YRSKjDgBDJoM9cY+H7+6lMBHmUugkEEFnv
ZfmEer5i670YveYEybzWHlB0iWWnhQnUP04ykHCNlZWoNo02RCjoZpaAPvD5hxfw
7FdMA3daN2a3CwCfrBfyP2Jsd8KA1hLDib/yWyBC3+ksw2Ig5616gDzMvMesCjDi
wuepITruK4zU7qBR6H9r2KwXNF7dpklaRP//Ol9jW9oqICQYyviRzKSjbE6QtCkX
4jp2/ayV7u8jA5hkDwFISUnmKmCadvgPxoYdYhibuuvZHRQt2uNNTyGBuFAMGivJ
ei+C7Mb0sgetAglfu0L3lTP4sSe2EpCFvRcZmF58twx8nL0QM4laba3SCzWdQ2Rx
o0pTipJRUlRWu2XGmuT0tD+VXkne7e7Ym3i8qbtbEOmGEIQcHhob6p8PpAMkMNor
eKUchVh21a7i+zRp41msdzB2gwoY/rbTBYfhSeMkzUSuzTCP+wZnyJ06DFE/2s4b
leYtylrXnBmt1hgOFloKzQgMp8k8JOFtU165MiXiCVhKD6epMy9m/wJLeSg4C8Ym
a1/h3dL8HbZh27agwRGJlvnDQ3uUnhqn72V06vAZf6GylTxafdXhtR2s8POKO1ow
go5U9WohG1a1tfT3ob95nFmPo1wsl1Unc5AGo7giB2QCEWDi+EySA+nBKhd8+8me
DDnbM5CGx24ikKNd5mhlBvrRHZDc1PhM8KdIwR/TuoW4BwvGD0KZaiL8CYFdcw1h
Rlb0SihU4Fkapo4oA3M7Inu6dPNeVNq3N++CxDivf9mqnXyRjl2eiynvqcOxR3M8
PGufZW2TDRmKgrtF8btTkDnfN8ruDvPg7h2Fq0Ds5Cc3peCkhFJJGredg2JFlTO0
a0YGSV0akyKEqGeGn1Nfj8YmQUZmOi8WADId4Yb+yJT2/Ly2NYvzrbWiKKG11TCa
KSjhLwZjlU/cO2wK+L8Qq0tiQJNVde00OuWxVkkf+HHiz+gP6DUeEvp9QPwg1yFa
CBZeDKK/OT/m7y4zy5HBcoSaVY+ayM5b68Expqr1T1jJAox3IYt3QV3JjgfukY0A
ffW/Msx3HJF1XGUN8zvph8/nBon/RpHy7cXSXyZLRSf5Y2m49Xyh9V1j2unXAkOl
P3aRCNtu0aCI3EY6/d/PW5EcZ+zUzJVwvOPcwfGc0SU2RQdpyjpuoIl1DSI4Jy4F
UHAhawHglqArKIdFe0wjF2cBdL8zYUgO5L0Q8Om+SSA7UVD9kC8BIwWruFJPN0R7
MhjQNn76Q5rd6E+oQZXgWVYvVyI3teNTDf2niVoNbLpO0h+r2IVNH4G9vZnCUvyc
CLiM5oVTuZUGdKQE8b1JStJ7CN6DX+pi4t9AQv5sZC0RJSvE6UO8/yE0x56A+SYC
mC3mHbKdopk9LEJMZJmsxITqhevAr0eiM06lz5kOiGwS0xbM1wzE0ia8UTmMDMun
8i3Z8x/kWjDQYKVc4y6ZejrBPUSNSmAgcouwA6Im1+9RbGaHTN6Th4RIo2kbMFQz
EtbIwQjx0GoqXtaWKtDT/agVDmkKa5qOf4XN0ODdE9eaHL6usmw9nU2OqyUZ9xWF
W5bLLBgY8eWy1UWB9TkNzUoCN/EDIiUkmXaTRb/TQp+hPF1JgD+pxznZRN7aJ5RF
hB9TJ7Q8BM0Y0hCuz9Suxbc4LaufvjdDEad0gurR1LKIHQ0mEQdNEE9jLx07VmCt
BUipsuc15Y9YIxuYRJ38WzKCeDGa0AIvGIPqyYIIyQ/FAX16roTZ8d+XLKBqI2Fa
vS05O9Gllz9D4Xjngz/y3uHkZ/76ntbFk9h2zbJYyJOJiBUrG1iMwsFyogg/IoYd
tKECQhh91C6CKZtAIBJGUJ9jzPQP81NGys5N66pHKMou8plBNjuEUttKoBzDUvHb
u0c1cxmw6TpNMqgp1RDqUm4xTFMQ7VSD1RP5kObbGYPwWyUqF47YqqNpKt21LkUY
dMWXTh+7MCoOea2JbEdFNG9qyuBs4nDhEHejRQhgI27qUsb7h0xLP2u0hcy9N6oj
M698x0AXP7FDnODT9lf0nr36xw+zfAlyG4A2MCVBNLtGtCyOy75rAlHq+neiVUsS
CNvOY0BfUbq1l2mo30B6Zl/NwPWr3Y0JY7pdNLCILeydRSaZ0t+xL7jJZkYz3P9B
/7H+W1UyN+4aUiT9/vmrrqXXMmyN2bBuvZt+xB2EV2LsMrW/ZL9xKOyhPXtKNyJq
j3IM5N/TsVGANt3s+HGAowqR+dScjQFaU7AvxWMgENVsAMDvRb4xS2J98oTCtq83
OanSJ/fLRcmGVC75BBKu9jlcEh/sJQvfAylCZsLbpakRMw+51N9EGsfsJ4hnnmeo
ACy8sck8AErq80EP6O92aLf/8HRIpRUdXH5iq76Ol+ty5SoTPP4SncMc7XqBIuca
ADnuGxu0/zceiG85p8hU3LQAMxWr4s0WfSSDCrEq0JV2jTeWC6t4yd2A++yF/1yO
/pC6MA1oYaBGDBsfyegMn8epRHEvv6fKckKflelgf6FEuuHeMr3itFwFPKHIaPVe
2HcL7JwJw+XG6nQN1o4j+1RGKDly7Ifqa8ZWbNnSPxiJ0KkRFdAf2RKYsm3df6Hd
cz3fnk2oKj7L1ft3tGTY7e2TpBuvuFYb/MQjwiPeNrpCkKARlK2BpzErpS5/TYn6
2o1r0T2sC2YmDRtq2e1yKlcK6Q15G3iopcXjAT74W1+V3OURHWuS5Ta7rwQ9I7GY
7LZFeqwQS9eqvuV84+9XDBWdL7Asg5Ub/FH1C8KyH+wEhgygR5Xl8oLg/cSvYz7y
5witogTigOgf3od6m5V6r1U/IUFgiNgjspZ3A0qJVc5XC7tpk2/+gPa/kIyeHoGK
FyQGviyAgaj6jrgMwqJ7sQFeJd7+3u/3CU3nxqzN1nTo3rz6syZiLa7w5ZnSsykv
7Y3CJ4ojiwbaHXuaeBrOyvt0uGjy8xSD0YpmJQZhcPRjKkT4sEm6qttKYFQFrKyo
asr8yC9Dp++pO3bxGW+aniDvTsxkLNZTlZPIp8TTpu/bEUxjdT8rVOtYZP8ixfa1
KZplCxL67A429PP7TXyqnukro9JbtTPetu3RLUWIJJx3YfzO5/JGgXAewlrjqSQ4
lugVmud1KE43L0oChvcMQ/94SB5fanGeSTrIM6TKInTTvn+DCwQGoaDzYWlq/Z7g
DyG7RT1YM2yKL4o9Uyl64PQZ9rNZrOQ+XN//INNPMe4o2T6aSFo78H05yX7GhMS7
2sSZZNEgzYF8uklnFWMIIO0tcbkoejvwHNNvOMd82knfqDZ3CBe4TgBYiE3VpY2C
jacHsGhpnkE1aL4K0X8fF/kw96LCtMkkcePveJ8oaYOa+KFLBlEvP1bc0TM3xpK3
A7VTcxlGOZdslyBKsVjhPQshXOzR+tak4dKmDtdgBM3aZPjZm4ClGY2k04EtdgI+
FJ7ASt3XCdDM+TxLiHypbG4/pptTWF3ZC9lITP78uddmirOfxQ+CPp11TDvWUAax
WYziHDU4tHGN+y4nL+5PuwcYiGeCcGMHyhlFfiRVx0wtCJhrYUXm9CDMYHL3rX9L
F6eSHAGXUopkuGHd5GcHrUz67ZgNfa7zSsTJ3wocHX6rwIb0JlMCMtyW5Mhz7LsA
R699MYAENY7blS5BRDd7n8WFnJJRVUrZs3Wbo2X7YlE6P1d0fnb5dmoqLhpFL7Ay
Sdjzr8YWe5+Z6mGuvQ0uiu+eRsF4GvqxmS08EpLJu9rQu+zyq94zef6YDmKcDsPv
NqFSBkexbwSg1iCCm8X+6rYVAFNsonhU+10CknW1C+uhW0yUaOrfyaD5Gjd/NNRU
kpXpO5IAOMk+FTpCFg2Xlm7KiveVj2w9QVlNn0Dl4HJeKcAETvRofjBS/mPcYTMb
dlbi3HpG0kd7sYbF+8uPKJMEe9ads7TQzD6hqBbFyavMPh5MiE00uXlyeGxriuQs
Vp8Y7kGZpbXgJwA48+ONZu+DaeAxOe0cht/J/xCjpY0vFEVrmk+j0y78k93Y/9jC
38RkdE18tsC7paJV8NiyFOM2UwbVrJ1X07AN1w8ilpFFItnqtKU4e6pFWqnyMmOu
MEhlsq58l9AjGmUFcx7kVL1sXVfcCOZtGeeQ1JytucDV1v4aItt3/UIKBAemBqqI
GP5qvkaOwRY9AqAE92eZumyBfxw0W9pX1sKKjdCLo3Ao/58XwZIDBOe/+SK0pBbu
Q+ifandIYMMylUnt68I79yV47VWXNAwGUOrTVkzMImEUsxvQ0F2hkkCiToPGDb6/
UEPf3ZhGR1fdWwMPpWAwO1DVRLTqrrHrypTiT3LphVRFIBphBdRlU3/vuDMkuL2l
ZFySm12noVL+Yg2PcklPdvymg4PMsaL6FEVvgsB7lXFUbLz5kzZcWmzcxiukEB2V
lO47tdXjFl0pnXopzrQGbFvu9iM0ju/yvfGs1nIoyZbr+41gIQWo6ghOly/RfPX/
BQm9bgGOl7EyFgJgvu+uIZpZIyua6N8gziZ5hvwRJcpxro/hzcGeY4cM5f5D+RFF
QxyI5/ttKMhgpOtAmbqE8wWvOLkcr8aAcvitc94PP09gjhrCB8uZF+u1h8/dNpIf
wF3eou6aVcuO8Ed2JBmhbfZ6VcAeV6bX7NrBfCpnv7lp5JfjHrSrLYNplVZTyd0k
WkOwjhgE5kMiTIoS1XZAZC/GmMafiTF/tvAh5nOK56F7gYWa2DRoL5WD7xCF+PHP
BrQ0eIix4huJCVJ8war/GXbUIJEbJi+xiBHjR7kqchigZytSyJabtcwEzglyuqja
29BiURtdnHdFh3PPtx6f9pNdEOHoLuOXdt5whmLDgOm+igtKfQ0fJHg85Z8hWuYA
h5kGfeHZ02CmqLgaK+WzfJ09mf/p4fjjkBNsOHLYp0OAbiUCG8txHba91m9wuF0Y
+d3RLt4Yaexge51Vg8FrocCRuv/lOkYURZhlbS8ijxhxXkIqL8G7p3lw5a9NgCoy
mwvUQSwyNiEFql6tNy00tA/Fbn9gVg2D7mTN32aICW2Meq8zncROlzfXCvTbZyZ6
r/UooT1vR26iBNIzQf4Z/rYolgaQaTtKiNgoV21WWMGKG3Crh/LtHwm7YTAfBXTC
DYWPMEeu80vFuykziz5DSH11QpC+9UlCMGcmdQhghYOX5oBbLDO4wPRLtwB2T3AH
n/DdQwUIbc1pEIbciTJ2EYxynj2hQZ3KAiCa1MtT/ivff1HjJdU2Aq0u1Kb5Fsxm
Dp/7eXMc2gtqah/DM0K037xRAA8KgVhYXZl9yf7ZpxkuSotcZwySK/P2yDdj2DWg
wzbW2GcMKdfeMr/6Jmq05h1AFtvhbAYiElz+/gfJU6DMwdN1s964HomtshvFHYuM
UqXjmIBttchyvmm2Ox9+/Res4xdJD2kzBrxBdntHP9IDVhoIWLWhfYxeUX8Xf6Rx
gs67+xoIeexYVuSNj+tadJD0UACF+OsEJTT7s965u2ORr3OaVzut+/cmGMT+gOHd
oUEIiIO1kOm4Kio1jUOC/TkxCA/hTvWr4HIIpVat6hJy0WNxssndV/SR5Wtv7Dny
4KSoMycKiihI2qiE75jCH8Sz724+npqczVKuI9qdC0lA1cuvIi74NSR/EHFpL7Vi
Yf9PXotUCjJ4BpPKpDW++wJCu2WiaVD4DzViRi6tGE9btv2O2hwhrktztkFf0bZN
fvNPj/2EnuLn0iZgXQKxKZNOQYWEwMcdlgeMIJFttJPZqF+tnRtYHeWXLR7Un8qC
oPFwtKijRzfD952RNeMRFYyM1P+MmTqqqmoNuV+RnCzybxOKc7PHagqqWZqFm0DA
ImEfR7niLN+tO/CmzwAdPEb+dPdIKENCT/4rHSsPr/jfLn9sB/pvOngX3Vu8e/wQ
HWObsxh67DfPq5Bw0an90Vblvz7RXNPREqH9t58be5FDI2jf6+TdxdpgdYO5vVGw
VIi0/vVqBTyflfV2Cu3npJIALU/4nAUV5HILfm3+GcSLMUTSg7eP6fR9VpN50Rjq
D20cWEpfkTTpvo8PoPBQYm+mcmjdtQLrZGY2qnQ7s5Yz0ADX1NIWdTjwcOnzhVzs
gUI1JWT0f5cx6Em4/I1O/RTC4yZ0OQIIoSuEFiWfciTPisfhVwyB6rniKU+NRmIs
cJJT5tSRgIf/dhZBrTj/1gXZl60jNalHkzSFqClMc3LMmppNcovTfp9c45Sv6kmt
NVtf/CEnLuH8zXZ+ygQwhT0HoFSZqONpIClOtSjk4vmRabAMneWKvysdwMKat5l2
akKEEZJxg/0da9BPNtnuSOI5Ju5WcvX8BRKx4nk/QS4M0ju+86WzBC2oM+BeovYD
nKnyCGC7gVttAaV65qGkD8Mk+1W6jfHYCgW1G/nJgYkFvz/GdOqIUDYS7DnE1cUv
P1vJfrKs6Vd0TrajKlT2WHzM3t0k3mGzroEmlJ4wBRJc1fTrXAlxNGwGJahFM3si
lCNpUZAHOOH2sk+AlpsgVb7JxXUyk8jHYNRj8sURDEp2Kqp66p7z4oweLQuFtMqd
jxQ1MTs+zSFaCTcBAwlVD9nYDODNkyss+z5AyjcfDrT38n8Sr9h1SIxtAdLD1plp
/nk74paIC5JBhDogFxFI6KS/JmajJtyfxC4sSiZ2ewWiPjL4i3NwQklviujoNqz/
KwfhqCMvsmwm0Nj2tK5LuFmCMg242wRvV8+go84lrHvaK0r+lmJF4AYIdGDpWtro
drTScxv+6/2xtQZ7eATQHCFD5jai84vLlemYc+ngA8BsfKWF8U1z8TBFi0Fm1YHx
nwJ1nWEZrd6H8PLIUrJ3njsz6UwU2v3IME3h8YF215i4/Izx8HNdnw2dtE99G7rM
7IPrxDgRgWMsVR9I0LiRP5KFM0lhC5tIyJfFswErsgPPPB3J5cNl9P8HawcLWLyT
YgKKql37FCXqrngtR3TtqIAIMkHbSfRMTKkUnLVKovkFdHDw9/Gk7iqaFZ6HoxS7
//CpLkB4z8u9z0fjMRC7ZTFTh4tkN8BzcjQpAp1ElOZSnBRKoeW0cwWeFZPb8e1w
ku8/DtgrNQ7HPHdjUCIOqYN9+dC86pJKbRR+cAv7f8D7aqmZqj6eGiKTFEAawyeL
93dwVc71Gns86oUHdnmx3UomuxqBUKv19Bj9vMMkeRRTRRywzMrMh/mraESuOSDW
KESziNK9HETUrQhfyIcJHM/Edk5yuGVTuZlz/J2NilfHAhLG/KHvZekaknifk+XQ
xV0o5YVMylB9h1WHJSodrvEjl26QXN0VkbOckV5hocr1u9pLdN2rTDi2rvBTWhW1
uSi/2n6dfQsWN4Ry1UfElFhj5fizqry4J9XZxYth+VwPsYwyRhhU82o8I/8but1h
OrpizEkD7rIwKb4BrKgL9KDIsgQ5DBVDpuaTFs1MznGP756TBcakVv5/BRCIVOFs
aFEaIH6pqi610xT+IlXIQlEGLoCcppGColMASx92WK0EXBZIkz2RA1DyicnsNnFZ
wN6rHIal1whKFZllsgbsGhUNQDuEwMqujg1Dw5ASF+1WOlRFvWzW0ZtWFjKRCpEC
ySr2/VxvNH4gDOKSe2JePpZ3bS7c/zhCk3uf+eV7AAWrGDgOclfjzDGtUjHOPgZw
UMbrRWFbLQCXXnYq3X1hKDPaDh89te6SnmhwiQ3fd2iJJSwr+D+YIQq2hIMJj/Eq
EK5vxti7sdtyAQNO9UMoZQ+/luqv6497gN7eHnDG7TBEulFJgtLWbEv1c9zPWQ3k
9hq9qGsI9K1cGxWuq9IKQBME9AdoZCxFUX8FH2tVBVVZMeV6LVEdnsrzcrrDoAPi
Dv+a01oqE8TIZToOH698yhYCkqiQsyymsLbwDwoCNSZfnd/+q+cbq0GJDXoQC8oE
+WhZ2lm8H3KTk6zNGmLEyvU2xrju4lphkqoeQOZz9sJOTVldhid7EyUhUQZasz05
lJ1B1tyJ1VESO7KcR+W8Wr47RvZ72592CZOYKBx4b+cV9Men1JtSPj0XYfg47bqY
r/pJHu1AVHEglVWKkyQH3K8QgNObWTmP69UC/s3AUnxOqkgIo3flF70ndZUKZscL
i0Z51+2wozC9oWMemAcIAQA786nIxQcLNHxrXjJdJ2LVVlRHIP59O0ddA+iq0t2X
6J9OtT4/lWa3pCOOH80gTWaClXjT+4JDSoTVuXAQowAVUi5SaLA02hntbh9Cv/55
fh5tDWtM0GBnhoR2MRnSj1QSoXmKFUINGrdR7lJWRvl8sS5Iyd4gxUwkyt2S3T27
I/4SRyXhKQM3SOB+CUcagJOLxryH5O9+na26/y8oPYfmL8WOUoiygfTy4zLpqPGV
B+kQJoLNcfV0JU4o9OKzQ3xw+4N3z2Vsq6PhiABqPAaFRgb7/vOJ6vJtpVb4201j
O8r50+PvnWRSLgqu+VRxl5BPNxZzVJbo7vheX0V0geU9QWfXc3QyBjW4WjRt0DF6
HFV8v6JW+cjQFQ+IsRO+DNQq+D1kPuuRrT4txWcuYKXx6y9b/vlVBxjzWUdo4gdk
Hoy4aBHCuVB5rJl1siKuRZBnKBKgJNyRIksFUMKTQSQUqqH6+gDwXqSomGkZhEJo
pN2OdfbOD6tQjVzKZ1CVtAoghK2u/ry/wZEpCiHkKKAZC/LTpqV35ob6aYjHFLh7
/mbS6ehy/1EG+qhWVA4jjIFNc+klPMNbi5b7bwZ9E0ef/hfimhhYl2C6PdqgAQii
qGd8VjXrQt/ALW67iTIsev9pnXHne3T5PflzDOVEWS3uT06iMy8ZOzYPG03X+y32
bcuDmc7n1/InZAuAUq1/mHUPhIqa9Ce3Nr26oU9ckEf56EDNJoX/Enyt4Mlq9MFN
7Sva2R/ElQnwrrC+14mfg4o25AqJvAFvMPdxc0BZm/4V18hrLaSrJW4rb0ptvOvN
P2by1ML14OzSCM4LykHe+/YgxXDzYtneAVasxBHNYXrAKN23n+f3k1j9Tqfa7Jp0
6zD1DYdN6wogrqVGu25Mj5hkfHbMMhwLzrx9Z43t/+dS+GrOUZFQW8RWYCk3zWHm
V/SuJUnmEmZjicc90lQaFn1PfuzJQ29kahTvuKuhPy1D+crtYapW9aWxHbxMyKVx
d2qhMV/XvlMTImJP3v4qwuF/oS35/7f7MUrI+3Ab2oRGGpKUEsMTXs6LB9hwxlh0
c2Q9IhMV7yM3dEUtnXW8vVMYSGKMDKTr0m0zVZbp++dtkcZNJPihL6S7UyKeiw8J
PtRJ7z4mq3JFhfu4EMoWyRpr4zmMrIgXFO+oQ6XsGuKiC+lc4/c1/fBgvMaE7l28
mbZ/SFYaPO5kDTTOGXBHJ8tnn0H9C70XRppx5Ar7Vh3n/rWEeyFOiWJcnaZP4/MX
aFozeH5ohs2z8HBKDm0+zmOL2hQ37Cy3NSL/uzn5eDpn+hqI6+KyGoyprKM0HwAw
voNnddywLVGtlCz5q9BU7F0BDC8PVksrICCPeAmdHDn1+AjrUl0nED28ZOmm2jdC
Za2U6SVaLFJc9m8YSjY7IZv6LQG+zDvrnsTRiEXO44zTrfn/D7TR4amQEwWjoTog
B5XpBAgBfw/G1yVE7JGt9RG9owu/ROSPyIHx9Mr80HGfr7HpvTyaoasKVdvVE4GC
R+/2hjof+FYvfHApbqMFeivdUHc68xUwXYIiMxxu9svg05jj3mduwxLM/FrOKS8k
KZz57TFDOiiYI+0SGeh3l182oMrf+8IFhsiCrzILgekKPdYbC9iDT9qVhgyUyWeX
Ikvt78ceAnK3Saj9TQLbPK9/YmXj9yKXVE1NHIHU74Ec0bzaoFAoN8T5l7SljADj
K7YRBbaGT8tvS4LVH9FixlkEICyjdAq94QSi5oS+UkoFrkN064SRe2wPgNhELvOc
la11OMjh7oRewxduvyYMjP4PgRBcgU/pgQtTSA2uRvtWBdqBKJKlN6CYEbTQA0ep
4MlBslqbMQlIheWDpDrDMWgXyMloSJDrQ9qK9mrlgl+5a8iw4vPPlUW3hscrCMRi
5gAvCCIJdZPY5UYN9c/XTpkJQPxBrbx1bemzZc2c+9wBkZmTsbCE/sU9ORUTII1P
mBpp9KkDHAZADLQXO53VAooL5lsU0+x/jhxmfjaAuw0m9GbtXckUC/pJP20xB065
lqh7hKJu1mvBLSBa4BZke0gjIyk0yOrn+sXMDAUwzbbIe/T4eXFnaRsx3keS3geV
RYD2E2EP9Qbwog6ubnsU2sGWRii/qyr/fqe9ChQoadahY8TYNJCp9suI8QaoXfyi
MD48pziJY/tdrISFlbJRB14g7MTVy3HmZwEmU+rGXnzK2aNyBnpc0o83mx0WYTzU
UKT8Yf+tznGlgQ5doh/JboJZ0G328Fqz8qSyWkFQxlhrDfXb985rqp1eeRk0SRj4
8Y77XXKVImLRBKYBK1cRyMxE2DsBGUvTtc9ANhZW6HDzvu+x/2i4TRYrIRJ8TqqT
XKP5yC6xJEY4gjlcXo+TGoMp7cmjKDSchsCn+sV+s+EmhI4Zca7lu2ev7w3wWVdf
3gpsL8PjDHZhclwxm1VvAjUqCiJGT6exYB58nqETDbHHRmHRx5u21CrnEfIDfaDh
FLpFOAFwk2+wTxBdoOzAwiTSV0NNt4OknV97wlLHXR9rK4M18KOBbujI+Sfcy+2q
KRFqyMGlWqmrEwbzBpB4xJK9ZVEHFVwFV99wwD9ZYDYd4J623WpQdi2QtawgK05M
wdDkY0GLjpp0tCP2Lx3QTroCtNTDS4RedhhCIjG7ggvDxu04jN9BKnLas5WKecB/
CXLBLl2Zn2pg7gvO3zsia+hjNeAAgNzrqlilbfBaKjLVp7knga5U3F14g9aWQna4
NdlcCocMdODLzcLIY+f/U4TRG1WSSeHDlozKC1ue0J3E7Xq+dCaW45t3+HBJ621v
qVKXqbGnQJ9NbjmJ0wFllVlVzgV2k/Nu/DfS8cv6WRLyCji39yfIwZBbAy4Z4+Mr
PhNH93gV8ovr+53NhR2Pv/bmH8YsuKEW+L9neJcgTSKeXxPSL0IZE2B29BPed27B
UcaxGPDcLenFhDON/L7D6ZzjPa+PbW1Mc+xhZtZOFkyulKE6jTFdgRYOzLobhDkq
TqB/uxlmAE2yMqLV0Q5/skU+q59jLno70EaObysR9ObQG2qJUMOT/9hBfHwkdi3e
vSPAQCgGlv6q9Oo3eEcDEapdq72vP+L+wn9O8XxxaLkq+p9inWFrQ6ccvfoWTUbx
g+fJB9rcU1pgh1ON2+KmdJGXEgCAg6e8qEgBhoQQ/3nxVrPjQWy47NCt0tRq+a0P
BqNv2k98m57iWFHi5dyTTgeRJqv+ngPCMBWTs2Fdt5OPuS5cGvroXJ9HqdBc75lB
UNnT/0VKtGz6laaYfUkclHxr7kOtVcKrunDi5eZl1HUWOJYm7b/alMtu1ohxZPrJ
V/PJBQnAH47gTAAPDrEO5THFlwq/QhxpAMkLNcHxecglTVIBOqSFMo3MCrEuEfPh
CLkmz8PTLuK+L5ZKI30Hmj2TgGVLEnI5hXARoaLWGEJcQBuLCm0qyG/qU5xysYGt
Gl7s9Tu/XhTHAJIKtrgIiEGTlujYNfeFS+ZfARCcfjDweplvQFykQQgHEolLX0PH
cy9hl8apaVMABtHCdbStyB9yynZzZF13jp0JDinTUa5EGD2Y0fxw4KiXT3Et85Nf
XMW9g7ZqOx/31mbBrJoDxiQ9/i4mWj59m5JunpNa9PHowxi1tcZvYcQ3YBvvursv
lHUtBAEsGWe0Y/pLdky/TbUe8D6A1UlDPCXM4+tG6nArzYiz7PScFU6fwQAn+DAC
LqPoBKGrEdZGPJ21I/502wT7Z58LtaFZMMhTcuQ2IoM/nh8tE7fZwV0cgUxp3cAB
lOp/8KoThCd3iVvbsA0g1szdLVEfJ12LTTlXqn+GYObq35respKG0ESoWstb6jn1
/L1lL5QvXW/T08izW/rbYsygLbkvvAW9HpKlpL0qisPB4+OCr97eP2fs6MGDX1rN
llU87OInfo+13158R3kOgkBdsZoAlkkXKkG20AksA8ekUFzYK1uC0ij8t6mV0R8D
NRyWX8AhavjIhWwSBmq00HNM19u8Q/ugrfQ7v2ee7VH1XamuuRErJF3H9+4fyjKH
rg4pZXNR+k/emo5xWic2I38fYUls6bkIPuQA0rk5Og0U1IjSOP7ajbndAaaOwgXw
ocBHTtUoTFlUSOqsPjGYCJs/JDBdPEjHvo+VfBKuolJ4XT8yNsElQ4CnTcZUCtEE
z/Ec6dQ77qZm+VnO9bRAcPNj/rBIA3SM1KWnB4XI6lToEvUTlzfEexiW7gMHfcJq
TS207lOBB+dqSVTn7AAyaZsou7n0s0DIgjDZJARJuQkLG8hapRlqS2PoPhXRECGT
Sk/qsDMH5+dqdKqRIMH/7AVMiEZiH3/S5A9CqHf1Yz//KM/C5l3ar/moBkSzxIAt
YOUO16gXQjrXz5bpoTWCk9axtCv1uQlFhx3c9Raa6vBbE8ygnmmdhoudYyck3vDl
U8cGn9JOWInEP3rSOY1HWu0WU1vZ+gdyCNvLO1Qn3y1HR9ejZdX2RIuzrrB13vmi
hVvpmiJt5lTq2i4nqnA3ZKz6s+EQE7Mpk3oobSY0gVp+gPljKJ0XZv1B1+ofm9yI
INgbsz5DgS1PpPq9ldxzBkx6sC8ljVackt3zZStU3GAKq769xtAE12dLUpmW0wJ/
pLmYkE7L0XJB8Wg2BXepf4I3S+0rV74DJR082u5EwsxcX3kBVTjCWrlJxsqOZib4
kRl3+1phWv3CJosKJNQVRa9SsJoi0c5P4O3PYsYCN6deeI4zGdwaggqg7fiwEbgr
Zw+GLmMyczkjU6qZcBdosAU2pD1m6h+UeGblG+FglM/NXTqXsQU0ZXmWNb5rCGg9
9NaM75MxI3zSyvcJRstTljELIQaXQoExF7r17jnlezD1IFnumoW4dIWpWLKfHLZ0
gFOyCgW9S6DbWsS0TsVtObEMJGyOP3v3T6J5mVJy2gAu3zdFBH6rEMxFIq1WR6Zn
GDEj5bFjQAdNoJNsgQhXNA8IAjC5b9W4A8UwChLLtiSH+wVdF6botjeJSFEm2rsp
GgumNPqtQN716GzzyQ6dHSQepVaNsHzoJ3znPKo0tDEf6DBJkcNgkG/K/rTPRwuK
3v0GW4jUDQ7JYyq1aM02Xao+Sav73nJRBNADaj1ELcOF5N9bJfTdjA4OD+qI+oGY
42nsROx+kQiF8/eKRPM/ClojRRCKlOtjgLeiS3GSHtgOCwiudO4eaNTjDgsPr3Ul
OBkaMDPalgEUniJHhe6NPKTQtunf+15+vM/W8DL9hxSMfRXs09+jiyhvupIgjjyo
ZSmUpeThiNIKL3hxR9yg0aJwKI28V2meXMrrP1sjiyQM5hUy4j2HWnPTsD9sNXq6
ouuUqG2o0glHC/vvzAREh0+SzCePbHdUQvXCCI8K0XxKVTO0weKde0q9uusWIJLm
XVpLMpj6S16oA5BfeGnHgZWZZlSUv+GKlxR6jbqSwu0aU0QxBHZA3bT8oe1HwH/Q
YH5xGbUbgES5j4R+3geuVgSgy6dTR5qitT0BgAmQtFPbTnHEXY2MEGG50lLiRy9l
QMYeYd8IIr9vVooOoGr/2xOW7H0ToTeWZOxjvWK2X3VXuqlkmbz5kZJTizMyXOtW
fZVkvW/DKgfdIPydodDTN/HrIhFy2QfPz05BYxE8397xECAhywwi3nnzpxm1FcSu
+qHbWC4zF6azrcvwnq8ZVg4fc0wO8HTPOp2rSxtWBhARu6NbhUCE2x0KOac1H150
UFBA3SMGH4uKmHWhSGD+4p11eq1qAKhy7R/i1RtfeT5BAWZMgMseG+rL7opepePA
GxZF121ZNDsD6oO2/to0xqOf/l9VkN6dhLEP1TFUDomV+03XmJdwlkyvzSIi+tc5
20/4aJJPdTAn8/DX9Kr2z5vVqJ36dFEzXk9svUK6XLj0rD2UK8WwtWbB8d7+iCO7
FFC+WOZmpX1ADTjrS7S/C8lfF3UO2/J/HGR5u4q4+/8Y+XFO3zjamukXgL33fo7U
Q39D/keR8W6P0G8dKtM7rlT6Y7i5DYHDF1ZUZToiSNM5jAG2Glc4dClr+yxKdIFQ
5DYo8bQlpwt+uEBPtHtl2Ouzuly2H86XB+cqYDRR3NY7GCVgCMChWfCGkDD5GFux
HgWM/8AIqBrn2zQc3j8fvffeISfL95Mvr6/YUzItc10CcqESW27yUIRu/imdny13
KXOBRZp/U7Y30dquYUa7+yrOBSKg+R5ToMQXQR3gzVvI5GalF68h9ZZCwV0qMeBs
JUmhZ17dcIVFoFR8WyMVIqmq+UUYjL8d7Ys6uFYxFUd+yAGEoh6KK69W0CjdgkpQ
O8/S/98K50kvrKzoVZMyt29z9K8Ct/vrQSKf3ZiIqIUe6mVkjJnx1mdFaMNFKyYO
HQ3Ew97a5x7okR6dPMuc1zeLcybxNu5AN1pxeV5RsYAkvZgXP3+X4NbHWz0oY7cf
q08fkni6ous2ZmUHvAjm2LSvrkWPT/gzfWluhxjJpzGojh7dPSGtKJucSkVbP8rE
pCnQHiL1CBi/IPq/hKCOh0unCE41OecACeZNmyaBntLDu3shwJQAN+CfGD2ktmLz
3LDPA6yGgE+1YeIMUTdHrvHE3En04QlpuIo4Azwg17d8Ek6dtU6h360/R4IDdvTQ
LM2v3FgM6ZzaobzCBWotTw83xuouOvpZrhNKEn3f6D898wf6w402kvRoQXacktKv
ItVCgsIj1FjV75NNvUOU/w+NbXZZqMFFsusklVoj4Sfw9y9azQWmssoI/zv4uWzO
kP0HFB380/K4xavAfBMF+7AGlFtQjlPMNqF0WgQoJda+pP++zscO6kHbpZuv6woz
8I5T6y4oQ90GGQKux4tY9ZJUkq9FS2w3iWSIRblOFbgFIMCYWrwHUBGRZ1fOtn11
7jQ215aROHesMzeegqc4xzGPpC5YKPmCJk2f1gcxXRZ4iFIPUrCi+LGHyqbdY/tv
K8xPhgCiuuWzW2j4Lz9P8J+dDcqKz5rsZGIPuXP1oeWUi7Aju8YhVOZk1SAluruy
BuQuMPJUqPTit4xFBM/A0uJr/iwtZ1cEpuRdegjK0oBPaC65ecaFcHqOou1tATRe
6guv+0YgjfUSI0vj4Xs0vhOz5DYg05VKyqHYsv9rcp5bUNjWfBF4c4JL+cLt0Hm+
YDzKG1REBpvvKqz4YUuHMVKJuMAlwCcHTAzM32q4Sqz7AJHP3xky5vSixPBvcUA7
77nGiU8jYqQIe6BQjQSrMDfcR0VNLMj73eUbq9NVukrmYCVS1ntNXn7m874CWUCD
tOnWYzgc66bFPlEG6vM0cr3ZAiku4f3gMujxdfrOBPTYWf+cHA9nLsb+o2gRqbQP
DXZaG4sSA/wbNQyEcU1iljLb+yXTdeMUrDRs71tupYLGj6102CP5ZWGvHHycHWgg
qx8GbETjJvIthjzDrZEnMDMRDWyAztUuleE/coAPU8ctpciAbzR+YliSX0Hx1sL+
9ZIMCxaCxU0G6QaesouMUnWbc2QHw4NSAULwMAICGJ4Yix9XWrWY+KPbI42UIO2O
WQm59DzxCg9T2ZSDygfwAiGVaLmcux4wRzGu92Bz5616GHPvw0A081JC3QO5vRYk
7CebcKhxZC3hg4EIw1v9OCaFH/q489MDdilo1FXxyBzQZqTE/ZsnQ3T3qG/GOeyG
SPQbtNgfmgq3UlEViNx87mAyvLdrRWsIiCBExElSy8MeDHIQgj9veF8ibRpWTtul
`pragma protect end_protected

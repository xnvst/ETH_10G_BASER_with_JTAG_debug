// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g8vTQ1B+nLRoHUXzJvEmhYgUuHV+HwrYy8u4KfW9lPO46ruDuMb5wGqx8Aa8HguY
p46fXx2YEbhgyxLcvFC6Iv1958QsMe3sMc7Z8QHRo1jgEW/1KL/WGyqFsDCWM7JU
t7AVdfwH2gv+VeQSGdwarMaCFDil/vCuy/i80XIz4Jo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15824)
xq/A7JIExbSh/cIY/ErPMt6kFWSNaoe9WiY3+N6fT1QF8kRqxmgLfPnN+LDn3QER
4XZ4+E8JdK2SGN6+qZv/DIQELcNZuKiq2DtFTw/iabb1AIvy+zOwKvGkN1jAddgJ
WZvoNUQwHXYFhJy9tQZe/NP0Vgo6TvNtbVJxDLCazE+gv8Jvcr/x9j6hwrWAigzR
Jo40bU1iOoLSTo/ejS/Kjpo3EFvGTsfMYG1MVB8ysY6STaXfS7vpfnuPELKK8eDx
UNZnrRIRcB4KK9rjGrjWvY4x8xfJ7qlXMpPNZ0tRPjwGi1Jm2Zb3dNsWpNS3+hiS
//u556dzDqkYn4eFotiSnYUYxU1B5skswzt52dHTqqi/WDZoKEKMgwrQcnmlimNA
9miVx3AlaDJ61UyBrYrWds0pp2bxn6aCWB8JqVKQF+sh5fMfJps2HeTqop5pGvYf
3F6T8YeqtcCEWtwe/ZeC0mWZ0zUuVyitjih0xaSXiu7a/i7ePcmSOQ0y6vLF4z7V
rJJg/2tDGCm7Ew6eeTb8dPFmbY4IjM4m++RabewjJkuPuyjSFXYLEpMZyGYsLn8t
IdsaIrxubRel8JAQxm979lTZTfZJPq8YU0GZu82JicOJD1FUSm94eNZ5gjdh8nBO
c6TGzssV63cJ5hQBKvgeSynLqfS/IQothlzz9JAswq5U5e5vbTCTOXOfgQgn/fqL
dTP61ndO5U2MVt9odU9RoaDOe+fY1I31enklq/B90unai7xY4TsrvWBXHCMM0obE
1JjCagWfx0Oeg+F19V7tP3ssquGM6XsgVLffVsOLyUVmmBsrl9v1KGyx/0bf4t4c
8GhkzkHjUpiRCRnEyU+W11aYAc5i/KwHI7eF8prHqWh/amQELeRVFDNuNPSxS6Jd
/rDXiLH9f6oKq5HEX7IrZ8I/MGq7IJxPEspi5iK/9rn+qLXgbjB2WWcEcP8Op2j3
BKqGdJGOzCbvlkA+7T/xUdvHHPXwkB2kh4Lh8O3KtOnlKmJyY4EI2mTzHbp6iBDV
jpHuWcrgIVHwYXtYuPb4PkfBy8nzXIe7h6BCl+YCyP662cPBQKC/JeRYdpEd7yjC
itvYyf0OkgrMbv01ylu0w4mp8dCajO0h6a4b35e8Lan3Gtf0zu52R6x1nSV+8YpR
fv0Rkj8MLhV0t1tbijUq/TiR4PkOy1f+TWmtJandcCsVTcb+DiYDQ+awYYCdU5eB
Nsz3Vm3R7U0RXh7EJNZI3aQQx7gjhX8vHJ0drWQ9I4+/tQ3nq8QYUCmhKe7i+1Jv
jKMBoihmGb1QVxmgAsTgdMmXYO7ZqS9xy6itsXioKTNrAvztAYrgkmYq0wyZWKvm
BECitK/uEA+kuV14NfwuJ5UJ1gpVAleT6UPGXBuh6H3MOSoeRu5KnEKiyduumONT
MezOhBaKAxkCLenY3XV+5+Fk5MaLHxCLhV3BDphp1IENaMM+SGPyFpLIUTTaOqM+
Y4PMHd6vWw4Rh0S6bfuKGQZOXVEDN8hEPPYAK9l8bwG/wKXZU5f3f0TvHNaGzotC
3jJKOhcb+mQ4/RktRQ3sEftp7qwE0kZjW/v6w5N3WJFdgTpuMrdCLt20X6at6eGM
Rd7M5MmjPy6WX4ZifuELFXksIrLOVaDnFa6+GYsnM1M4Z6St8BNFvopE0Yu1+7dr
0ZuwAz/f5RRCvLrVMGHk3H4o7cvZVy8hsE7nVTKQieS660lXdc+m3+huqWM/HgM+
w5xIdcU2jzWGyuCQf+peme9LtAa1wtmccQsxzEO/xWsGdgaEsO9NTC3RTSQ39R/U
K+97BY3TRd8QneFH8GGQQ6mgw42EsReT/M2vjGLKj1wmmtOQj/hOHZ/GbheGORg8
Ejs63gIPitjSOxxbkk70DVfxHfFhDlkjDF2RsDenkcQQRNiGfD6FT69ENNM5bAqu
8x9lAexa0h7kh8SjLdfCXIEVQe2NRHIPxw/5cqguUjBDD/niOSHfAYFoZpmUfgf5
KO8W/Z5bBxRFwPDkxDlA0nVVH39ucGAhRs7ErWb/2JOVfnHQ7NyytjScTtPCALUe
PefDtKRkqPsgt/XFfrjBXTb7Pdt+3lMKIfLGS6ok7yVS12n1UL2DzY1n1rhOGJbH
ezsybpOaqsFe3zwvwnEPu3U7O5r6ADH3XQN5Mgu+oxJtI6jAlzzhg3TyDJeJ1FUQ
cPsYhzZqEYL0Swk0i4+qoyV9kKLJHaRTPRATrxxA/gz4zaTULcJkP8+9FHKLD4+K
J+XtBUE/9qUSjyd2/fYqssB1ir+vD+fMMWU8gFPrKM/99C9rNOmS/N6/2hqxGJfD
lFaE70nO7wwHRWrsJ/m601HoyLlYW4qMcWeed4ik1D6koGsKZJBd5EsCBFG50zds
4fPDwyNpzjAEDMb0n3oJcynOVDNg00fIK/50Qq65RyO9bVHi+zehe6+DVXZMKes3
QmZFhnTL9q6vrJsED1pyb5S6d+d+eOetiYYX6jnEMxJ2c7vSDjZxRHinCkzusDyO
OpwFXoqBh1MziZryXVuX5PWsZxPFd/hENJo9GvZbN+8uI3PFLBf8vgRI4wMHX23Q
+pAODHASmRTKlEc6sgSzz4OifzHc17ZD8l8WAx10uSRdiZo58keUR5xEyC+Ddc1q
XJR5ckTrjzqd59h77Az5bGhf3g5BsYZJMw6xqUmeYfl7PgF6xEarWoxXbjWCG6A/
pMhg0Q3e/3n8IlBCtl2gixSRr36Azgn97t94IOQh8WZ/LuEErquMjza1G14XXnx0
N4P4xvOdS5kShBsixjOyfRdGBRqN/nR1ZHGCKT77jh/GqAK3+YUyK2BQpBSKWG1o
N9XlZK1/Hna/KDdUxUBWOa/wv8QEW9fCM8zVCL4VHJI8uaHOSsGmsDmRynx6PpY3
xXu0AuwTy+hUvQ3179E6TbGudXO51xmcqY+wkFO7qO5h6SqtY25UHURj6+O4P2xH
q0E1NV0Q1iFxaH/1ODPaFxuk4zozkFlzS+Wf7G236K4ljbK4YcaydMLHTqSaNAP6
CpH5y69A0x9Q/BFow1wYAFubgtnMbOEtMR50Vx5soG6r0d6KXe7XWcWiepZCYS1i
J4dvN76rWbKQG70AcgfVK4EBqUu2SGw2+5Eom09suauqSnX73YruDEaQr1DTsx24
rQpV8TI115JSrAw1vuiB0bASVjA+q5kQqpOxuASv/t+eqvcTttGsazSrfIxKaOdM
oqRQWyyYUV7Ke/+BPOyYhzV2sJ4Qqdn3rTXf5t0h9Uh3hIwOmSBYftm5Qq8FOyo4
UuCRx5gMrlXtozKzH3fDhQXIsEVd66lbPMh70t0npcoLgpcQBGImVl9Hm8V/aMlM
n2DAL8ZK+PBTFToMylGg9sQev0LyI3TJ4UXJOW6uHwUuU9kUaMVgLdkJlcv2tA8v
CYDMlfXrNgRm0tAOAcSFjb5UowiRY8GhSFvwC5L6faK+DAjUfCsNF/ggzOSrXE8O
AH1cfJxf0uTvJQyKFc1q1X4eN9YcvcbQf+wQQJUudgYukWBW2rT2GS9U3K/cTRyj
cWFntXlaVBEw951qRvuZT9VPD+QYlk00nJzu2AtTbR+Xs42yqO+ohK0s8Cuufcjt
Xr4n7LeIqaLO1lj0V7m2fgwveAagGNgDvYwYdWEVoB4IDfcoK+cgnfJiNIWm5QA9
Fql6fSpQgalAUxdsmSJrvE2ibZR2t2aG4p5RNtoX40Usk8EKG0b1gu0a4PgcMN9L
8tg37p8A5B/lB7YWBlLNzYpNmJD5cFk0KRWnLCBNePuAioOS0CZCCUzSL/4GQHJQ
KOCxLpPNu/BVjglxHR4xntr3Et9QBn//YPHQahIu5shtFSwhKvRPsOJACWEtm+Ah
OApDUBa5sIcXijsso5hkPV7MklJtKCE3hlzzWwUcCfunFSjUDE2S6sllBXjGFD2H
qzHNeRtUo1cRkrAeRxBMvVMolTbHUEmJUw3MlNwjP7kbCgZyL6f/k9VtksjiZArC
O90EwPiXyO9OTUEOgEFJgZ4WR1TZnkmdtlfTZu9FK+nI0p41KBGBTb3Sc1dcVdql
D3OEKLMkSgdh71mUdL3dstguU6OIaqzB5Jco3H/xiDRKU8Tq8UWREDC9FXYLjeW2
rFWGFsKUnUykIQxVRx4coAZkHYoNl+WiGNLpIMCs3ZAnaDMBdlMaLgysft+eWXV8
VM1IcTjEygW3nx/1Tjzmc57EogE/KuHLmaDMuo7veeKtQEyhRj1IwYFd4HWdv+PR
ZI1emUT9nvg2fkZt25zKP2XyO8mEE1TI9qQwClryKtwxOGk1eYs58xyb0PljPsY0
tyIArTTDz4wqT98v0IJbNA78VMV8cR2CSyQ8ie31mcE9oAp8zl0DxcAOmz2osKQQ
8wlYZJqD1XAYa7qJVCTrRe++68ZKttHpxcqYiHIOzB4fJgrnh/1MldGPkwoKvcV/
I0RZ+9MKqXzJ4fxmc/vy/bX9Cx+MsNUhUS+lDAPkyTLGNeWOCwDKqdiaxZtrgA9i
F1iwwMWI9KIQd1nvehm9OBNh8ANkoVdmNbtkTL272tG+570bjdGXz0DnArKAdBTh
3fEeIwyVfl0UwFd5fBhspobmFcD0njdK6LY6eUGk1cVXWiSGBUdq9CpVUrLeAmQi
kk0Kqglb4kqkhUXiW57GpROyTZ/AnXv1pdsZBleNGuSOWvYmitG/RGP3hLibfmIF
WwF3MoH7Tj6YY4iGkDoOWymr8uWoPa01J9rPuFUJIVri3GZq+9Nfa7+DsySwJ2rq
V8Fb0lJXsZppg0Kmj6RNI4SK5XlcmhFbSvprdxkhTqYj28IK4A0nDczCIv7kcz6y
CnTtTeuqDYLrryP17is9KyrmTcWGffLgQZAO+vCj9QeESx93JSGK6ZY9bqz26phB
NqBlFhXyDVVeQBrZXxvQ5sP+cPeYEUOgCU9pV5Fi8tzEzWlXJdcdK0lnqTgqqpth
XLmVEkQff3QeXlOK999jdVZJgOMUd7HXv/F8KE0vXzhK62v7LLPeWkBF3tMr7W7z
oU8lRdJMGtRWFlSrxcu9fD6DZyRXw9Mq3PQONFViiHYYshE2qSkU8yF43lxJA0nb
dvzUDDJ/EJD8/Oofd2/w3XK9Ga+xbkdeT1Jq+QLq8rG7mnsS8OgrtKezaQUmeS8x
IQuMzGRSwlimHYD0dvKCF33pDuono85e//JApF1I88hPnYKX8FX/2WgQDWZ8MpEm
zRVFxrgZW8Ov62xSJqO5A9hvKDP/IuIBCmgKofGksNJr+lxUefjIESUlcTJFdK2v
yyqalWxfXjnZtoqX/OU5bkO+h2ub7xjJyNaDP/6xtKtrzCyVLGBQHVZMgH1ItfKN
+fgcvdozUrPfWpstVfWt8Obq3Z22N4bnkkvV0UCkD8yRxmIOesQGxJ0/vQ/vENin
Z/lxY4Oro9Py3dELZoU4b9QDLfQSJS9XcCvBX+Sm6qPlYHVVFpVlI8Vul/QD0Goe
TrE2Sa8V4vw+JilWTv6cNlYlM6TJv7Y8JBOz5qhD2Tns1oEo4hal4645jUEw+y/Y
yHWsR7L3MQO9e4XWTKui2viyqERWYnsTAca3rAf0dsd2vgwm80X03+QINFItcuQx
ufmaAyynS+bgGDa263XMf09M8gVjLo09VET0DfaFmUw+roKkzbwL6CrlftM6POQ2
ct+b3RdBRMLHklDb7Q9h9FFtj/BC90ZTEHU6J3KrLG9bBEvMVZpsZCXcC6IL726X
G3i7bzhub0rS1SIeq+rwqLMKkp+ijrxqBYOojGv1hhcZzCjcJvC8bNpL8YpOV3sV
a0gc62VsQW9OcHlL9ocBM1dxS+KgKJpbXN1lKipsnfxy6hY7qe2tnRcCSVs1mss4
Kf/uwKtwLEuS3tAk/AXUDdJl+tD4DxjlPQv+lpbSKmI0JIf90jm5+ihxJ8MrSQ9o
Z8RLKXnRvUTGo2CtDn/CBXV++/motEcdkUgN7Wrrm47uMHI9J817UBDGo3D1vYoB
aSwAPljY2dgmx1KZ153ainpwKaarH7+gVM+5EHFijIvu7JfuxCwFZ4RgpyfgHP+Z
07N+4P2jXrpVYvJYtHyDSW8zCvU6spnqrUfvK8jYY/HeMw37xuh2OI3Mp3oZYtCs
fkPI3r8BnTDweFQZaUys1QVrYPAEBJ3FgJ6ai1sEljwuGY9os9qloZMJ5btCu3t+
RGlaAD0nit9oa4ZZOSufDCA63LQl2U8ss16tlIhMeusjcNs4GWLhy005cYjTSX1J
sZSNQ4IvhYb4LxqlzRZDKHRa7Nh1RyPyzh947BM+yp7VuNUzhFRqpP29PfH4Dmdz
tVLb4G4TgZAvNrE18C+w7ndu8Kyf7Sn7Z5IcfNykovDfN6swWkMsJSfh9oqlaYL2
4Ki+RKuv5kqOl0eTw8yV1f1LQq3CMTbTt3GamwauQColI4/UQZUQKhYgAkNAKpkE
0t0d2AOecThM8Hvw67D5GLZuipJs/j4fS4uWHFynmvtsUbUIqS/C2qWEy6DmTDFY
S3ZU9s+W79YbaiK/DE1AgtIg26UjON7fspdIDL4CewpUdbaZrZlaJ52m25tSpZ5T
+CkEsA6fmT5ZGBPH0sobZd73EXPHVUgZo9gMdtC0511ciHLL4QuIdKq76UTfwzdX
A9ImiZMXTb1YpzzkcUw2eoe4bpgnROwvJoTtHg/lqK8BivQKWj+j6SzAErWvUhkH
LgJ1xQMc/LFkHhULKmhhoENm3BwRuT4Z0m1DwmyHwllLKT5/tHqaK+WOx1EwD2EW
yNnwqSjDbA3r67fTclH2rassIm8MnspBD1EzwHu+nWOLOwGCaXMWjcm/N4FpeLFT
hGDh/Ee4SsJ5aGZFfD//tBI/8tXAWRifw5EDHyQgp7zrfN0uJC9HEm0groDd2ad8
PqXffgROZFKi8rFrdS9CHbrL7SVuPnKVrpm4OmAQcA5aGE/H3wXMBzMQVn199UJI
pKbMH+sDYK6JXZqa4IUC+FNlnVGXUzZj7XT3oL1xjV3axFajCEdRAmpXpz6yFfEZ
D1142HDC9hprHAp+48SdhrTFD84FCA1qO4JPnoQ4Grn1FdPFdUaazxmB0t9ItAlQ
s9eOCOiJVjoDbpkgVEaBVmG+swrOh30JKr6qhYI70wbymxYBWBCkwfvjDgA9W3Gz
fJJO0mHsyYGlxSRTYdjatjbSC8ZJOtysy+DJosdvBUNWoQQ77Aam8xSVk5khB/pC
v4mKoQeE4h6rYq4Mm+wA4Kp6C2WuzSPBuY9KWzYphyYhqyIzuRUbOEbz2r0C9QHc
rENmuGju58BbhI+bmWx41RtxhmpdrC6R5XH4KNl1oiHy/oP3GBQpccMlx6vePwla
q19WKQakue2+qD70+t12p8J8u558wivD4FTZBDWHzY0Al4bo3ehS903wYhTmZkSR
l1TW/bXlGewYszEczvAQYtqTWV3F0hGtyHd9hlu/ops/xatjcGWsc1ADGsq8TLQp
+eeIdVWJ59AX+i0+EntaL7nsHhPdGuFwxWs1OuCEAO1aiRNVjQA4Whe+bcn25iX0
oaFzB6dnY9PxVv7EVDcX897+vOn3WSBOoLnM1nIJ8wXDqY0J/2XEACyjMvnd5rmR
TFNo7g4HJ0lrWLvcOysVjFPiTTUSBQ0ItK0FoFZqMLZfS343mxJ6DrzwMES0k4Hz
lIF8ugBuztCv8sPyDykZThLxoQeOpapT5/a70nGgqbLjENlMYKqNKG58GcMmKVqJ
e9AcY7PjA6cQ5E37ZO2DgJWYiJcaY1OKPkZ2rIgJBy9J3U/M4nk/bjZvpOALCvqS
/+3llHs7+7hdzKPsqrZiJyd2T3rPM6gCuxW67Ol3Y/+4TEEbN2nBOtKjyeazFBUH
dpg9xycYghEYa9vEJoskMva/jyLR3aLSGY8C3DE+4T8NO0XhHFYcXXLnr1Y4Wgne
FGHO2BVdsQK9w0xg/ihc4BYW44rZSGCFTPZXhZEPfVGW8MgitN/ZTL3ucZn+y/tX
mwRGCEtZs24W6mPM966VRC9a7b2NOoZp4hpvktuHzygSEzYaqlabJUK9DsJ9JcwH
DLCX0LNQ5EQV8A8XCjt5kRzw/cElft8fZXN5akF2CrxYsEtUeFYM6F0j5U94Ujl8
SqsxcJBvLIvrYWdRAXXBW0+2BXLvkMD2M11GOWIrOlNmfdOA5HeHmUSG/Fi5UTUo
jzeyJvp30YyREC2y8UDjRR6ODVyM3e16OkRB/G+ad/LI0uOHqJZ2iQa/Fq9zfJsb
NFnt1haHwqb35d6/k33i+v1s+KZDbAmZQHreP1gPXRXWt2F49NcaEU19UHdG9cNt
MZV56dnbSlTgNRfUusaFbSDUhJulBCKmz4Lbnm2hF/RB8WyTSy43/b6y1Gi+I5ej
IOyUfDRUROmWc3hSSndehK5qXn2/jO8IBEq3vncHHFj09jxrRwPyBWKNoFj1oPQT
CTqi+yxtPoabawtpz8eNm9H3/RiKF/sgzk7tn8B5NkP22a0daDaIM2qzqtl1GI0X
7YO+l8sEEmF6f+TL4QpiIUaXJXKmpumhBzKVxotsJ0eyHfxOE4XxuWM180aic6yT
chZ8VfvT4kOeuU1GQQ8BrCuZk3jt/TH6pP13Jj73r4NAB9ImnTdHVZKG7jTwaxTc
zlvtkJKCniIFmwj3GyaV9Fmmsgz5Tjh5BiHtOHVFZigxoT1uVsuTBC2r2o9QO2LC
Q+cpYBQwygIJdO85WmDCNPa7wqDO7xqUd8ib9GEX9Ombko6Ekx86uOZcRiflSSVz
jvi+frlSHOhG0AySwnSIVcLhg5Jl4cVVuM4WvGPGH3Cl1z/ZIICGi8sEjycSChAF
W/5OfB8JyGAWsmkusDOZQgVOMucEdVA+DosCvJPinqISRprenqull8i11VaAO8YD
Ioqm4ki39EFfuQwQrsLeEDGK0jQEvsE7ZhWOlX5Nxo6qpha+jEgpJUpEgd/dmrez
mWXyB1j9LeAjq5W7WftGWyj3ITUcnZUQqYs67KuTCjiZM+oBZsX8AxhlUB1wjKf6
x5s4Fzcmwm3nbjwqaNZP0EqNUJqpVm+tcJ+NRueeOSvCKVoIy+zt2iJwAUQFDx/y
XntxUQ4XyCnS2XcJGtJz8yJm1MDdObb7S5sfbxm1mEgaHZW6s3F7GQrKxYFR2UQy
AFtEDn3qvdfR9gkgU7T8HcIYO/6KsyIuEKfiFdKM403XbzGzxK9LqZ60wfRr6fwy
zL1Fm3r6z2+/NmTs3LjR7ifMD221LBuiRA8VZSm7fw+7Lqqn5bslt8SrAAorTu29
QOIHa7XrM1Fs7/HW8tC0+57FsNI267xa3FqEDsSP8JNR5bGwki+MyMlt5vfFeb7I
Z8Co5IRDRt9m+ueC8zhesJTc9EaHncLmCj3MbJpMsgNj7tKRXZvzHNjISYdtLdjQ
R9Mrve8P0WQEnGXhBgZCcYYAnb1C6VqlAX4xq8IfBZKcqR96JKOBuJ2c0J3TwCw/
7ZH55mLT3zdw+VzDAPKjkNk31Tp06y7PSHgczUzEvQr7zrIXn0MRzrEAnt++nCBe
iB2OROoUlzvR2v1VEeY7YI95u0VA+f3qYJt8b9V28ruxY3xnK/QUdf3sh1S8zAHJ
D7U5+h5Expd/yZNYHKBHKvjIrOeQnSzSgreUiRGNuK27HmeY2Ke4T0sgdsBtw/Ma
iitomEXH2rHrAITPtcROAPmzUfAqi7CW/cpM/5HcRirxyOSZXVweRuKRZavVwsyw
U2tLTET8p1FcFiFqcdrV+T11bLwAJzS196aPGeFyfwUeoIESpXliGOiX2R5S7uaB
eKIV5sQlN0cmTl9IthlOY4VVmrl0j4Q6E6tqvU/lW8n08Zgs6PN6L0zLlB1FZ6UL
q+6xK2YekixMVA2sMDpBd6KU65MjJHd1LVUsvwne1csj/YiVctNYTm2Yq71m3kK+
JwYn6aZsbfe/UiWq1tx3M6LOyfjD8o5GXagn2oM+ylzSSTysQ4gs2DpVxSFgNo+V
Ldxy3xsYG62oEcqWN/jptVPv218Bcizzh+EtSLKaNIjPRJWhIm5BNe+UbqQGU0Iq
YAjG3z6RHbw/cbFYZGsiUE2E2L6WbEeT0ooikvZAMeYSKcWoNOiUgqQmByb4wc9a
DpiwYMoItQmoqt38CjRZUxQu8cwYdh7xwqt0RXoLf51WNvGxh3cbuu+ZZoNn9YWA
1aTSs4d2FV5eLAUsW+W0VM3ggsRVkqW/liOMull/8i6av27oiVGDtfbyRCrW9lH9
T1V92LU2+js1NP4MD9MlzdXLbT2oQGayogjVvZPd70j8pjZ8wUba+u4EqUyW6CdR
cdIJfJpVj/T4Zn5pr/q59TwXAFC1J9DXlarL/p6gzvCS3isfEagTa0GPD8dQCUMw
2e5FPTJz1/PL9WQzAkKtOdJGqT7LZrC13A+QJ9V3DZpY2tq25j2kp2ycx3mZTUOR
SphFKLVyHJLxuecP+sCTonGkBSxguTXrBPbUsHjyI4/cfpM8kGkxuiuhZcW3uh9S
LHbB5+zdZmv1/c+z/wFZWZ0LBPjncdFQoN0dnPsMXef/JLAvnIQ6gzqHb4ktFt5H
Y0T63Kkvxdh7INb2z1ug88TqrqdThsZ028QK+uJ1/8NNSAWJC4Ny3rApJ6nFFDEd
qzNkDYz2hJg8cFWYXK6dKJEDqt+haXHVsj6bNiBG0tmjrzSi/aUreXW9g+umPvCn
HWNVFUqRj7tv4VMviIpggKW210pfNJzjv75MQxeizvYBqBmJM34Yt4fFcj2gkxw0
vcdJLxOkLQ8rkaMtC/x6aMpQqIafDp8O0bNkW+arjV3KJMNuscExyCTl+APz96mz
hu/yNq3Dwz91bm9HvOTkLR1WWhMlNLnG5ZufRBmn0hNaVACMrPp/bN4Vdlujp417
D25K7quuJeCHL3wCzidvSl8DcBSUYOAYr8b3i8jY3U7lvrR0aacr4B4aHevThGbm
I8jO0docnixMKSr2veygErMLB1LQpKtP8Kp712QKLrXukqyMZE7UNykuQyldXj53
XyRwMKxNmHM0v3XZ9U5BcZCC0p2xePZ6hq0edlORMOkPPQ7IzvHCDZRdYBimA6JU
/eS6DfuBF7xQSgOY315U1GTuJnx6FMGHH+N2k3Z5McglAnesYGKPA0Rsu381qnfa
gsC6ciT/+Z5FaGw1K77F6Bjh0DPSHMSdUgaQYw2s/zCTg2eR8YgCtS2lgqVQUJiu
eXFS6zR4O+BvYCJwFi+0KfOhem3KJAKEJK+GdVlcjPy3NgO388laUXuRr/YS7WnQ
i2zKbywfKcEryhuS0LS8v91A84nZcINs1WqUxzZ5VgwI77UjAVBBUAXWAmaTDikJ
V9M44EO40fXjG+wsxj0aintP4XIC7L4SAKiA1OMj8mkvGGeTumwD+GREVZsFAZrZ
pimTXAN5AbM4PFqENUrZfoYPHHU5jTf7eXN8hihdJ62yM7/3Isv2swysksIzw7Gz
Hu2mlCwZa8J+H8ZKlPlraw7bwr4dnM+/V0pxjByHybFlyqeDv8Qud3phseno54PU
cYLuhi25Xv2FEBomR/OeP9jHpbMsH10zFcFqnsU+NzicVQv6RbU8MHQ51sY1YQbr
OXX9Wp+5K1MavYEbkVYzkn8pKrsi/WF2pGLV004gDk1ew7+Zt8yKK9oPsYuSVaEG
sWo/SVQgIv0eBlgLSsW0wTTSNd4ZCWNXfjv8t2d15plWKrer7On7gwhTlOpiJAmt
UrGnkpWWD6y97uwIrkoQ/Hv5Il/Enty6h3Y+iNHgHqa/nMIyIta1dzLnX9MDf71L
vNeyII2F6liSLRuoc5Wmszb0s2JvnU5NXJITygU8WzHcc1n+mzWGxWIG6oIlixPI
zhsZCLccagaGabswb3LavVMNDK7A5pLBes7j2xmtJSA2XSAx3rnwd00QdT6lMbTb
jJgYAAjtDpUwQVFRSjqUL3iMHHu106OdshoI3UfPT95RTwxIL75Q7s9BKm0DiQS1
tA/ljiNaH1gzzUQfFAPD99Fy5XL3btnHq6d7sm9dhxgkp111LqjjED6N48VFSvsO
6hjv5aSrI2qX4UfMqxZKSERpfiR7m/qc9KQTYo1HRks8IvI0R/dvTNbUvmrXC8CG
8cCaQXHI3jTiH1mJvoc4LL9Ls4RSG01Md39KpTKJfvZ62lVey3zxMSnYg18Yi+9I
S+Rvs5LCPXEs7gkR+yh78tLdUZZsBdnPFFmCfoNfrGInNmM4Bz2xRYX8vbH2iC5D
TFLO6r3PnhSCv6suaytXgKCOBKqfdbnd0bUb3YLOjGHoNsWkmU8kAjKF9ztVfveJ
UQTTs0+01HpxctxZtpqcM7GKszc7Adj5LZsTiHP/EXjzBmAy6kV4ATOyvYiVM0U6
y/DF0ZTfo3YuTb6MqMpSnZR6IATuJQxLTJbzhHApJMih4emHjctxKFU4lGWV+Xd3
Z/ALdPH7E7h8lVvPTb0JWipqKhNEhgkwTXmmhP6H6KPWXz9DBfVmZ4qo8cOODIMt
4yTp3Za7sRBudyEEENx0ic8bZ9js0Yq1saqEDi85E9kcENMd71uQIZeOw8xXViU+
nbPKMVmEBWCA3xa69W1mGxE2OcfO8CiR2pYE6PiZ71jHICMafKywq61e4gsQMebN
IU3jrtzkmJlAgbGM9n/oE/18QgytqXzH8MBokLcZo3OKhQq06E5BBhXYLER7oG2H
WXPRjCRIcUE6WKbWpbmkQFqZkt2ZrSjvkePpD881gRkWj+caNOvb235IApM5x1is
hYRv6A2ZLsjSwYzxXHagNnyWphRMUh82KL86xh7QZWG876s2RZK8dSja4k0OCObT
LcoDYAlKl4YoTU2ygKfU0gEDh107UCv9n7EgksgXqjOkkF79Vgrj7ZyckdyCuosy
VVu1YRI3BEDzrAF9z3OokbFXLh4x3zC33JXe9woyRl2G3AASNH39r4LfUboFuJx3
0jzDF46vtlwAFu1t0A3i2RfuM3W0dkyo6QO0h5ZhEQ8aSRiBXYh3MCOgMt9/U8SB
1a0UFf677zQAkJMTlsLmm9qxISpQSbLhx9beyoedRrS+/icK3IDgt5EnXPOQcZm4
oABTDkTp3EqTQxknju5AOsowURczwN7FaKQBQLMseBNlV4Pdj2Ux0AYbEwZKEnM4
RktnY6VK1PXr3FDqvFAPeERH57WBOGiS8UYdAFgqnQ0Bcpoc1AIdtWSKPMPWgB/s
3HaadbwG0sbfmt53rjr8GvAyrIsZAJRDChUUHmqLp865YERo/zEv3YBnNEjeDtvc
SVDUH07Ud2SqqWRE8FpmTiBuXuOM8AwBlU003S4H2z/KwOt7XOm81emqesuTOns6
1qI33ltFJDZ5eSE/l8Nxt5pjSgUsV3ns6S19etclliCo/Bgz6K3929159oMMgP0m
RO+arVV30gT+A2PTSbavGZh8UQj2SUxmC6961NWeeLyxNGmhpYVIPNAdPa8efbrf
1ySrdiNjF9fpX5EsH6bSDSJuutJFAqvQlmrVj2TDlwvT+HyzR3LjCcT1NbGQZftJ
ic0Lm1XuR0Efz3Sm8EFlZFMdosXQNB48/g/90q5oTj+PHxqZSwNuzzJIl26XFV62
5AtUi2cPORbhrBK5VuTBqIlwxfqdJvJNHugsZUp2jnKiCM/LmnaV53pNZChp5C+e
Fwy+b9VRhenanJi/TtYo2ZXM3xMirKO6Hjv6bit8j6a9MBYkuTDHq+vvIpZdzLJL
KrRrXc10EIeEVBIsBrHa3xOnHQQZiEGm5G3a/s27f7WUiCyQIDj5MV90QTui1ztS
Wld8/Lw4d3BgEls4iXMeeVPWl0SgUJzKa7XufeRwQ+SuDRcc8ssLDcHhIWk3RE+F
szCwjxnAbWLsk0zhQU5B56ieYWVttwcLxMGbHyNsXRVbdlUA8lAOMxXwNajeYasj
IcTJSWFGIEPm5bnthCux9ki9+ryu5tsVdUZPZCJYZaMerAxVa6Er0waTpl6aOVyg
bLElYLWSiptsW37rW1kHl15pvhfbG+Ja8m+XOuXeI8Av7hoBPM7A1pSdLVL0vr2H
y2vUAs+aBnv/dykPcOta3uSei8gB7AMKA6iqCN3+8Kcb5gqPj7TjD35VYWMGKbHr
jwLtKt6tsaN6lhMljJBudSAWdjz7WiyC+Wc04NUlsXC3e8/OwT/VZoI7QyL9IyyB
TU8YPaegjKfkZw+Bx5ofvYFS06g4IjTPSX0euv5ZKvi5n5TAfGnM6rji10Tfv+/p
e26sBZG+DiHU7OcxOv3qtd05U0sAr3Bj0hXwnvAP7OKGy4jLA95f3Lqtz+HWZE+Q
OPg1xeGyP3kKCUc/Rdpa94O/+DD9acAOSGS7288ze6zF66sPiJeQeVPgr23+PfBb
FnxGfSomTLb86l/kcFCZiWqcfFSjr/ss4B+SFZG0G1J7h3RNf2uNi6wR92yLn8kN
+63Qun1B6cHMn0sHfbLvNhKcKR2u/Hcd2TR5JpPQSatTMTLhEZYLoV8GRyOreev9
YeeY4zYe0jM/5opn0HfH4GKz3t+jF0boX4db5Q8ixeUvzuxiQJtdvOGNEiAs2Imj
VXD9RXp/MXnFKCzgF/vesQ5AxWdunw0KVrx/wqMNgM0ehAGTAV1iVwkRrAWzWiGd
cjbqThfF9Z4HcOJzZzeWWREVb579IzHdMmnbvkIlNlGjbBgrTueXFv6UhurpTZ88
hXD7AHCoBxGlxwNYHCUqOF+WECAfI8zQT10GpJWybMeeZrElNptgDlY2ngvsWYR0
UKZKny7gck9NyzrHPvaNbBU/vynGqEjtAF9vGiKjvJ+VWbATxZzyzEpA+Ap3Cv3c
3o5QCoulDZ9vH7AIddRrlcvhGD8tCybYL775r6v4YJuQZ3fxJLaOojcZRYr49sh9
o3GkKAKJiXv/h+RMhsMRERmW+ujVzMf/+AJ6Ba5DZlZTvhFZb7/9xwXiezFEv6Rz
8rv3wafjzWXgMb1+5V2Rgt3oPZHByRgsNWvOLlm8xo0gMuruNAk2EczMhyElvboA
lOcSs8ppQQKf3HwyKRuA3V1W/wS+dH6j7LJeDijtafbDnckpV9vy4rFMUt7L8DIG
NnbLv97Mi+SVOwoRfTJ7d8l+vjhF+snfBuEwYcskVxsit6Xb95P67+QsySItj/N9
T155TfVrVdZLqgdwcJxUzDd2sGErZ19YqlIJpcvTgLAV27+Lb1uz/UfsG8Az9Jkw
9ULWVSnAzGKzOTO7ClSmMary9cAOs5n8j11vvtzvWzWuAwQKobiwM1DRzAhqDrfF
NHEl1uvRGNd6u9yXuncFiltZwKAkmHCju5RcyXwZ+yrmSVaCeFzYw3dXjmIl2dDT
OsWFowgOXazg2FXBst7AvJZaRqNb+ayVoaLfEi8rwSiynU4AsOyVpwPiH6wGcS4G
cN++6Okx5AOADeqeaReAEYSn19XFlOO8dCeY99UditSmAKn3GH+fs2Z4yiHvvuWj
KvSG7/IzRyTCQ3S/hoil0rbkgT1pDy5ldqCSTZmbibQtE34psff8DcoZtTN1TfxX
nT5yvqtmnvxFQkoMGC+n/GHPa9PBE0Mt2ZHgYJxDp70WF20ruswE9hZaGoNLpX1a
0haa5+uGx8ZKpInQRT9Nwi7iyVcRZnJpcLdHRiysjM+WvEwhB+fGD7wVcztzetHR
+Aol7bOhrSjteBEW/P5L6HZJLMBJe+DTf5usN4GPbfe4zvftds7CSe1SGqutHBHw
3t+ztoa0y3boa8oPUzFJMMiuAJUMBYv8bXwMxjUSR7t56+e9e7qgjg2oTr20bkO+
n+o1uSqQ2qN56HTSxpzmM5TQ7rcw1xAxOGgcV0nFlr/MB+TJ7hZ+bUCNw9CUQw/z
Z6RClJMJYO7Zw1RGT1kCeFOPVBGZzMQPG6L3Whmc1Hgn0FWjwDeVB3++QDaw7/lM
dtLfrCiGNByrHWOViHf5Rfw/JshvS0JBQSysa8Gl03eNHDcn1EyssqKVkeE+PPl3
rMKBUYc6oXtjZGdyYXjciGyNVEuTsfgtYF8l3BJ3K+mBnE3Bz6sKr7olIsdg+Thx
ZGzQUZijOzL03oLSX1WzNb0tAqnMPlltFLPC7yP30j8XS8XC+KqokoPT9gIHlmmt
olkXvDIU2Wdk9PH0aHLcoPCeUxpUYYVQqUL6Ji9QNrjZAOoU9gQ1jq9Q+it94OTz
BO9HQNrEgIEV+mJJDGUVkNes0DiHt91qAO3vhb8CLh/dRQNgDJ1H87EuyEiB1JWE
shSVydxJ2GI9wbSaH+NcpLLrg4GR0c69KHNO4UXetgywbsPvBh7RaqrFekK/HqoF
R1OiOY4XVAph9H22hnR1hvyYF3YF0o4Wq+7HjGUMqq+TriprvaobinBaCXzwVDU8
F1DuVzmsO/UqVFZRnPl2ZZifwk+/P7omhY3DAQwP5IKkn0yuvmkebu8HPG2v77q8
FOlA1maYXoEYAArs4ME3ns4p514TvDwWPAdMdnDgym5tKHYKIDNGuUnUsxL0IEhx
+7cdCL68ZjasVMJTFYdFT8UvtdnjXcjAEBtHARvNsBXEnRKvtQaQUeV1bD6lV2j1
6atbQr38eqjinjBHV+KgYUVXEtFPzC+g7zRGit30nUSJLplPx28QOSD2zJshysZu
Mzd3E+E9iKt2skjeWTQ1lppSezqPkg+RdO2Nb5yy8e9sQWIJSxHPoXnfBqwRvIYk
moYzkgAFEOU295mimzIm+PyqYhIS+VtidruLU1Y96uIb0YVWSvoneCHHCE+Flm0p
snsH0eXSPxibk79+Q1lko20mWnSeWundLLlFfzlOUfEAa1vkJqi42rvVhBPrB9IT
u087kmZm6oWotCnywfu9tYwGKNcaugNJDUhthvGStMGcrS58TDYqdMLWMAEdZqjc
YcVtDp5smp+M2+mvTMW8UD15X7Egl/Avb5YixfHt1lVDnuGQTsaxGxg232Lf6HiT
cCVjtXCukWDghWjiO5I2numInK9Y8rA3SAaqaCBfsCma279my21QsAWN5L+0kbxy
fk7fhXhYm+/MXCrDs6ivhbxqOlm7AyaZO6qSKuqBGi3bQRYTBJXFnE1mlFK9D6gq
s8LwaYNb/1LqFaYSn8Xbar3uEfjQzn+GOfMUzxbQnrUkXrHMfdA7FCnXTwNN5ix4
BmtuyclhkihoEuCx5Sk6VcIUgBuG9SKPtRaKue4pRIWAYZeKIgF0umRomGniXAJ/
ShkMBfF57GLFk+tRrkYpiKCQXkLoLKSmGEq1dN/IxNEKHjumUoOWwkFPASiZHOGw
eFO8ZwlsCpRxLH/FmKqnKues/rWD53oIQT1oDhlPvbnghGI9JCVTmOQrAWcEDP1g
3R+eDAJxUgE3WdBBn4JbzZwsnko9Nb8s72IWxLPlY0zjK1DHA0sKcZaQ9LYVFcej
OWZjQ7+LsVn+V5FXudchTOgZywhzgN7sTqzJRSPIsA02I1by1qvEsZF26EF9B2ny
KnqcTEWpHtb3cYQ+K4nTRRUPjqQ9WNgvEownOK4ryP+Z3ppfemV8X99qfqe+CgkA
FGbVwkQtr1N5g7lXTuL0ytCncGENTLr87ekjZlKg3oUpBQln3KailwBejpcGO1r6
qvDSE3C05Wcl1TCvasepvFEJQu/sniSCow865sWQPxKhOJi5VRCkh3J4A2xzN2q5
gZLlf2kCQ8JQxpW82BizH8GPauKfLMifR63lzJuzVgwrR6Z4UIjwaUl7rS8s3Bls
+zVI+2+B25oxUsEwPAg64KPEHjUjdLoYPTq4xfVZ8XwA5xiIuBbYkp3i4uH3big1
p/Apqhf0X/y/4C49le1yL0ZViS8OTsRlQBLlQKoVKu2NU0ixGApgvcTEKT/8Jmoe
ELL9mhUVAx/aX0D/1d6uMiKswYGPxhVosohmxGek3oCTA/AcukTKIReOCEctCZHc
Nh8Wigwe87g06ioOS6KKIW+y5Ic1Of/VGOkzHJSvrO56RosOG5HHerrMUk4s0YvN
Q3DQqktbsVNX4swtOaF1GMKcpKk4pTRcy0gC4XDlGkrg3Ir45jfHbjgYSR1L9P5P
ffVVmxNp4zq3GHNhgpfLwQHgINwJIXIZtnHYutNh1UxvJM6BBJmjtEIng7YrQtFS
2+BVJs7jrpEDSMH6HLaw3oyXFwA4XGg8wO854xcarmh8FJImDL2muchT4890DWyU
EqEfVnjM4S5suOiDcv6czDD4KkaKt5Ds+QaVlfZNf2CoSx3ciDXEHCOqa9I6GOC0
2DjKyqG/owfbK3jJVDiJ6sn+iuFPpahbbGBLJw4AVgtYTdREv25M2lIWawn7knGc
WQodFTstYbuR+jkctSwsfZRCuA5MbBiKpVdE33dKXivnsZpz/NF1mwjtwjGF25+q
nFqGjjP3n9FpLtWlOATOD5xge5U+t1BKAydxEtsqTURPlhd7GiH3tHU6b8rNpvSa
YxttAboQRO4/SP47WhuXDWnGoySbitxIOZJ1zJ1CJCte8xs0mv/mSnQ7Mmf0RHfF
TFu1jTKMEICLpC2skQt8nYgqE5pc0O0drECmef0pFVW1YFm3hjNfancvsFNRnlhm
kMdnAyAvxxeMiOIeLyfmq0Fjp2091mvlGE6nyzrqFaLFCLZG90o1UremDfMVwKzw
yosmUhX48APSd8dbmiQquxEWSAMIulcfhqw6ryqySnAZuKXvqbir6DdjhbCTMQND
aGGS3y7xXqEYsoafOk8UB73oZkWMo1HEvnrB75S5UtJkO4eDBB6mtoa/2Bqb05L4
zprRwqtc/erSo9S3mFwxWOUpYP/be9MDCY+WR8q3ViYjU2a8J/QS+rmT1vEQL/Zy
zPBPOfehcckLt+Drde20oUWo6lWpfYT3nQz+sUBKfdNK58gRaaULi9pHNTqKsaPs
9c87HK8dMpPrvd8oetNpXralnVSraTUhciM4Rjx3n9YvivuqufUQ4HD2Ty/9aI0O
xLCYvrW8OrhI88+JJt/hT9hhQ96f2X9/jCnXxskvVGjA0MsGyiuobjIbDcX0yAZW
oeJZYIkQCJf/NKg2iD94nvH4dlKTyH6YwqZAzug2XpfswLBeSQ2jjKNvIeecbh1e
236+9OrDyZyhHQs7YVSocbI6ookX41Mt5z8NZbMO7JHEVVm6cgDtXNevkZPfzdF6
2ihrgV0LpmpZirsgkRIOc0wxWV7tYUaXZ4WhZajRI87yn5bOmJdaqzkoAe4GaB5/
ikZ8RHy9HE4jH43rUuBon+bDD4Um4+GqVf0xNS1g20eOubFfWiwmyzbazYh/faSd
ee2W5ZoBJId1j4EWsmtLWRXuSM0zikO4PA3ntgEU8o4BvEBNShnt+bQb8jrdXY7a
yCE49MDWaCgSDD/Vc9MRmA8Dq99IntglFVDivORS85rBTrZd89Z8dkCs4tvxSWZo
ATpr0PMHV3ojxr1W0988SvQX9jzAHBJPfDUt6YMIuiO8XRBeuJsDjX574E+wDcxc
BLPFkDRMUT6V5AOelMmoYBeYaZobB71fo/bwTGG4r+6PfOxMSLzwev0HHUKmpQaY
9KMwhZtfkDqZhA4sjq1lguO3XhKF3FV00RU5X1FA6MSWN76reCpgZb5sEwA9p7+w
vFvx17Ln5EjNuXFzDiuAueEZxZIC7FiMU9NWa7SNDhqVslppVLzMhntEL0RpX1sV
UrT5Vjdhe7KPksbbci2KzUtThiWDrBpIUkKQXJOWUunmQea7keBlUGUmCaOGCLIY
/qdqZ7gkT2M3SEo/kOgGe68LzBgPIaZ1HSc1+qt96gbxDMZXuztS9ObDEWxz2Evn
GRlcmNHRzNEpQilgxvyL88uRdiVji/H2P62utdpJOequ3lPqRG05QAcYCCcwYzCU
MpEmM6W2Zd26Dy5ptz85iYjsw08ECm9LlsRTVAoXVifqhUfRZOeDSKejk9dO7wEX
HGOP5F/xeBkEsBi4Uh96/Qvau8/loV6v0CdVVEHnSGFnjSh3IdMO8BACVyvHVTUO
EYFm63tBm6vozNTKPG6Oo5X7Gso33ZmVZ79uZGMlRqedj72rvZju/oG7JSXi5dsh
lNVY4SIs2Xg30Ui1797q0UtEUaTruDDhpkC2RTkSdFAcqdIjDfQUA8JT7kDXmcRW
orH+iXtNVDNhpc9wQ44/5LUZEcjjjqtA2I5gNYYNPbRGWsaxAbqFVYVGtCsa95a+
XHewJH/2ZaZWoFhbuCJdMblxBj5uuZ5+nfTAnI9xbcRNzytkJY4WdzsR0GGnrHl/
2aQwHyJEcHcM/+Vvk/WSPn+4lWset/zq9R//1boBZv38/e7Ub3yLNa/7Lnz585gU
W9BBgM2Yh5L6YHn+jXWCg1JQNBrC00JwHVx43JzZEO0KJKkMpav5P8QKTHN2CnbS
VZrAbHjGIJFEijtO6XwPl6nOvpNkx793de8RhWHmJd9ttJ4jtVQV6wT3qnNfNPhu
IVGOzLAeJjq9qU5dVJtsoazepMYyVAARLFhtv4FSv5PDjskRAxUcte+taDAzgqym
enyMIy8TQvC3Mbi5FhobnKrjnaYkNfeXevcdDTO+st7pAuX5p2CQTBgUm/W78Z4Q
PnRvK8Bdcx3OESso9OuHnMUelViDcw4iJnUBumpw9jZcLvzNf7JWBFQLBnzlsVZI
viMZ07tsryHuJ0JrQmqLCvZgKAK7qqgdaVb6J/v1l8EOmDSfAW5pZLh07PQizNRV
NlvfMLkw0I9+C7TgUHDVaeUALe7D1OzzclBpBqQl0r1+EPNYohAA7kYztYjCjLF8
yHKRSTFqSxn3wSqVYQjzCtzIzqwHzhOxz6RnRzq+NkkasnK8djP3n2mzqpsm3p88
myYtNztNPsDPeKd54llrkuuqzeXODWPcsTUpnZ9pjkEC9wdeDlzdalQdLrZVUA7A
fttZuB3u261Z2p4yywq8sVBR+VIrx2awWZsZ0W8JWa21XTG9i6sYruj4/BDyQhYe
xEtkZp1jD+E/nw+S8aa5z6G+Mu9nVgKcW3hAcNL1tMmStD6QtyanAihCr6qyCAMp
W15/iifwMs6XHD2Q0Z8zaIJWLADlMkmLmh5mcFivp6dnlsKpi01RtGy7VbKhMsut
6fNXVoOA8LTDhTKgt6zWcezZGJT+5ht5ljo9UuURlZhBVTVl4z9/g9VrCwbv4R7j
GqpBRKkAZM7ppIiHjjtFZuThwxBxHhmCWRcR8xReymnNsz8nQyi4eggKOOILaXjY
4Z2u7UPD/THEa1KND0GF943J1l63epd+OQk0deFcHXw=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:33 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G296RDFAw8whPeGnbEsLS+alBp4ruyP1QBU/EDg0Ty8XJi0QOjl6pxf9C5DtMrXf
v40yViNKev/C5ydhY/PX1MCwWpr0zZNFjGnuQbnWKEkL5/H2HKmF7DOAhmOCgwxb
G8uzyAv7oOAjQhMT1dGDYEsY8U1/rSMbxv1Q/vTQJSg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3056)
yZ2+A5KliK3TI9Kx+4yCVx6v99vulXHrnUVxXMpp5W0eApI/HjD41CkfxqoR8e+T
+NqObdVMF/KYWSmLIxTIk7eV2GOzG6DFsWVkhKna+MFQFzzjwxPvBrMRnJ5zkWtI
SGiwIdeRYFSCO8F3wUrQzadHHzaqkVv3bFRBG7S8SZ6qWyyFFPjKS4fRusB70LU7
U3BWB9AFHS4/5LbgM4pShERt0xyQit+FFlQw5ZL8d016EMuA9JXYedvbnj6uEoUZ
p3232RSeI1zEl7J5y20cHdjwB6OoMyuzHYW76XSHPVDLSDT9eP0lwh9E1V2mtn03
Rk3OcUiSO0u+nnG7oqiAAJVvtz5Sh1zvDXQPuWLNzB+7nefV0uOxjdbMYKH6WXMl
toqg1bdF7aSGah9CyQBRw3MrRn/GtnSWWq681cEqICDlXh0356h49zS4y1LFhdy3
ztipXel3ws1q9YwxkS449aMydltRo/fRQq7xuulwkZ0oG53UDydZI6rA7GT6CF9U
f4a4v5doR27OxAluzKbrH9f3rwNPEQchXErc9sOqcY2FrduT0GJTYOsTn0ujz5Nh
SospICR/9F6ZEb1NUh0Y9UcVGQ4DTmfTsHhwdm8Gn3XrTEyrH8Mlnn9f9a/Nwe5H
z7G6GJGb32BYjhee2uWyMMfu6euWo0vbTym8tk1NfyGZNutOdmK4Ln+Uur9xw3cD
2of/c8b/ysbNyQ1FV0A5hiSt3ywhk82ZtNqI9L8CVewemX7g/2hlTothkDP601RN
88MgOcalMtkedixf5VgGO58lHDwIm73KhAv+Lh0x9Lvu0GLFYccDMzP74jPWTPI4
VWBFOBFj8pwSM8t1cpbvZJRggan5j/Jbhm/7belJbPmz2F6EffdqsZOjbSi0VFCE
Nes0/bfY6HisXGMo1jDbk8MA31KZGEN6TnyKctif3ZxwZtuF1KiudzC7BNq7vFrn
ncnfmXu9Fy12TaxbY00qjDGMVgjvVozRtoK5G76/0nQcjFcVnZVBk0NrtJXEaf3A
6yO+SjDopLUsfot3XCbM9iZTvKfbBunkl6smBWL7+VCteRYqKJV0XNw+YeEtn1eg
8QcaF5JtAEV3ZfGKWMmyK0lf91LoalYSNg4KAGCGgAt9EdZ1o/3cxwdDC+XE0b1b
EjCrKJEtvp0Gnw8hGUfDXkl/YHdPiAy0RH+8cdbCJLxrZPi1d+9r8xnIei3Pg++V
0dn4NVhvk4zGOxX2AcR1Qsk3O9OK5gCVly0htYIFk0C4M6WvVqytauhBE+HavbSS
CfDl/gyvQ7J2ujtGQodA1tQUfYNvs2hYrieHgV6H4nKGlTm3qpyX8HC/jZWhMrCb
7iF1TETSAQKQ03F5aGWgoOiJATnTSqdAN31GfHA9zH/Z8w7h8mRTJPOID7MfNHw9
wvIceU9bYp+kLZB6bHC4N8gL8Prd4A+I+skGhDg3cwPEWJH+V/OvMf4k5xVW5jXk
bW1YGCJbIGI5++SC//mqMPVa1Ptsu2Yz8kbvkmZ/i7w+hjjZBzQs+BEh2XdRcR2p
QZC25TKd5UJY6Y70cAe4PgK16/Xfg3uIXohCPR9f3/nrdxFzq5sLVuOli85F/SqS
G+vAdHzwcLXPyEWlkKurKFwaTG4wXwldt8j0yTuZLQlBszT8aFZgCxtEnhDFAPO7
G/nP0bkLFYcJEk8RTUE6TsrKw7W3ye5Zoq2s2uWgztkUDNojyg0+xwtgAd3jYmax
S9VrjSvIhH78Pyso4IcB5duxAzJ7w/NLbAnXqvnkOOvbNmNTPR2SbLWxNKB5ie14
1tinccU5dcNvS+T/fwn0ZudqKe945iesY7JoQ+thFKsqFG3i5KbobwaN6JdtuE4O
336/+2jlkZ3MtD9OWSNwDkv3a1xyGA5J4HpgKRj2dyoGMnWv7W/xNcQiM7oHCUxf
cODi+SBknfzVNdi5m7Hv0D72Nkpsf4kD4a3MUQXuD1n1IhyNkmhOBK7IsMnitSdi
6hM8uTVgNNVNhoZfsr9lvL80gGERATx7MzGWobp6wmjAU6WwqZMp4//pGFP5klYe
+Znxb9q7ckNRTcxjU49MZrB33mqgiiDUArojdh6/+h7Fx6AJvIH4TWcZPew1VO+A
5gf/xFByjqOZALdoxNmr4YPlQl7g6j5NqGsN6fJqtFpYHgaYwPjaqVW+3K3nQTa4
lJ1tLZ7oTT40qDeaLbH5UfWkPIUtatHT9CLePnkGlCBUCztFxZeR/WxTZd8UENZ8
culvAfN9+u9DlVtmFnak0z/VWecWm1pkTYVxgvPSopTvr7meiOT+KULZWZcaGSX3
uw9xKi45J1dJjPwZhJ1dtpoMg1PRrOpWt72bg95McnG0OfRY+7TIy5JJMws++q+M
T2lTOIWp/TXY6+vcTteGnL1PLiYoTGv2Et3OVfvZc8hoTQ7y5dxKojX0J9gYtRzK
6Xvcsu/KzOPV9v6AAoeU/y3ZWtLJXaG7ilHQn9wb8FJK+GrzszkHJ5mzarZD5z7+
nHS94SlD/Wnw1Z0wKjBGbOHtHN31TT3lbZdSRsqrNM0V8tSt0lGsl7KqcY6S7DdD
AMMwuzvzAoAt1hoht9P9DDSu2KvIPunDKNooj0MvK7Nbd2w0wAzarBMKBbW8X+ge
zYGJOciJJCegYITySzF9fSXGBvJkYvfM6cr6s1jVqQJ0DBxd3rsLqCLCBL8CGCld
mBxYLHVGSYEW4KdMRpimeNakhk3DK/6G8Gp5QSKerIPskO/aBGaeo1NLjsx0ldt5
DsWiA8Z/bb5icu6rJYHZThysFxccrH+TPdXIsASzhZQe5YP7T9ApfmGT2FRA+n6i
luV/cq2YLXk4CTIjjNwXjmJ6ZuIyR7wM5VSbPjKOk0X80P5OhI9nxlgzidwoM72D
Ihcl8dLEkhbNKN4oPwqPN5SkfriKI/Z/l91/7jTYcTMdQQrwVIxRXP2xT3J7YAVO
jxB9BDgtVtj7W3GC2rs8vffEo+TvxlJMIliyj3i4Gem6o7WNRu7rth22OLEGN1uz
GNymOcF/mhDwkWT8q1PzMFAstXiBI9wu6Yih7zYTIUuHO2eja8bGUcghgubhoKFR
j3tySJxXU6cZwyuT91FJjic9lJH/LgIuwvxv41eVSvTgFjNGR2vHNilIoDMl/gYA
QvwVuyVtJSL/Som0mHQRLo2N71HgTjG/H6TtJchEqTsvfwW486IdYRDkY0yNPAa6
Xmus0DiKlEBXZ+/mrLikLa4FXar5OpZUJW19Dq9bJKhY06u7sJPzsKnXrNjE4P2m
RSuT12Mg6OSYN8m4uTZzQ9LhsR+QQfmvYk45Qf4Wp7Z+Sf8jSZvLu2rtMpppEM+w
hXdtGSEcnTvMYBk7NaYuiNTvJs5M8pusczisP1Z1B3MWE5ECk2z7MZcbGLwokNr2
NAIQTBAS35w15aqZvWxfLvPlHzlfnO1oza8cUlCaqdpH59+SsCYwBEmR2Q0B8OhK
wxH5h72yM/M8Nj7n4fHgqbPdtz3o4tM/dsMn9VlbcFnaCUH6dfVRl5jK9Ffus0ZG
9cg0UMDTgR+cmVpXQ9Eu4RkTVuQES+2LzTyrJl/gCvQW33kmiRY5pygsJK3xw2Vu
jKXdMNvry19/PyahviNYgw5zjSA1+9BVzxxcIjbBPVB7NIZpia5xZPeZ2pUO2B0j
ryx4hbaCS7X1XWlwPOAuwaiUZZRtwn1PmEnL2cQ3IKEcf49HO+cpR2zqFvRWsHXc
YdY88YyVuhPPBQmh7A5BaeDdkTSifzqoS8bg2Df7nB7FzF19EDR6TxN05CSqZ+1Y
ijixJbrjzdqAYEDEZm9OxTKsRCwlOUu9OpbGJOLLBYBfCD+gOh7NhPpqPds0fj2D
NYJ6CPqdwfMOu8JA9Sxv0pqUnWAzuY+oK44HGxFa4j4o91u2/0FMisEvTeSATswU
9B+bgdM3xEmQNqVF3GbUnqnF9s6ax3dwRtk2JB7GAg2OC2IiYx0YX3Ds5R8SSxQi
ERFsYGj0u8QU4oA5mMaRKDECr+1iuB8IiY9oEftFfS+aSZ6oE7UNH102RrOE3bVh
mji0X39jkgZ9Yh7fxHhZcsR0k8Hu+MXDcuU6iADKpXM=
`pragma protect end_protected

// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ZedPukJmJgNmmlIaj2mhpKfjKnMRu3gJZ3UmvRs6QRNqCDHJuuUVwMahcWP8S8s04ZGJXOAMWGmp
mdubpXvDSH2ooVJ0WoemRRaBNdOONVy80+6Um+r/Yzem+F49fwgcJRYExAOHUMOkBDlbx/4zIh9t
KIZJr4dxNFRUcTkhHpaEMEL1sWGmbK7f9gwdsw9K1x5UgQjdZlCLcgT8EKabTZsDcNenoic0LNTy
MGo0HsX/PAiMsV1P/md0gdWg6dfaKgssjZJBQicPH9pikkWkDFs9n98Bck8GMFtiDuQr6BT8G6FI
dTYh53KiY01PTMO0OcFfKoYpKHMA9j6C5GKMsw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ftbDSQ6U6/mFH88qruX6H6+FE50SAaxWMjrQrNCgzFNA8f/+9sneDLLk2vCloQcgIehw8+Ks6IHG
4iexXeaR6bVRf493/kBjqd6eGBs2EPSH4auW/I+FINbFUIPq7R1xTK21TvNEs6b+WBq9fbPXlquc
VYFllO7A2m4Zt5YOzB1emGVs6rxFCEsJEy/A3G1yDqh/QXzVZT81Gf+WwymdurXHOqqlUTLCewmh
P+zzLC2NAEkqC2DX6oZ0CzajL4PUPy6aO1W8WPz/flAc6djRAYfW7ebPGtBJDPmUfATixWZ/B29N
ecOL/ZCIMybqV8IV+p49Y70AY0ChYpqmLbahfnoyZyP5j00Gcw1vPnfRShbIdtwSui82VtGx005x
kjqJz6W5nUYSbSsUYvaCqLJ22E+OUXLfHu9G+NWOBNU6HGFs93+SGXswqeMn8/NBrTaenCJ1+deK
As9qnWMc01M444n3xxhFZRb7SbXg9EZkBg/5zOE+eaWejG1fAZzWS/oyGMaM0mLDPd5r3r/834UI
Q8EfshFrke9VDw4NxSKgBjcSKLVzICVPebv8MW5t27qhA7nQRa1VZcp6JCdpeaC7hP7AbbpHco3i
xSI4XSpqkldhx9MdLsl5Yx69MAX6lL5M4cbYswiex2Jhj5ZU76vQRKIf2EBfO0FYfHbvmTOXmeA4
cxiV14rzYiZKECy9O5J2L55+5FbJS3Wh2kz8K2OJzBm2BUp20IrgEh7pv703MRUFLt3XkqVgX/sF
JDLQECdVoxaaYvRQUNjT3qv1oJkoLHP5pm2AuWfs7b5rvQpMqy4R4qA1oDe2UfM+OnivsSKu5WOY
7lL0QfkAWoHl5qOkH1jefzoN3i73Q9WCAGd80uUTFFJQXycl8tgcqtqvuNnDaIPKJ7+qG/ab0PbB
KU/7g9lZZLInkliqNNyPp2f1ELHM8Uwt6wwDuBAN3pd2uaqSSS596byeDg/0jvYuNCinpozOTtvv
NlW3SgIorNB1CkmIAOYjEk/mTkMMN56qKJaGdZg5Nrn5LyR6MeiMZ2yXBMVliT5Nwd8PdEO6JGhz
IfWe494wLHBSH32GdpNTo3p0iXiVlFf/CkBXoG+jnPbO6rWnyj6JJVs7FLR02s4WpSvLdA75CtRx
7YiSCUbrQyapSplZrVrw/wL2blUDFtDFVFsjIt7tKZ7FEkcoa/ZAA+vBEPmfY2LtgQc9e/Y13Gga
WOgzrHV7X9MaAsEc7k1MA2KvS7uRiH/wOifBJ6KWph3q+ve66HeW7/HO1Sk8NjOHnFC3ya5vVbJM
bzokpe91Ocbe9T3p0BEAgFQFh/003zRnHZipWDPFF3fBwP/GQwIjLRhi+HaxSmWyzEA918XjabXB
HJq8bOClZ0l0CyVpNUe8Hanm1hAQEMuwBcBwub5XeYbh6l8Jv38ZudpAxvKftJaXRuQEAp7c50h8
xiRjZMAWa2g7DQihLxz3GL3T633lxOFEIU9/WUjAHkTDA3hKGtawN6SiYryNbAVBRifgyG62OGNe
GWUazWujgwufbjyU/DIgHphMSvNAPD3zHd07RixXGKUHBNUrc56kZ+gl/uhnd1DSW0Ub+UUULs1V
j3m1uLTlpD9xBvKVr2hHG9AeMdzOP17bTg/CiHVd/L0kATbbpdmAjpShVLBJl3wfjOSnMFohHJqM
Hz5jh/GnrMGW8lyRbV4peO6bZYnctI4ko9C5WFSnyx16j7IPxCm7RB4zLvH+E/zz+V8epcPtDOc2
rIrWUiMLi/+Q0O7HvtFi0vZcHLNnQrZ4cXQm/Sl+kLMY+hxPd5U/jlhsPJcJf8E5aCuijCtMmLxp
pU+N48E34Nuxsn+Co4SmaqqEe2yTnJ2odiNK0MwPZ/LxWd29UbaetXPLXP1rcFpQ103rNor84tA9
hP68+SW7Z4YIhuPfZLgnEdmAWVIzX8n/K8oK/DXHfZ1j+jthsZLvojTrosMNoyXUCX7NMWIV9Zm3
BpTx2oV90pSgITS4defTwsfubuXheCDl/UZGEumjudGiejxEHhJ09ogTD+c6BhiHbSw8alr7X84D
e/VyPcmSiL1KfVcsu9TDX6EbAK4xgxmpnKtjImnmQjiOP200Psb+eLGd+Dke0WC6futFUWFFr3F4
v2vXatkXtS3hF20ozv23zhJjUSmsGscThBb4nVyFbYme5otlt4gYZsVd7CPsS8zNZikzKwTlnVBs
AKApDjnxNrSpy4XjfMYF0sdMxah4Sd6MtFW3V4JhzXHxFW6uJ1oZuqbd+pZKU2hK+Xy5H5SuOjBX
0CS2wrY7eKyEL6WC4NzU5qGl5toEzzZ3OIv37t+d0g7Tv1TlXmSBTzILm90c8THg0lg9YL7VW855
G41S3KVgUwJUUDLwnkB/9Z92l+DkNgaBvbTkdl1c/5u/xzpSdKad/im/61ylxoymjqbEMr0Q8m3P
IU66DfMe8P4wOesWRGyuSaqJvwL103teNfeSx4vBgAFBSQO4pD+3bmKxjiMAp8kYWglmWcGR7+YO
qCWR1EySS3EinQ9X1Z+6LQtlVznBBaAlOc5OtH3DL3dDa7sjnUuackHvbQsNRGulOXgYWa5M4yIJ
1UYzCKVtzoAjK0342iIzmI1tUiI2UXFDYi+HYViYKm3XjHLdgwjyjAP56J0DjfM/9HFg554PJm//
t57EjenX/dLEFSAGw73OBQrUkDfcz4cfDU5XXmQZ8D/N2Mb2OOQyJReSyOO5iRWo37pa7WlWqchy
IphHgQjbpolbiYKVIQwaMFyzn4uFu5p8UZAqHEd1YzGFbq3TqtHyuigkyRILEt2bXRL3PooGZCmR
sxGnmPpipvPUDAoXDsbqVpR2cGumUUSZe1/NEMzTnd5lZuovRGPb6rhTYurSjIs9MXKwI7zq7mdK
VEDFuKV6b0jC/WzKLKUUx+65r6+PTRq1wA5UaVT/nQ1cdgq1T6roq+VVtrTcrw/o4cZuxRaD4buj
j2bQJRwoia/RKvMMpTfJC/0sLQyKmGBvDqpjgR6mW8PSTVYUb/lH/QdgH4pxMi7dhSzBImRvCfGS
B8HcBXUyPoY8ShKKseATnWI0ij6MbBgHdOtbrqptcN9Q7ygNn7ZDrN2TVdbH37cbMqQ6S6Jbv+SP
0CSedvKzC/GBxcexq2Rilx6rO5DuQ7J0PMjxV1Ctt1gr5r4BcxtZXXDipRkiggPtc/KrpftHc3CF
VAa9vr7bDEM2TUjlud0IuuRp/0PASh48vCwNf+ok9kq8zW2PFy91fTwRVx/QMHPDqtuDbTvwx3o/
u3fXNrqTJgztObmdNcu6wA6udIJiQol40IamrOJQFJ6Vxp1e/wtMD3bKEWABe4WL86AeTVsKZ06J
YDc/65RBscz5NMpv4lMzjAW0o8hgr4wDo4Lq4OYA/3RMD7buhwezXDCLb/xOPUDeFE2UmI2C7GG+
+c54512Q/qJyQgBFFstJxmKvircxUqrpdW8Zpe/e/kMjkqbVsSN68g/bS+9my7pthCfc2jBADXZY
Dov1P3LoRDoMkkKXZbq0Xbtw60cz4a76PMeruzwYciScAilYb3EVMowfl/Vh/QoemBwmbavZvE5/
YL7ovXcjZHAAJtvZOLNdjV+6KaaoztyK49ScEdyd2La9We3CsOwGZ1qrhVX2CLFnFxQjTTj1rKdr
tLwWWQ+ZzLbHbHLiejRA7hy9va9QVGVBkJWiWeuKXS1kgU9h7afoVO3Vu5LEPzkFrSKZ7XQFsrtq
iKxn4CQPMW36HlidWTIdm43SP2bMja9j+g/wWByQWMd+3cE3jI/mxAE/rth2zS7kURkGYHLWculc
7GVBa5C5Yyz1nvSxcgjfVyTyd06hqqHhhg384EULC7E26i4uP9Q4WqGbN8ksEauo1wyquJEbRyVx
u78MxNgRgjNdBc7l5LLojE2fFKOHxrh0Jd5mfOJQN4Pu9vP2R0ORdDEzaUK/kiSNOyQurNQ0BJM0
nkMRdZGTRbVw7biFYsP5lXMO8tpnQpik3GhhkHlfJZeNbmkGSRb+q1lZHy3MflDThVZTPWnaJEy1
K6jAytExIwtIS+3HQjR9A1coNgUVf4lPCUn923Uz7XoUpg/i5xfa3khL38G/9+J6mSdpNDpvC0rh
IiE0RHB6TgUk6fLvCRoKP9mkX08cO+SKE4YqqmNS7TUbOH6Fq7VXGMs1SZlIQmK+UTTHkWkwUuHE
YxH89Oqtb84d4ZWA+XlP6NBE2UwiF35+4HDIBKLSnhmLYHenynbpuIs+X/Bf0BAgv4vIixHq/SlH
CZ8f3Lm4QGfydxpJtIssMl/0b+/seKj8LrpELBug4dVwXSpc+Rvg2XG5i0ViCFqPkk8pFdE4N0kO
kdLoQF3ZUugmM9vB78qfC8Iwp/Zv1Y9/yzrtGk9aXZCVfxR8XkQIhhapMyOmDu0Sqn3sWpMqUPa8
B7oQofE0KUsnpon2fAqFqPjcd98kyNJEIM7fZgaqElvH1UtLYnKO+yT59pjuaLDE3KopF84wLj4h
G0yCTQmhs2TQAiUB039oMvJSGaH32BcxTcz92sIt9jd+EkZ1nJEuHpx+Yp0AxDz2MLWDA+Z4aZAM
NVfBbBxytYe+mRfqnwEFxevS+fElYa9xcKVvQ7jR+HSEsuLBIXZhPWxVltYe7CnhPP3BH86KcVVs
t3rqF0AdrUZnGh23At2TIehHGJ+xBu81HL/DyObwdaKVAxM5J6UUX9kOO3F9+JHHMAH7pvdQ3lAY
d9ExpH4tqLiEmcAXougWDmmlGEgIcpLKe9H5PKTep16sCSHVOQgcUwrW/edyVO9Umb/bquvu50B4
bmANdP+cz5dYPQ9MZ+Dle5SDsKJaJbCENd/CYbCNZQ5fh2gA2zL1+ihyBANNtvKITteAYeRIkjpJ
vhyVNbe6fXZD77bEdBh7UTkV8WmHbXguNIws/pV3rGYmFICxTqQqlK0KlwFE3BHhRagl2iUhTTXE
NIYvFKfNU6SEFJDhAFvPcvfRgTw1LyNCv0FaHW+VROEbKcYfhv7CpCHPYcNJjmMPak65E/saOT4C
YzWDchaQ4t40JFxAMnpXlhrkUiBjfy8V4avfwzjsyrDAl9JHIjVeQnRzbB9SXeFj4kKzQFe4418l
EpwyD0bYzhw3r3e/unkaD0rlou1NM8D+0w3+PWcMH4DxXBFNY0b/Gl8U+9bS6JasI3YNild8vbpl
GqVGbxsh7dxOvSLIyu0zpCoqBZyRB0ZPVUrV82DMU0oq1u1DcbILuQdHsGEHobtKE4lhbmhx0ebd
NXsgeIpT9cEgW6IoLYxoF02JD1xMpqRYnHl8ZOKFBXepomOhmkOFlEb9Za7fUsd2YocM1fibqkj/
aCU38VCpDKr1VX+PSDYmOSMSlwES/uLyTcCRPPHBO2K7jyiCh7hNod8gGLFm2QyLictgweBg/zKO
RdMNtvGAALVzH3rnKtgumt79YX0N1S1Nj6oTdfBPa8qTh74fQl0oivGE0Mh9CuC3qXmFoxOoY9ID
9CFa5JytKAtM4wZ7vEe6gE6jDznzeJ+bJy7Jwad/t/jmFQDWQCdrLITkmor01kPPPIg98cXDtX7O
f1pNcghtoSa2R6RtscgNyZnSSiOqsAs28JuD/ONmqzSuySICmpdAqClsVXsw6m7LMPx1OqiJSiXg
KkN0rf1nSCuHr11nuv0LqXuFaRCus5z75pUnNQNmwsvZ8KFvfilgKmK+xsHkp8tgBeLJD9y20fwQ
I4J+EJVTCkU71nL6xnkNDrncCdFkuehjEL+WBXQP/RLdCrIwDlKxRf9XtwLg8SUYrDeLoD8CWhmx
o2PPLrW0C7PwEfMDpKpdkrgvgp94McSUzzPOKj040TyH0EFH+vsHV89TbjDUzBem+OidXt7VPoCh
cwTyVL2BHlWLevjgJIWWs7c6956St15jxFM7Fh2QZYucVygezT7SgkGEORiFItlzfoCyVd3ePyFf
QDOA2N9TTXuHqKx0GbHTxL7G/y7Fc1ug3gTqmzC2nqgby+cgVEDn2mmccxLKm9rxH7FNbnezq+1H
Wf9ORpvBGMvsOt+1tk5dT8DI8KNtxQmxry1TXcP9y6b8iMpUxzebbExGjbLYFyXSaJssERo9pgcc
neWQxbSBybPIOFcucFVWfLJ4jiGXfPgOj3v3P65A1p90AQmgd13JibiwRw0hSgr5dEE50gHClh8j
QWyi6F37HuE2T8rjL5F9F8mC9xrXWOXBhiq8V0PcXgg9xjeWGoglshWVjF4+8vLK0Hdc1UTMFyLX
AYh6pP8Psy/GU3/TsR4Q0TdavP/Um+HZUdK/KxebEKUqrVMU8wjvJuxbjLp/8Ixn54VyTsTjR8uM
crrIljkXFTTdJ5t7QW/xACjRqESF0jLS5VueUS4RTWv9doW1kcbBfI3ik0ZQf665Idfgbo/co1SA
2CzIIvMAoP9fEN173l49Hg8v04TTRo7RQk5HhORXdelzgdlEeK42WyXL7DZIQ6KcbOkOrzkQcqsF
hwpbq6+9/4a3pCfcsi/Agkqj4JVf0l6EYUwTLBya1kX82eiRO4EL2a20vlY77+xYqq9DGPa2vPCu
HFwWE6nMQH7rqxF1aZG/adHAc/kh8H3VY47a1lfoWBDR6qBz2oJ0lryqoHrbHafu7QhweON7145X
jXwjgjmjN2jltrms+IPeR7d6eN5FhJh5dem2pnnTfx815bc/ZNGpSrho5OVZPTL2WboQeLtYTdBq
5AFxDN+Nla5JIxzF+JiLWLY1ce0G6w/uxPkuQz+PWO5eA0LJuX/6MwSZUuB5BIOTNM75moAnkXGn
hV9wzZcgCmIVNIUrGckw9KH0muLEyYxUDmyJMF66kwWNJb0ySIhnWeyfvU05h2xKYe6wDMtfw7SL
AJ9Ac6rYRuc4XP97rIgO64Ge8d7UlwAunggrTZKrHTcUZ3m1a/7y6Yt751sJaeEi4xK/0bWvsdC/
c1XJuUBug3Q4MZZ+cleaPnr8P40QwEG+QyuVG2VB/ms0GS6cCr/N28lXqZv7kU8/zu0GrKNY0TMa
PQxfsON+zOtE2k8DhIRlQ+KCLwjDz8Im8OlERzPFV7PbMOj7xbI4h2L9y6llmmK2WU7VgSOTyXAz
2fuEEp9E3xrU9VCH9ips2rg+2SBgHQ6tkax0z7IV7imITCYOwMq2vfhJ3LhifuMJYIi0rzn7ztRb
qZfi5Iklh66BEKp303BRrX/w1wV1lhzCOnQ0eeHES9PJoMhnej71d8hPj5S5vsp4bOJW9lWJRs1e
I68U5d6St4wyLxSpvjD0hyd30j9e5e0i/5BQNvRsT38yFr6TUwtXUDLlzM0AOzfO92Pb/1ikTwVQ
UgP9MC+DluZxmtELVykJllcZD0lWvRVR165+ufBn2BVbjqwZ+evUJgzBZkJ+vvmjZPxH0yN9G5dP
/PVI5kSfQf/cJ6NYPzBvE241vZm2wsgd1I1umV4p5kaZu8IlA+ETV23J9elg5vOvmF1qMmj3lXAy
9ANpY28ygbfmepPa6546EB5U2Yg9YaiVp46LcrZkuH/Jp1Vp9WjPCM/+SPTkeYp4A4C5USPptM/J
/Z2jyQsGD1nEJVxwVLnJUguLHsLcMA5fkYWxnE1m2aayXtI55UsdVk04WzuLjYnn13txoPHq4/j9
Jb3T42GrsrLNR2UKcPVx0ibmiBCFnM/remx66dKPLv/DBqVIHayTJfR35Vy3Xzbwj7idSdFwLCnT
ooUPMoC0kJ+RIWYNvT1GuL1nYgbPsDiDDnTQtJsp3mqBEygLdIz+K6WqNyotsSanqueKruNg24TL
00JO5ZgCGTA8GofwO7ivOp+tt0Ktxr26Sycy8+Nr5ta34D0hsPREyVrinCgEsjyw+HC4Lb7j4QaR
ekMqRrdecQF//dZQ3abyu5WSwN0ZnZympZa21QFD0txbRdgs/ZlE7czZTqkROMIl7Khl9qETI88G
igmwC/zRakQUxzp8fd2aox8wCPQcNogYX6FyTeyvhe7dEldv4Ypwn5zpgc6moTzVp2ahHssWk7kX
TBdqcVW9lwnsdoLS2Gjvcxzwo+UxMZ21anLzyk3OUPPTOiIwmHvrebKaCejPI8SDvSbi/4JO8yjl
wBjMdt1vJYrEkOdlOEOu9nTrzwJtkaw8Ks79/iVFemmfFF8bI0amK1KEyFWNi6H/r72+BQ8lzwUE
IDmLg8yuqsHRV+EQjB06d32eQa+6Ys5dK0VPP0Q6y48ubiPhx25ILj2j7a5iqNlUedQ481fL50C2
JZAedQ3PgKghJzSHtcx/68ju1vwtnwQI1OXMbXWgVicyVern+SxuF7UtCaLcZK3Dx8LWahGT12rY
u/SAsTP6Ig4Xb3FoGzEYE+XdpDlUyuY1wPY8klltxFA8r8FER749AHtjswkfI8v/wi/hy6Au6SI0
3gVKsW7p5eZ/06BmR3xp5h2uFhNoVSnnoDXSoGWBrGKwCXkhSBox99iFfG7IdPN+ihR6SBWhXlYe
UrBdzN3OUZpIUgjY8GcjSxn7gkvbYkHV/Mt09RvPBp+9ZsC16llXTF/z2ICjLSO5IXa349zRAl4a
WDg0Q3SXTp1FMigM78Ns7V3M7NYBc9Y+h5EhuUiu3F2iH8TgPb5478yfI+qv7f1zGsv0BQoSYYd5
tTe+OQiY/TkHBMOVvzKiuQj7F1R0q9d9XyJso5PlpzmZnVUnZacyHWbj+iwf90MBlaSuIbt2rqZO
90UzadZ0P0o1mIxc2l/PRg9YIBS2slREeXePymOSNVvEqvOxy35XpI/DIF8nJemsygM/tLPYsM7I
yjk9izayHsVAkH31UU8f5Spx0/Vm5UYbUh3WucgtWt0xmYl0/3yMkc7a6UQy/qVVGO+g0X/H/lJa
IVI5+gLFUAjcXHsmBypYaE0skIcgFDCt5ZJ1sb8AOi5WUlbV9T64+F2JwpZVT26TDmTPB4hA+aR9
030qZhCsicSFGUoh86wqdKRaYuqNWXw/SjGPk0X664AB3hW159QACLMbh4d5P+b6muRGXQrk7W9o
bjrD2/NMNut8/tvNO3+XYjr9kctUvezXNubx/sx7xjX+DGrj3Slb1WRsIF2PZpPQJlH2MhgjXb9B
bciGfsxg1d9JgVVwvP3DeviZMia+tReGDHMMgBofq965kaImvoGm6T7QOVKQ4yQpPxugN0OPiPOK
5ngMB3u85n/cCHzru+nxvqpg2v5nU1BFh0PC+5NBGlFDRlmA5Qz4hepppfXpN4SPckkYV2AOQ3na
Koj2KudBNZc4fwWmRuydmY0V0P2Sg9lAV2RK/9QqmHdswak0X/0i/V6HZ5bHTzhFKEap3PhlH1eb
jQuuESp3wnFT+fdoPIk3Oba5DLsD30pP4M+ic8I3h+I17z6qLxuYGTlAqEZpr1RXuEME2cyMRLVu
Km29Hddq2uXWAde3YkWmPk7MbBNztzfDQJZ6n6mQ8N1bTF/G1+9MaqF8zEgqOs5FqRpohCHxTJdd
THCxOK8QpYcj1LQFjBxastxJCGympi1y9ac0y/IefcwQiTggQloihk8j3ZjWNsuAr4vzlaoArWR2
by6okbxGcQEQILbQs41ENbb4OgaKM3N5xvTIwpKRBR2lBpVVoX2Fp5ixsHusLxpvAcbfhQ0GSMVZ
HcA2kmCB6sjPR7q+cC8YVKZXlk8XwkH7VvQ9AL7np3NWd7ackpRyp9v77tjiLAa17TprNgC9wWP2
H/AHBFjMA9w96KjklUgJk3Cs+hFaM/+geFC8Xxo8SawTppH6HoHqEKjunPKUWyu6x3lnVfIkWpfE
o6cx718JycfVzJ0PHpAwL5g3riWf+B6y51J/SCJjMj1F1HHY035P1214y+f6QKr8c0JeFfLGfLVS
fUdnZqcvWbBmHsFzbyF9/CLj+ghvLZ3fsZ2Ls2V0o52LqHT0lKNXojpfwoR0eUmvAy7KYt0uDHvQ
wwKn91887Bh+MbgQXJWicZgq/OpJ/81d6Y5ico5ZDE3aF+7nRKlb2jvfszAMEbqYvx3sUAmZ9cHc
BqKTFMoYJ/wFIuhWfP6AtbVy/CYTm9lvtqp5kmXZBcaO2TujITdXXqh7Yzzx+5XBI1rirrNMxdIM
y0iQ+5Nauo2FceWfFGNtLkmutvZyooZHj+/xOdINzt1yQkV+uuKU8TVG34GeOZIPLR5EVahQJvuw
qyro7GYjACcHkzaPTL0NgvAhDAecGRkHEnv/itfghqsAgU2q6sJwMAsl7LPRHkHgisKt33aSh0xP
SgCU34fmsh56ooJ91YZt51JBuG0Tch8X+1Qi+74O3w/kTg0tgvrrSUSKOYsJDx4An1hCfQIBAkZK
Qs6RSeI/+KaWov5OHVTij8t0V1rFTowIpCZVeYrchqTl28TuvbzCITKu1F40j2SWdj0ECEEz5Xzf
FRDXwOMRyX/3r0tkd+nwi3Xn2g4TC0bF6IkFhj9tcsY0fj9PNrQ/Q1aryEoe5yBivd05GER9sH8L
UWBjRK77IMdCUk1sxe/aXfmdIajhfvAIHsMgfUvxJRRFxLd8mLUey2yfEegDB+UIITPs9ovelocy
D56AbbcgaposRoPuwV+rhagDfHQlNvbXRAo+MiK7ac/mTqjXHO6gMqdQ0OmjQ12Cb/zX6w19159T
5wyjw89cJT1S6ZMc8McGI9a2IgbYc0YDQQmMZ65curp36U+i40wP4p7zKrO7sxf73tjkaJzWXHN1
hvKRW0DhYHZuNBs0NJbraoMjKJ6AY+8Av2E6C/oV+b5j2vHyULtAUSt/XuOXEXgrrUuSL92y8hXI
w2i25WmZIJRkGh82hrIYvRZffdbAgLTLT3VQvHC+00rDjVUg5TyKX3YZC20Bt4ZNLdPS/EWDCJvJ
UbQjVi6ON8m99c4k/gfqpB1iCSWheGQL3JvvuGj5kTQsyjWMKZiUXDoyvIDvSDaoQR9uYdB8x87U
fs2czd1jUSO+smhb/tzRqv1C20II9d5mCOKfH/awu//ischScDMJlGPsVmHFmNUsA6iB7iH0gK5r
QMwAReXxEEPJniqDqDEVaii9C2da2l68OT4Iwi5KYajFuVgn1Jp7i91s+9jKoQaitia5dvH8nRLu
/lFtr+LM+VsgtnZ8HF7mj0RFolKK880erqTERmM1PVjcLfK9dWY7lAtbhwkp1Ox9CcUDl2LnK+10
FNfZf+rR8lyM+IOAr5ZOFfDlVemtuytukZtbWy2YlDCb6Ae4r55oTwDvyM3W6s7hWik976zbzH11
B7ZVda1PvpJo1A1PYnWs/efXzbjIwCKGDXnxs2Z59RVXoN+NcZQ1KUyQVwE/BTjGd+gQT7o2dYaJ
JZIw9i3im8ggcDnTQxj+i3BL/QvJ+xmkoY+jpKe6zzUQBD+DkezTYv6myGIlNWiaY9zp4343qEL2
BaXXEygvdHSguVnA2ubB929Gn4wI6NqZJfQjQFOl7jY/XKM/AcezHitw226XoWO3RF9Hr5Ckti1A
zXtmLGNzdU5AFBdlfY9h2RYRyBUmiRpMFWTHWg6lzLyc8hHP3XN2so8yahPRRn2SzkOA4KMG0V0w
3aPDpghj8ZauxmZaSRF4Jk1wGQm96tBdJOyMZvFWBfsg+J8UVmh53aPOfGc+P5jiDmalMmq314xg
gL/7fFwoWN6ABjMHToTZFVAw42z0LnOrkLa5ZyjNMfkz/fNceAi8RnTgixnrrdoHhhT5dP9PvphL
m2MqdNTpOGQDJq32xJMwV4Ur+fzejHf3lF1NY1l+/A/J5ho3lyXmRfLLxgaep9CnrdeaBtMMK+tL
pxCF1TixOyTSV+AiM9gGNhjua6JLihGVgm927ItpAE6hcgtLjvp+n3Ur6FfSSvDPnp0kqNr/bI7p
n+6vfPcHMgZ2LZHyURVNEJvSragOwIrSQum0tsmFezYEjBtFpCr3Au4dc2Xqnnq5C5+di+Jkqd9w
erP6N/YKAxy7LJrBoITr9grm9mRB/x1tRwSc8HtNbPyyJIveFt2ZAEvimirC1zBoZHBgT7qSon/K
b41LLtBz1zpxs7pznHWvITBWgS0IQcq1bAqLBAhIHGvbAa2UR0R56OJx1ZbP8cA72ag45Wm6wi5p
5RECRXcT4GWvoIQSv1qO3VoK3op7HELzekqCluveQVV72BPKmhsjgPWoJ2Mir4UvBoqs0zM5AKzP
ZkGOqh8aD7xh2+2iVaqes+yleih4LjrWozAdO/P7OqFcDaQ8FqIJNjSD+3LbvR6XOsBodCEPK2ef
Wbp2uG1XAI0ufJW9ms2zDyxDH6+UIF5+vYnzd+JjZ02sclwRWjPmVOzglT7OWUYiH84MXRVJD37N
KCaQq1Mr7ekr/u5+1+pCaSlwoYb/tr4j6SfsTpaXs7SuRcB4j5zEJicLSurQhz2CNCMm2uZ9+QG2
JT5BechekqYcWHQ7gI2KagoUEmlslTNkNyFDWi2o1xFu0oGdMXugyRaPr4dl6PaU77nQjE12UpP1
ZyGZW9hI8H8TvH3wa0kkSNdMqoGyMyyyKIAbkml3u9q96biD2LCgyva+2vpVcZ1yajkrSPg=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:28 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VKTPOwpMTBKvhS9EyRta4cHwvY2Uu6QBts1Jd5MVx3qGrx3IWEoqqrLTwvwWYbcc
i3kqfEW106slOs8VoK3upJ79hd6F6GoEg3P+uNYkK2dD3Z3EekNm9Bm0PJkCZhZY
20iOQ3KMWuxFtg6OqYpunh7Z3EPSEfL+88bNuiWT5v4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33840)
M2zUIzyUZDbUuo1y8rOz3v9oOM/EewMCLSUyR97UOVFKA5Llf8Na178zut62hh5S
XPdlsZctR4RQPfhbPsCCcFLFPrj7yhxVPBA9ZVmyyr/fIMl3lIDVVG7MHtNA/s66
bfO3Q2xNw/I2Cxct65RBNRmcTmyPsLfVqDWOoD1j2qRh8pXgKWMcLLONbIvqmHzB
+28+uZiNr+ngNX2BZ4YA0FdUF2wmjuZW7e8GGIFiL68IkFbdmjCnFq5CtxPVBJpn
PqtGfVJr/mORyy7qJmC8xxK9/gv5lu/As3OWI4McyheauHsjO3TPC+f+hDDQ33LO
XGOJLqtHT/2Zl+cATe33Om7VliqPX8cTq7RSER4v05L8vK1CdVkRzX7Jbl7IrU/e
9Se/h9nqPCaErNjdB/SkZ+tsIjl0bSThfy0VqZS5AtnNuXYSaZE0SJQttoZkNOT2
9EkoM0MbC3x3TkOXfUyz58DiOeWJPtzi9sxfFKISdfOZQQ53qYd9woAGB7rHie5g
nNqGTINDUVYTvuIT3nl3GM/cdtZUwU8dwnaQ302VkuTJDNhyfYc2gafC6Gaa5/qV
CGmealul9VuhjDGyKma07S3NiSBpts+YeJGVuvEqUQopWtwO0Zg2J8gZbwfgvmzV
PI4mNQpckrqD7m/RlHgDRQwdq28ab70y4ZNgvrauJ2vW4uzjJRWmzMWs1JcLqp72
Eysxx0Ixp1RKkYyBazPnOy9vOXZFsIhV0/K2rebjXycaAACpGH7TfFfVGCOsllpZ
egamFP2DLDH59ahuxHIEHH0VPNC6b+W+RuRT8DSxkUoPFiCV8fyyz1dr4d3aKusO
FFwcZ/QHiX+LwNiKcLbBgJhHUapSDinyY8MgbIEOZgIEoZobd4ntKt/jzr7h/90f
/IZ/K9EZSglRkMJEafh3bG5PGyhNlUzYmqqN6ufhmlRhvMivRhMoN0jD7b5JKIVw
dTirOLJ5Pf1kvAKCyAlKbhAiZhbWfLjHH3CMhrCq/nLDC8Ohze7YtpFDTxt0OUBl
Nd8HljPESevFOrkadai5tch78ojYN5kshkAaiv8wjknAvkUomBMyrQcLNFZI7Cmb
ml0PVHQYfI2ooi57OkbN+7EuFi8BFY7B+szWiVaaXg2VhipGxlFsmyD8SPm8BKZn
wKQAJsOVpoVO36gX49KAL7ec1PAHiMCWbR0pdmY5C6PdPcLTAQwTIN+CbgSFkY9J
aNPJAgSBgJeZ26UW7V6fV/cEEch7x7WwlKIhRlnQJ11nii4tp6ndUXfZpH0gscFY
eEPGtUtazxQmfW42bYAH6NeEki6aLBXiqC8DzA1Tex9YJP8lK+WSqz2l2+jxi+bD
UXWiG9/0Ph65p5zT8MgyW0X6WMyPqhxwa+wzodYcB4wECCW/NNtw5sgnoqaHLkMF
F8QEXaOqdbjA5ZP9P/PArjyTQRnzAGEnF0c+6cSKjRJ1eNlnHevLXmwIO0WJzXm5
djvqK0Me2yH5UNFtKEp1cjr/L0ccolp3osh22zO5wTHDXnKdwMumLuj1NJxTQwe4
eiiHA2kDuPJWJ2tem0w6YNdGdbv1oDqhzy1fnfOCK/ERA8tJyKJ61djg9Nh43eR7
QVfqts6hL0yMoWavzhVQIGCF7ppCyQfDDp+IyzxWMP9KxnubzIA+EkOgAdQqI81s
TIPSobONyR0Qdck9mMnSdb4Jh9nw5bp3vXRZq5dlJaq/6yb9LYbayuZudrlsMS+/
SkRhubZwU6cJY4gO4T4S/HTNoU4qKkDk+3DAwTeHG6N8UoFgP+XTWkonMSrik97d
00GJktHuCWdWf1zJ3oYEuMfzrl1vmCZb8DtHy6WJzRZFHuiKPVV8gUBP9DJt8bQ+
oPfmpuuHzV7yKSW0Ms/lJ0mc8zWXKb/a3uLYIjQP9Dm5ythCST2V2ZJx+iglICIb
Qu6obHjLlRTLE8HiafyTYwIN4qtg+FeuWP8oq64MBwbFnLdMEOy4IWtaK8yhR0G1
4ow9+zh1aIoCFNbtlamIo4+0n2Bdql3/Jf0fVUSYE84ME881pIEy2DGxklDKwitX
ye7JZk1kEvSZ1dgW/LE6m5lrblnHbt+VctHnsO+zqT/EAFpo4rOORAiemfM80rC4
MdcrzTjvAVeOA4Z7mkZVhqg3fGQenMkVFIoOddWySPCSLfj6pUHhFVELpP3pBxD9
dUV/bikUceXvYjD0YbcvWGq87wjym3FWdNEQMxj8WY3sUXuf5bhm/gKKHeYPVOT1
IwKWSHhZhuY0LJ7p2AaXspak2sXCpzYPe5X0CO12MHPK0FsWrW0En7N+GEyp6B8k
Iaw3gRWx53/UQRQ1G753B6IDi3mUWvCjEe9Tgh9tvBFVmOOpHJWq9r7yFIm+baTX
Gk4eocjr3FufQMl5O+COXjZqoQbN6fG68b/ToV37thtjRRz0V18wveRt1fTECKSf
qYke/0DtKIG1StCfUO1oUnBOVtJ//2sm4zq5TvmrRjrnw2DE4vVLIoB3hfVHAjOX
Rapg+KkeeUUHbaUiQtL6LaYYcme8N9ZFk78P2HRRyj2Hh/lJK/bW7phIH9OXNipn
JrP7J9sicqjLSYXDtpLNaq8xlUc1GYRuyCKd4wlY641/jF5G/qYAe9pkxLRsPyII
+5xw346brs9w/QDEP9mkMtJoc6SafdShVNH/+8XKPwcK2DgOXQXIvA1B8r+7jMHE
u726rX2qgJJIYUMA+ug90eVYe+LHl/K6KgFDBCmxHupz6366/4vc6mKUU1sxqh19
NrCfnPQ7dyvmledyf0DaZgrkTwFGoec2YbS9LwUOnfZ9ude121PedR2fyVTJHQcI
sQ+lmCU9NbDLiKIYWPAKs9nXX20zZQnWwFowWOd/rS4N2nD/O6/CAH0xJgoJa9hq
yjiDzQVKVoS5UCuUQ7u8lH3T5ANex2HFEMRzykC2gSmShpMIgJhmAaQhUMs+01oA
fHnEe73INGQ8TMahONujFQMy+P/Vw9uorzQYizdpDLVE2mdAL4/T3Rnsp3znkhv9
U6wJSU6Cn+N93VqSo4rfV7ogG+L7fm3L2RiCiNpKDE6Xw2a3GaRHmNO+cW+BSi9+
Bgr0+z8SjdfGs5mX5LV2bAjt6OWnnsZoWIp10YKN1DyQFhTzoxrWBkiFIMCZ6zNj
erjy8rjUTzFUl7iZ9MK4pEwhkx6JMWmW4MzxZBhxcx6C+ki9m1B6Gq89ZVY8yuv3
28loWFX1G3IG3S5T3q7obumTITzdWBraSJRkedcHv3CyA6mYrGfQUpprlshq9XmJ
/ws2pBng9iMHvE30t5c3djNVuLYLsPc8b9CZ/8/MACke23Tfe/5Kctvh86YJFNH9
jEK0tYCOE/OFwtxGbx48ubDt4qgMSHrDg3KDlD09HIP26rCiHGfOkdi/DNo13i/R
nTGv9pWktuaNlZ36ockhAVKkMLiLAia8gw84p7ilI79w0bODux3P3uv9x3sEiVoF
baGJTvemM+pveMzUaal1YvotwzVv/gdVPJLwp3CX2ohC+G+wK8xbalT7A59Dcov4
erevCtKdOMM6MARM7T4eIQZKyeIdXE3LP541qm8bOtbzXImVSDASd8mo9F4gwl/H
2AN1QYqVY5tAk9g5XpkQ+CjaG2Zi9/kll14VNsvQOB8Xa539yBXM0W04FTM8OS7H
bJl97Bzg5/4U43843fZCe8b45kheL7MZ53VcEjjQMfHBDd+VQGmLAn4MzGG3iojg
8zuwCdXPbWkCST5N9ThVHilknaT/sTxV/MJOXnSLPM0Dd7+rKmtxqjgGRQVgM8CQ
fmM+DUu5IOnFV59jfzPxNM8zgyqbJ1OOO0WA48X3CjOgF493UzERSj1uzmUjdhGq
WM6FXrzIuBhlHGwNGmR/HhOZWXOLapLNEsdHhUB5JU3OsPfv9Z5AIk7zdRAy48dH
eGOqvPPQYxcgGsKNhDmCq6QuCRwByRl3iU0k+xb4KI7Virf2LbZ6yHvYa7pTr1LO
5WbJJ7Z74mKzaXkKgV03PGzYyRkHPLWcmUPkibZSdl08wiD2eeW+V8PRGLB+rHn/
lNDWQcSiC8LEulNWmhjP8EK00V/XgR5qBFBHlyLHOLCLuEN1IMPQ1+HxDGE+kFLA
BMVD0IRSEZNufn8bM6MX8TGymdjpad1pEVsCTPpWfSNzSPzJNM+wHngGDKPoMWGZ
++aLKGa7G10HnXNFNQaVpZF1gZ+l0MXj2gzccxroniFxxtJCPzCcB2qZlxsYdC/G
QxUDpH6OZhrNw0YDMFEiyo3jiPJz1HIYsk0kK8jup3W2tRWc47yth7tn/3Lk7LXR
Ypz8ZNzerLL0xdDxpOtZrzogu8+hKLVIYmnMcr88F5nHkqJYASHVfTw78RSWk1oS
buPFFYd4WtV8g1jTU016wARDZo67nJmtKDk4U+za6cWxIhDhbfjgyOp97NmeaqNn
9VdYYhGuOnxZERqlxfpQ6f3SdzD+IXuBIP1hsCl8NhoYQ0MehMTmxhm1eF8CZbAN
pIMQJQGGKB4rVmr27bIQxaC2n7az/qFrdb5apbiPM0MNLDM7jwFOeUg+hmH21QfI
dHwBWEaiOzpZE2zQU82hD1eQcjMOKn+ggedVfMyHBQ2YmVtSiuXV1+Z8ys6OJmHs
hxkogPDyig1OYRaZtR7pyhqY9PeBWgOpw6au6AbfPW52IEBGMI+FPdXnyfo3tZoj
bowF1F2HUiUTQTSk37BtmRHl7Mqf9Hk4gk0hGrY8h8qS0q0jIvYCQtYqcRA3JXqm
5wOu3/1Uy+n/Fdt/RqgxPZ3YJW9VJhbpNbADe/7B8Jug0qtwqKSfVa+Dz0V1ELF2
AupMrTZS/s3W7Jo846KHBmWP+0AKl70Pbdf7go+swQxliKT+Jvwmsp22wikknPLt
KSiu/L366AUgnsJL/Z29txf4xgk7EdaxYWxOf6dUCk5Pzr+k2pYBAdkjAsnmWC+k
WkXVSS3JPy6Ri5B/aDbku7oXhTK+4UUde9Yo/OA3/Pdoi0AJD0XxqUIuVJpYaEfX
BHjyCGnfHWwI8hWwBOCtdg73eOrF6uTQm8Ht8F2UZ8suKLhrLJsGR6rdDx1v/3zj
Ean9fwx/g/h00rhsTiW0qf6kvVbg3g3hEkZobLr46q7b5rZuBALHUVhPktN9B3Ke
sdGUUe7Agb3gCmBZR+NaNz6n1FXRpyKirMgOqJRjkrDTU5L+/HyNOokjTKJLrwv8
ZbIfym7a/wXpCCQPH6Ylxybw5HYbzncxqqNNtm1TknZs7nEvKhmqh8hOYw29EgrZ
mJKmFgWLHWOAKrKsRlc5bN6CVOv8iZ2mOn1y0IM5BOK2m+VhVzmbBIVq3Un1GNiq
mOZLKuNujocYgfCg5jHHfz/iYUE6RmWkYY9csOjF5FelYbbYsj49q9ql51mPkVXZ
AKi3Z7J1IpzPoM67B9em4MMniHU2Bd+buv4RVYx/TkFdOEZp+9aL9W6QlTiv6qbY
P9asZzbha4sea/aey1+F4qcN6/G6y/YA6/QQ1ERgX2u8exWEaIamnw+2gTLoz2lh
AdUUI6uHAW8ojlqtRW4xWfaN8bSB3Sawvwk6Jg+QTt982f199AoCgc5IqTCh7TBr
VgeeaHWcPKeQtGi1oFF0Ytp/0Ekl1YNx42XjpS4QsYZrLLMs2154hJMPhOll6N2v
hhLwUk5+3bBD/BmSOLhad+4ZHaanebx5309ngaBVS/J5VE63FYJBKAEXHsMGK6km
UfmGFUFuUJncDmAutSmPtQaIPx2AnbhYLYc4rKufV/J/4eGEKOr1YkA/K0kyP5+C
5VhBSYp8MSAFNehfu021jdJlm919FvnsEgwnhe+FB+Gtb/rVTDgCAK6CkXQATvj5
lrsAPNxX6xERDtqe1QwPI0acqWgzXt5xk1BqQRc/xwWlngL0yEskBvrftc8vrXq0
RjCjJAhuPQJXlik369isEdiE8rRaBp4JJfarAKr08t665CfEi20tCR/UJ77MkePx
TLqSrWkvdWFAflctC66PUKrQtSmKVyChIQ+wjMiKNdgrlzj5FcBD43IBwoxpr+Y6
7JG4+tAeWYZwS8n6bD7cYbbmAdQNmMVEoNllhVDX2Yo8Bo1egmkx8F8CoUc6i72w
rAgoppoZNg9QjAvm+N3F5X/Zd+vsi1l0USUNQyj4p/dSU7g6l/EG8Ph6PXvEWHvx
DHHE/MtQwHZZfqJo2L4d0f5913ImHIUdynLnVUC5+0CRUR3i1KqZ5UFmOa7aOCD/
+lrc/kseq+nWu7yqmTV5/pHmSPLnYHCnLC78V+I1Xg+1b5yvGvBS20kjbm74cX1a
wS85MDkacngmEMxyqsJGyFOweTFgPkUlMymBuzfpqLiwdVX49iPK7o3Ho8dlyuWw
y3cMZ7qcE+B3jULvKpqGPPFXONZxxnrdl+pdIznlQb94G0PUPZFuq2m/E7Lgg+g5
PVOI2xWt8ugaHWF/Ey2BrXQ9nJoRSZmw/4gI7h2DAVc8qPkPy+HQ/qVwfpM069yS
sKjH9qjfZS7LGT1GC9I845equ5WX4+oMLab1OYgFi8qM+/aCLDG/nmIdFk6hVr6o
n/78RTaVfhKfYNvQcMDWro0KB5hDu276Il3V+MXvGQ0V7eaqpbNViksga0iYn9xC
wUYEhJ//c4KPx1mXz3PERHw4t5s9egRvo41PxWnebuP3pfDpc3BU15WEmMNo47z2
emRx3C743PuY5lyjH9Od4+d7R3c0huygUAz0vqhXC9AyOv2DAH7RzUYcACXlY3O0
HDJiQFAYBmIHRBplrEsv0N9Ycpjc20qczGCbWw8n2MIEcMOnyBji/eDxI65bESVn
0Y9FzNA/Y7d4Pl8UA0k4ZtZc8Q0Tp6oWlu+jTaKUWUjd2yueRvrE2SImmorQgnrK
18G1yN20J9rQNDtgO5WkQTq/MvygtKqx1zKgxS38k693LiaUlcDNReiwB6R9egzd
qBbTkuG11H1kwdnUL5tjNdyG8wbXpR9vAmTBlp5YhaN/HQ1JCB8dhZJO3FKuerbr
wkXAnYXpNtaaRjoSVdKWuEjWEemJQxI/7StpiC4FVfHDvZ1agIePZ0KNc82Y3TlA
pyE73ULQnsnyDqi/9qCrWs7+vN9mM9/qa0S+viavL6qysSzd/Lzx8XlCNf9hB7tw
v0qGfZ8Z1Tbs33JNivD+oSX2m3kX0N3PjZURNqairF+ZCupLwrL6Vsgdas/XD9Wz
EgReDgQbb+Xr9PSuSyhip9aIqz0JSAVMWIY2/xNCTzkvCLL67bHOWhwf4Opwhr3k
Tm7OOu00CkSWobRvEBEkZU6E4KSWUGfNHIEdrcXDXoBbpS/aGC5bV04r48O6YwP3
fr8bjlMOoCJcty3p7/sd/3QH594jA1NIAKGphkRltoD5RIW9GOE6GNePVAzcWjY8
R7bt9xGDYAwhwo9LlVmQA0PkCFv6KI2SWmFvaekbs7goq0FztKiQEJZNFyAxLXoR
rfpBvgnnYmsgJC2R6IpO9f7Y1VUBpD2ZUjzZi9headK8fdPbpVujA1ztqlMV4Um+
LalBLuRZyO+ge2KmBhUDYi86KiFFdYyaHyPNXY9xxu5+1uPfaBCz9hRZsnj06rOI
QUSs2CaWiWZtpjPdgFIXbw/0U5eLTQUEB463wez+mj/s4oxNSzqcOP9IuodlZDRi
rkuCpn2Qj6KuAMM/mZBpnHR8d0of13nN4gHaNi9ZhBY6ppkVqYXTKozJOwFUfg19
op9h/fTEwCvLlNremphHxirxsQkaTCy99yqnjUzftYVLgYC9F4HHDgI2KUUZkUQl
7JtT7eX5jYkCzk7VPD1lPmxtjepdclokpjmnmAfxqy5O83mwh0No+UxSkmvbqJuu
yxn0Zw9tgY4HOYH6MuM2JEcPJcYNdDv60Boo1aiAaXzJhsJOYmyqurfXDuxjc7eR
kZ1PSUiDCbKpSybsCdWjEKN6KBqw4OhLZzCuIKIabFXO07QIDuyzwZtaDDFlH/Jq
WhRL5MSW76G0H+P6oLK2h9gaqrQWe+zDggoK3xtRUYzww8L7nybyhxY7av0OW/N9
iZdfZF97EAgfY/2EiqqYfiM5ybCjDxkK3HMdaA2ky7napHb004NF8awtdNgtxiQi
oVRdHDqbrtJBEdwNGkPEHhHTaSUzZaWaS54McHtPZona851yJpGWpRt7MX8okjA/
0eR6Pa1tsAIMTkkZ3xypLE+yObPMhunJpEYO8SCq+zEtHPyTISudnprXd0EyCWuz
b15WajGv0M/aOH/ujSfAk0QFJ8+NO/D0mB70N655l0PF1PAvhW6ZFdJTUIiwd3v7
/DY/Ejq/y6tSuUci3i2AZ7ACvyZXiwkGhXirNeJ91XqpfJ3XkIOpeTab/Vyt1mCw
znO1aAFlfeLPZGnQpPxoqISabfsJWd7tZ0F+D+hSaW8Fm6VvCrQjwLTdSG+WpHr2
FC/5uQiA3nD2303QcJal492FaSXLqVOUddE7VaHggOMeWblBTucOE+f7FJLdZJW3
fOmuYIq6yatU76WQvdZHcq18UBFILAcWSPsK6Dys5Nt+Z/SvdyhVN3gIGOG24yUk
82+goCGTkNXR+4eMqFqiqYY+AsqiASRjDij/G0WVc6ejT8JSpoMJX+qrDf0RRBsh
BIrbP5yZ14SykCL9rkpdrNcewuzhP0u9A1k7kMoAF4AMlGZZ5pba5L07QEPA/Icc
T/O8R5msgua3KXr+ztFcMgMVJEovEqaqC9coaDA6uGkZ5FhgexloBgpv25ZlSezC
UBjLRVU5XOiabLCtpzlfwe5Gc5nwR7s4nQbcs87LK+lFYMmfpSptyFiIuyceHSKm
wqzRDvIiKgoLIibzkPsPGTsj33hPdkVD0yyOq5VljiLczhFXPp48/Y4IY+srDk0L
F3eI5chTPPS7e/A+pFT05ltCnjkNWiUuLCHirWwvDOGIc696VRo9/U1Zg88XegYB
3ifHHzLK7XCSrqGHN9+XrMolNjz5BrxqRrtsV/ADwJcOLI8axVKfcOUiM9tLguTU
cUcFl9qJBC9Id2RHVvdnEP/9OFimTlMVrbRGmgK/RhyKCyEzXB3jGf7VxA48heNw
oFBpPujZMAzEPKQwePCTbN3kc/p1vO0T1/azzfnn5Erea/kNnIypr5t1OFmaNVxa
CEpY2jeh8mZiIfmT35X9EANwNoSjHoEEQ04M69P6LLZgxa4BFfVSM/G3l25RBQVZ
DFwfWghDu1zTCcXKqcHnmcTf07PzfAu6K7eFENwk4VdH85B+H9OJAZN9+2QGp4kF
op8pcyWLA+6cjESOQWed2QPySwnSefPBU80e6cZraL4wzPE0ksFKSetvia7VMze7
SWw3zNnBnzZbJdKjwKW++cKoQAksleKpHqAlFYpvsqxEWQZWhsJcvLYmadCnPVCU
5QoOGhyrh/zhzem5VEnaLxYHkJOy8drShddkf6smuny96wZnFq+foLweLN0qD136
jVEkSXVwdjIdraD3LzbT0r7J7RECwYsrVPXygiLYtROlmtqQAo+22k67NbikwdIW
xHUvzZpnzXyxW58DXXH+b/T4Vv+B3d1JoDIV+6aspVa2gQTTo7BF6MXvqNUcSTR8
XC6Ag+T8ty2CAC5+D9SdluRZtOTeyHLUZKxdugWfa5cnnbTpOaXL7hWIM0KL8KAe
aFtM8FQiC+p7sgcyjCZvQLoaBdIfouVHy0M9q5qjzVEZ2DQfNlDz9N/0PqsL5wjW
EIYUzFhH7eSYfamHrNf2FYN8pa3W5RXkI/AKDlYs171RTuNdT27/CSkjv6crCwvj
TAN+GcOYhokICKQNQV07auTBLlQi2SEXA15ZjGiPui5dGsID9F+PqCkeicTOLRyo
SDcKfAlO0P3QgzpbWQh64X6MnTM4kObLG/jflI+/noL9FFHpnxuDpftZw2ALF4CH
GRn+TOk2cAcRxbpve98+Ffk6UphRIuq8e/FUosejfuAC1hYBFEfk7cPLmbYCp9V6
Lv+cS/PeBl/p98ZGQja1pEIoZS89oRGLx+FiMQ1stmFREFdVWKl3sl+h8+773sXX
0e1BQeKkuVzFoYZN1qUbbA5HZV4ameeTglRU6HAn73FgP1ZesUFD4zEFLt4bb5hy
lC6e6TKPHzyMwpkUaoHRnxCpNWbzxCn8nYMTdkYAEDKMWaPDIptIW7VNcweInUws
u6fsVH3ZXnKQFFKVK3nOXt1ZzxoaC6byxQOkd4eN5VF/WYYWx11hAuIrHUKwly18
NPfyUWEEmr6BozRlAyxHi+sekr5NH3pycM/CsEGrIdK2ukm+iMSw7BeAVWQ9eXYI
YflvEHtDffeWyPR0yXBnIXz/BmwHZ4qGum62vixbWnSdioSAvGRdT9EB7rgoI6LY
brfZkm5WuK5YML8FMDTva5MWkSpPWwtMmdAfE5VRwi5e7hdhGeiUvtfPhzoucul3
Bea7nmGr0p3MiW0mL+9l66/0R/5lPLg5lHre7LFKZDs3dIEiJdvj3bznxHi9EuSL
etABbEYuQ/osJmi1uEktSa1X2g73MAg5eMa5e1BOi7NpYF0T14/WXuJ1VM79RMfS
9E4oyr/L6B8zvNQ3L4lz2Dz2tp+FgemMnSadA9H5jNGtxfPWrgahbJ5bEokGoaq1
nVPUfWPKfCkrCzhYh5Xp5m+L+rEwV1UnfvZrXaxQI6lEgNWUiSpnrU6FSGG8rZZf
KYmja3cP9HO/8YhoaoEr8NykK5N+Nw4aqgvhvwsmukqpUHkxPDrsYUiedbmGOTBt
zmsr3Qu6f5+ETdtflyVukM7USAQf7X3J1tLNCyWIGf5trVEJB2k9jRR8I9itZ7Ry
uoaMzDlKgoVd4ol9NCdBjypxOhM4MfP4T7lBJzfuuUBJvwa8X1B05Yq26//GpsLs
qFIyldNLp3YjAOXrjdUT15q1SUL6oiKrQ4MKRNMkHT9RnGXICnm39XELRpjYvf9z
l09BopPEIVMg2mTMi4kL6TzQSFGAT0MGPHNRSv7E1Wb3oWCg2ltkWn2dmVWEKAd9
Ww0Wm7NX20NsJ3sQBC2G9yl4/49EqZYW8Jvs5Gp37yJHpU0RPOWms4JELdDjhHT/
kJXcuY3bf4IfXEBqhGIwkaL5kfM3s+NAlGYGEAb1DRSkob+0/yvIgCE+e5zc6uR5
dpw/2mKQMJfmxgcBwdHeri3HIbu5TSwa55cRnkLLUyB4FT8FJYH/Tt86blir+2Pv
Te8IQtA0g95Iy/wOndI/hBvM0xUtnWIx53i82T8ENF6kXjvCoFR+P7HAAFlCTMnS
OR0kFPP4Dwh3/y/5gqWBrozs/CfKTsPl/roY2pv9FEkuYR/9JEZ0Dap5mI+AIB2v
6wkduhVL55bhXgndg2hn29Uspeepij19/YYaxX0QnXx2LBcYFFmSznvYY7IEr08N
WVllapwfFqGz2mtmgaaF/MxZne2iWh8aotRgxEjxsIK+tFsD1heaenhYJbuETrrV
fn/rCrlxGCdAjvgK4/25xkJw+ed3myqVDhB0Fm/heFurmXcn13WO4STInO5crb8/
sn4Dih/JqkSjOMEGQTf1+uUbp1UR69hhMxmxDDUhp5asHxZC+juddxRG4sjuKE7d
8GVqXjF6Mi7y/U9ZDJnYEDjtLL6G7NN8rvFHJRQP/LS3QH+L+kabiyO/As6GdHEm
726gpXtIO7OjR+778LebPrM5QWaMZVLkgjPYZ4WHlzWYtBfu8hHuiFhWgdxoQU/e
7u4lm+Gl7SFzoxMNtZqhEGDMIycl1SHBLyLQ4YeVw8YBNumCsb57v0loprwKr/AI
3dWnlXO2IXUHSHik4BbST/md0zXDNoL3jtugftf5KV/MAqi30ys5G12hrZ4FoUzT
qzXrLuFORpS4Y5cR/y5ulMlE7m3MotDP5DZXhcayGd/9F9W8VqR162J3l54sG+Rr
nkYA2Xl6HOruB9dgijBxwy0g+TBxrz+9deSzQgNxkgqs9KLqcaa1Go1nirPqlFDq
LonK6kQUAOwdKUtKwj8Nbe/dUycqMHAbGvPndy6chiOv7obPdxfAqM4q79eopMLW
Ofpz5RiN/VZ0RQzrBe8m8tQpMlaK4iN0UKkOKQWI+ohSb/dcfkuYLi0aVwEvyvkc
lecuD7vF7cHkidQNFI9fIEvWV1j0HuTqTZ8JHbYuqHTkfGL1dUfzj86Gucgke9sL
McH6yVzZZCL0QayVG4QB/llLvpb4NLqtS8ZMlyT7aJs9+6TdOXtoDA5xFX8vBe3/
/HgDHYzTzqP2GGSxkeuHHV4qZ8I5frzc4N51hbof1JDhdifI9s4/PIHR0Tq9SwH9
bFYS9NNEAZ5bJvyhxt6IRtZd7A9sSpLQaCVIfUjRu/6/qTvw++HRVU3eSXZ3x8zW
LFPKao6IK6L1zTydwdkBZa8faEWkO3evBRJ00RotTHPzrF98ZXNdNQ7nU7/3XEyV
CJi2Ympb/X+M9zn/p65V5beEaxJ8Vd9q7Ku/CtvlKgI0FulihB1Rlf+w5hwSlE30
t0vX4hAen/OVKHL+PX0rnyWMFXRUOf1lm+ESqb3oJdvwsD5XrN3NKk7dpfDydYs+
uYHtunOGdugphb6tZn+r3CpHrskaq510uSFDZsiCso04pVBFASAlxQmgU/UXlP/I
rdEsWTQdE8EAsgqdOKN8zeNHNykIvuh/WJX+f4eFlJ4dxZIsfA1eZhVOmV5897g4
Po7ev2ezp85dg1n7IepwpGd0rbcDUgAaPf8uRsW+3yOvwI0ueOJgHv3u3x3X1UKU
8uA/iRFI/eBcKK0TG+tsosKVUbDPQYhDTT3oCcmckZ2lQO6MaE2RaqV0CgSMxrd5
WQdXp4oRp2zM0yyEwX1xW7e/WpsxwQcM5JIUGW3okaHYYfxvpHUL/gZPqlkTvk5b
EdcGWtmkWm7dDJ56OSQbZLuvWfJohzN1o/DGNG4W/l+hVC2syrDzr054Pp8OShrj
iVjgMxkbajZ56kahIrGNvNEjkA6Wo7t445yByQ6O2S7ulQ8ScHZDuEZHgG0Z5dzs
Rb+DL0bCX6eYUr1Rd5VkCs1b0z5ZQOMQHGpXl0acalDdPSF35x6Py2KLW+kVlVjt
Gi+nMm44bYarq+4qJ3fht2PlX2aVdN8A9DYfbNdo0pyeuuzMknlNSD0GSy+qz5Mz
0sHguVRN13K/GCW21l7BXkHhcM8RJ0Mj3pPgfVVa+iJ9douwl+oMAMdkutlhPq3M
O0J3I7bytdPLs8t+3jl3LU8RWvZGuH8rrhD6ieXqcRUofDInvM1TeNjVw0smabiF
iQeE6QBpm47Y+xJIjiUM9i/TYnKk6F41yPRsza4FsD8vroljTqXmDY+qPtGYE0Tw
memB7YSs9esoBY3hYe+eP5HUBaA1LEunMnK4c3pXIVTqx2BMoYd+gxT6Z0xAh7Y3
GYG1OPfXvoZzPb2zv3iVNwV5WPcJUnF6ZxzwQuG23Lar+dnPT6esPNTI2t9EMM0g
6U0RbhnJZb1TiKeWSIX75zPSfeIy5zNSUAHWHjsosHv0kN65Aqo/rV1E9LYCOB/e
V2wPQJxkcbTLO+b1tSM6nBfDDE83VWPBqRJ8aooh054bdqyPfSPc4pCkEFsznx6h
t1dTVirrKzgX8+cgAeFAnNLKEX/2C+HOliD1Isi9eYOLjTWM9FWOPclDrvhyn9E9
MSH3nT3unaaF2HwcCb8T7ctHOnq8DwnFj6XhGyhMy1ksjW1r7yBu+mPtOqs0WmZL
B/m2y1Lcwh2EnvgKC1BC+2O4dEj7NWMEGUGBfGjs3Bf1XgznelMNbkZQTKybRmUv
Xl0o54Wkxa65MzW9/7obWedA5IVBHoFvLQB+m3WHNbFAYPV1kl+VTCg1f3R02U0D
zFwwaKFLr4qyL2y1a3PCMaR5EHKt4js5Pr14VPuQ9mg+sCxd0yiP08ouJROtzvB8
dgr92Jimmwd++2V+nYfLsNMqs2CY16Qzq0Tw9xC3pmSgEX+HyuqaGQgx/wqakHm9
xl1Ywedpuw775D8ilu/HX1Vj/+2UsRWPBoqo1UQnUGs/ATCFu2k6MNNhbM0dmeiA
LSG/fgFZjUQojnt4FUhEbQ9kno8fOAfcIoEHlNIG+4psFcI/c8QEMFcLBgD26Z27
KA2inSZO3P+RwG5utroahLimOAdan/Xl03vVkdEC4FD2Ur9LtgA3Hl2AXUq3yZAT
NpfoBhOys+xNCtRmcjCzJY6oRnlf0rGeyFtnYXl1DDGUXJ17+94ZiLWsoY57e+ck
KoysNLDk5GXl/tClWzIQ9Fvhbj6j7P05Miu2BDbYysuIZWfU79Ea8WyD0SHUoyfa
cC6hn1dqB5KZ2++2wyNRtt0ewtYVMl8+AygzzO85TT5+TingeQjGZ7E+DnMetgF9
mDVeJiQ6Pukcn6XAgerTLdd6T55zmsCJtdBMKqXIvXmmhti/GVgAwD5ie0l3TWxh
7x4Q1fsPNfd8FF7GwZ+KzX87Q/uI30NII+42Qs9nNnyOJ5Mrm/ZNu6p9QpdjMrK6
M/DpzcWwRYx+oHwP+71ONa20o4ADLm/xiSf5mYhnyJqGnCAgJCaMvlUVAWydgbXf
7IiCNuzWg+hAIvXn3eibiHQsH49lV+yRzReiWQyWlKSfFkLlD99f/f2ktbpFsMSL
IQ8cem/9pMsK18vaTan3llcE1cRgmaGHZEUTGcy3iA/ELLO9gYyUYHBrlNvzWb8r
b0QcXfdZzjI0476kWpIOJJPETd7l7YkhER63aWcb70Na0qYyAyGbsz6GMgw0Qf9l
bGrzZFVDrxsdMBQMsb+bAhB9UHwghFxSn4OMW6M7Px+Tq/FrKGTlu8RGKIXST5VI
yMgbmClfzd3WdCAxGHXZ/dHRXNsPj/4VvO4cbifiKnjZlpM8er4mIKyukhS/lEl8
cOxIEqeDZ/5rkaYFkMvmStE6s0fDhUyhetBYCd376yVGtXE9K+C+7QQsuWnaLMzp
FIvT3w1tB3/ohNwR91LQayl9AA3LI01LpdXPNagxdAVcpYj8cI79ctvqjYl3Qgc1
O/VFbLFE0uJxeA7j8usIvI6hyTJY14zAj0eTeSwDK7YjEdbcKBH5wrK2Z9j7dPhp
tAmSQjlPUETKZ7keeu0MSZQIMGsVMmP8AdNk6I4C8cnzr4q65J7bEYPhL6PsleP8
gNYth6tmQyhDv8/CpfSBsTuKgsKuugCe1DZ1SqjrOpcLiW5f6Xp/XhK7RINwDALV
bW8Yu+dAia0C3g1WF8b0c23xsjaY+8CIVT0GouPU+sALNNp2VQnO01dUbOGb5jaq
iU4m0I45rWsDN53ZaMNex805yK3b/eFBzcNNuHc2MlBItxzckyU5TlDSnQ3BejLz
DWONKtqJ0/i5FGn0SJ59BsgxBdm2YcbbxZ1F8tH6LsmBKEEuc6fh4X3685lDOtHf
/u+NSAk7rKdY9GDSpHI6qLg/NdV1DkMYWx8e+uqKTas3QDwbMNs2p12iSjY2nQlr
GLggObbycc1ixWS9oNdQpenB2v7Agl5Z39OgcX1lJ1WnhMyiYPUxenwyEja1CFwQ
ditfZzEUyU6LyxxvYmpoh56g6M/3wiQ2wGKP+unME+UWyYM3KerWf5458pxWHPeZ
xBl8qZ40B3wpWOIaPOyAQAYv4zRgtK2FQ4EyxmXQ6/omWiysjtcdHvh2iSyvq8/6
oIb2kA/OF6yHowCQCB5AjZWZECbuKugXFOVcdC9HXaZZS1C2JZQrtAPB9areMLS7
ufJ2LdMNZsEu6URh3BPAkxMXePk8xjowM6dVkIH8OaHB9LmjE+tzD9BXgmrQobS2
50zqlmZW5UtA8UgDxRljYAdY7YE3XcY8z3agFyHAKPymRndrjLI44XWyPzpL8TQ4
tnPNt3OEX1Ix/gjmDp/b2Erw/Edry/tTYY1lRqLaE/W79BSM574Bjgh0AkO+RTn8
Wniab5cRpRerRvx+XKFOi2Xpvz97fQ7DbA5MPwU79Y4vZZK+uQGQaRuPk6eqECrM
aTVOhuuuZjZG2bpRLTSFTicElLL54i47jX3rwtAUp2ncFHgzQ6Xz/uVJEvVKGR83
H5uCkHjs/Iv4ddnOST1wPGqF9XjHHrFdyvlN4jiIN6tO84WXRDmvz3xN+hd25cPe
aTSrjP0D8HgUMAGc/hhlg4AUDdWRjbrKPXT0wavQuZyuTrJ0oPa8d3PhFhHLqM2U
5QHHWLHh1xDNcVslhalL2Ubk4n9hJdy3s2hFdmPuiZpGeyBKg2z2OVD+yrdGQFYY
A1TT3hsCf0cUlm/e62LO0HnGjuLCE/lImQW/H+HGFWT9xkztUxzYUn8vzfWTlwCX
RAqFQjTp2rEwKYGOLlQrlCI/ZukbWcsqgsfhz8M5RoBzHkMJgeC/+Y8LjFeY+T9m
TKLB+sdJn+mOpZyA6QcL8oLjYg4L/r9imsbhi/oLym/jPViU8Wl2Ao7YAVXxhV55
inCHpfoxq/ue6xKgjH8TSInYmhwSEA2HkoKqJh4Be+XyFnOvcx5u0oj8Nhu/utmh
ygxd6ogKcaEUD/hDwu/lefkW4nbaZGxMoK4tJLi/BSdusW6b/wu+6jod5h8I5G3D
vJx28CbQmpG8N5Bf80TuZBdDHEDHV8SGERMqydUJZScQ4Uk2cCzpaSlPnKfUQ+md
pGsYcLYZ4X1oxRFs3+ecKViAoPvVXNcTjlremywDcGm02Sqw7poWKZY35Cbyqhab
LMaPZykgXJ7175gbQ/tmVUEMZ4FPqGSJrLLKGNBzeUEXZfEbDIFpSBPIsGMDbQsx
3tqz1139agP7qKXcH8p5VJVvS6/IZuI3lItphET8LtNhopfY4afk7ejGBgdZvNYv
6xZDiaUOa1RoMBB64Y8BP1qCwviriqbUYvK0uAeFnoyal7S5izxkUsS0Q3+AgSGW
/JcEUwybYmyTVUeXn2jKJK/4/SWA9QB3SSuGvWhJiMha87tYzF6kCXqxdsz2i77/
bLDq/yo3xYcVQG1eWfiFcxuN0Iw3WnNUvzexkUgvppg/+EeSf3C+8fP8E7ma1w4M
ZOcNiGrwbmo2G9n62HnMuNmc8S/B3HocGgygP7kpPuoLXj5TZBFwsOhdv732Qo9u
7N5Bhdsdmb2I5TQXp78hpRn4zIcLvAp5Fx2/4MbZngInidnJctMCrStag+KdXb8q
Mw9OdsqGVzU20jNl7rR5gmvW8+i443xT4wu+zaMbTRagi9oms0VErzL/4SDEbFN4
vdpg4Y0SMbmc+CILqJ6Jir4FNjM8jsytXvPUyjb7AgFlnQfghtxwiVtRhoyRBWWA
Sra/3n/DnlF3eJNK8MXHl8KMobmUI4ANqI55ytlxqD3Y20HztdrFz/Z2IcjNtcYs
T424Fcbh0pCgNCAMzYegOEOQhuV93Eu/uIw/ncXj1LYM1iqmnJRs1rKAl5UDUh1c
tT1WrQ3chqy605x6aiS+V2O5y79HjXKyPZbP7NU8I9ZAFLybJN6e0FAN76xDOCJY
cHy+Tt/vMq3RKlxsBxlV7FDcB7mdvneW5cbRtFYRWKyTPoCVtnpjAK+xh4GYzMn3
TroQ+EJkJQ7wCo9vB/0WDT56vyZIWwZV721tJ7ZRy0xULqsq5QaYYIvpmowAY+9g
UVyA3aIeoNfPTZKbuiwdGmSK4xKLZa1n+ylXUVpmiMRH8d4pRsn4NRqcCbJQyrRv
+VCqIXJGoyl3tz3WJqMV3ngkoFgUHBXB+Bv8imQWB9jsNpbONTEwL5M7qNjTFIkS
K8IspFVu8duG3rO1BifShnNB6pnKwlMvraAuZSvnlgXbG+1KFtnv6zHdx5FgnIm1
ZP/Y9HY0StknwLckon7MMNUDDZD6THxZ81WAyqCeuzYYXnsGDxmO2xAhjcnUf3EL
+KQuRV6D5o8Ugkj2g1lWhApje+yrjVStyA6GGtLI3IWxHBAcl1+kN+tgqwSIDNZ+
EsRsASlV7efANa0fAOgF6n6G9/UUmKgLxGDwy1h4C8OYwQ1f85SCQSVougLrrZ+y
ExpiWBGVUX5cwgHQddqhbjdJ6G+HhA7RB5ZbFsoqdik7wxlgiIAeMP3sRDAlAdq6
9YrMbJDYtg9F6CKUmV7vL8S38LY2+0P2VYEPHCr5D/WKczNW/czRDKBs9qWQquk7
1/rx0WzPt6m0mWQW+LZ829JpsSLm/D/+XrDu5eGoDtZOWbf6rrSbxoFvGhlve1vc
eLlKZViBvcNilQ5s1HCK1v4Z9vacS3B1kuDTO1DwHr/6XaYORR+DFhy741kMdnCz
IqupctUjADW/tC+vw81qowMGWgu6RYSHwXbPJCBtUQBvEnlXYnZAt1m6NuVP2juD
ARhQ0cFsoIjegfdo3UCkZuxgiNdE3kJf+mToMltPfikiogNor3ceBQMmYc50iOe+
DYqyfAvqZa5NQ/oLVeZATDbZWSGc+ABssfvxG4LceyDcqKGXIp+N15YDsFtmvhFM
O2sT8zl4Xxgc7QZD8UgnJMB4OQ27gcK6e7m+671UiN8xhfwgFiCQ0mxGESGLPW07
zVWiEN10MP1g/9cJ0jCFicsul8PC6Bg/FdJCZXrF2Ykv+2Nf4kuw6TQ/00pHf8uO
o0eaYIjiqPMKvycb9XYeN3PRJS4XcBfdusqUeDMLMzts4/T1+ePogB3wWaJaJRQx
MeuveG5NeMyjb2pdxxwpACqEI3ErSa+w3aHHd35yFcHn4cxtznRTFkJ22WCURxoc
AXBtX8q5CG51fEOuzS5Mqx2/ZIG+JvofCyyTT35YuLuQnczCAvuT+9ON2s7Z8tnH
5HaKVjqmhmhZ//439O7yS6M3dMsaRmGgxNxASaxSW5P6Yfbtdy6UVCoUxrh64z9l
lrLDp5Y8ZFyrz59g1H2HAptBnNmwFZYfNvOdS+wp8FI9pCOyp6LK5HHb7RGN70da
/3DrOs3iSamuLcRwDFEfrTFlRR/4YuzSm9cvlOk68rcn32as+uow2ZQ50sGR2vpZ
myOKrQE0Lnh9H5p18FewBysmKrJrEC2bfT8UXZU7QLldwj9xMETMwfN1Pf7rM19Q
9uCRnDx43Qt+UulKH/kds9eIGUnfaITfkZyLOb8TrmLjd+FxlPTkQeNhSSLfZlxF
qzQpToaCR4A9Es5ekzdVueGd1lJ7mal+Tq4/LvZ5hd6Q3l7nsdHec1l0Jx2vKtUh
YHlf2iNonQcUPrX9PlSKYd3rGTFcs2ZeGOEfTIzIHcDwxKtE7e0Xrk58KTjRTh3x
Ng670H9roaPwCFnYXBvt+rABG0X/6kAPGVjwOCSI8ZGZTc85aKG4fudi7/DRswyV
EwbIEviSy7EaPBl8kmr2In0VSGSkyliG/KZik/DOX93FCwOFEjuIC/BaTYvntPW9
7F7lh/wE8Mujm09d33Y/l9VmXKH3MbvzTzQc7OYcrwniBXk7JsZPLQLcN886l8ef
DZBMNC2+K+70ns7YllgdyV9KtZa+31TRzx/UZOBT5XigukCRTwtLNl0TyJzdpMq3
kXnaRhvYNq3voY+5TUbznKCIYOR51Mq0b0YIWx6GLkzVJ64IGIXvkO2WhSKCXGB7
R8zSXSNEYcFoZu70yRq90TBCAHFfcPwXCsjGHOL+OiltOa2+fTlnVFqutEB6Qg5G
43anD0DwLKFujRDIpbKqoRrbaPp9R7WjC9Cf0L3t3dPK+yFcK7656a7h6DRpKm1x
T8793YWcp5ke2muoQmKZ1rcr7xfGDTU8uZWFRVzYANKp2xLeRwStaZ+E3VHE2dYD
ChSG4xDYyOpP6o4RTNqMMk41C4wvy1CfvxMmqvlkO74GtWNsblVrgZOdRHFE/msl
1kBBi0s7dG9HHgiQ0HV2fRTZBMLDD5MUm1xiVoztvag131+mmj63FenV4FxrznyM
wZ8zL2HSm8jwKMTSLTUfs6siWtt92YEKHfPiZNwj76hDN7stik6jA+kEE6P6hNRP
cah+WRwEi8qH0kC5A1Ik8VaSO+NxwAnJl9HI1wBv0oiNJqcV0q5lysTnCO65027H
OnXRlmQIW63Rqva2Od3ef9ZQngVReiYMoYRYY9DcJ1DGDiV3MJSBiK8YhZfkbHxw
XzmFwCAwsbRb57icK13hlnxUlHDh0qOnflgGG/LSS3KWnP8Wle1eV49Nl+BRwwD1
/ku/ofYNRQtcDKzvCjOYxIDyM0WMxGoiH+J4dkqzbZJYeC2S3xfNMJmDazyKc8k1
xB8oWLisUQqdq/QMMB+K18Da2EeH6QJHW/ZCHE1FkdJ7naLcN7k+BVdMoSKrUQrT
UUt4U2jmo1sScKdVt0Z2FV1My4EcYsAqTKo4zPZCY9aTr+kpDePPwYB39+1itS6p
d4BirP6xs2wZcBcuPxWkVckjmU4XfmGg2K+kr839c8pHbwK0k80UttXs64TywNKh
8j4UiBSqa2PhukPZ1ON7Zt3na8fXNQw9BPtFQ4ogWb49mXNHimk3KrZv/k/ZQLBK
OMn/r7bC3o94Dj7gcscuXNsZbrFawVFC5sR6oV4J6krSn/PiqK4HGlTDVFpZGmyN
qj77fGNjihwhQMYSz5zp1+H/mfEAMIjMKsHXMAMunvpx8Tkt2MJNN+qyU6dSlbkE
gbAYvGCTeN5X7jkDB/cAMNiGs1LqStoniAURcEtj5rOtmhwo00y3KgE1HpQ2gQ4A
ixUjGNohi1zDoXA6v3nPv0tW/wV5+sW+VRDsB0yfBHax0ZyWj8zLqvkYG92Z+crR
ZOqjLV8Tm9HaFj/KKVE/2O7srdFSzMB9X6K+WsvOVH39Wa1thy+GmmmdSd4xy/OE
JTdmRCmN1SgyA4w4ODAT/XOhL9D+gQTBH/FqZwUm+ZyMnzppnz4fM1EDiwse9NOm
1stFvPfMOlOPLf7kNIBMJTIfMkhepQsLyN5xgTaxddpVi7NJhhOi/eLiJPZ+wRZC
Ooo6mq484vL9DpjkwPtTBIFqUjUUR5lSrHodMK7RaGVIJUFUv89EniI4gjGyzt/n
qrfihW2yinhWOsmBYtEbhKaREgFmmZBE5fYN76xzikSWy75Zarr7dh8PLyn3ln/C
7gWAOU8qWqgt1IhjtJRZhqTzbzPy4r+M4LvLbZMUugL0Kltgzwsuf4793WLkmW2S
kDNWT6NgShY2Lmt/FF6ktRTfoV73eFmLgGXOlrxScb9AIeYGk2wlDilygLG3w8CL
6vOlXbk0jC8CnyAQbn7G94jciUtc0mULziNYkAFqImyCSnkVYwzdrwrhW2WQeJdk
0GQ6XFydW0Z+qMGgLpGK0uSwN8JQnZvAfUC+stU5//8xYsyBe/l47Za9fAeKEriu
LIQT74v+X/oU9ivBMOQikGMPd9SS+5MszEMArFN3YQUEMRrwhRvV5rBcWVM7pBuN
4uPBGz1TgfBxfn/2+PZxed2Tt+O3sbB2iOhNraKxj3KnXbV+4w1bAwykRBgtIYS/
R+O8xWAMZyFR9sk2yfcq/9qx6w9R2Pq/02GWet2l9aXHVUtJcnKzxRPgR4Tkrbvg
y4+/EonKV/v64mRBt0gvL3RE7F0zwvyinlRVa9TZL906wKQuHYQEOS4DzCqoAa2C
Vjqsfgt1qQyBO3rdqN/PfV95UqAMxd88YUfjZH/OPHBowQrWJtR+SSszPAdgnfO2
Y6IhpQrBox78vlrWkdvTNu/aR3KI+9dP8GLidB3Ac3O0Wbo/JjVMTIsG5MZF3GuF
P/n9USLu00TbZQKEwI7AHGYlI8PTsbQnmyYPO/CW4JMCPBM9IjUZ59hrPx8TgbTA
uXDo9+bqXvELgHFNnLJ8NwB3m5qe3/nXWILF8Kodvt6aOm/2ZTNtwOlJbPf7unIJ
ZLsfAyQVSxav1SU5sj7q/dP6ypf+IuAqd7iCVeRypjoogpWospMT0d1ZW/LxHPH0
oDVOsMkwo1wJOdVDU3CWgMfGdf9IlLyXgwCCBRKCuntJCdF2oe8e4ajeaFU0x4nU
Lcl4bsvZ4Lj/H4mcCB5RALKQws6c2SVlbhuiLfT3e3GfkK4jQQFkKqFtN6Jpb8mF
ldLpeniGiIYgOZDFKimbrfuIxLRuSTC/VOt8AfkRZzit1Mr94n5SPmntx2/52Pkq
4enm0ir0uXtfO5rCTf2HLPN5YCFmO2CDP59hOxR9RiDiSo8+Cr/YK+u/j+r7xxUp
DQoePkhQBKbtv+rbElyKbRzmg513J5lbxf27qu5b805ZEUpZvuY3mM5/lon2dQkV
P76oZXvFljWipEkYMY3XPrW5PX8H22A/sxWMo8uz7OT8c7KKGxFCSv8ATFhlCAu+
ihRFkGXiBViAxQAqfp3NKktxnWQwkAosFwQfp6YdjsPV2by9sHgGkTdHPUY4DYPu
i92P7qw7s9eJDe8MOu0VSqmTDSlwzdhyf9ZbvBFOuiemskwMoeu3fKLSKKW/7uIn
8ppn+1Gx7XpYMhWC7OV715r6UnomOauZQ83nmjfqLLZDfSIXIwn/DrAcFgLnA1Pj
wmMl74Xvf7wxPawBHr7lr0HYdESfsuRo+0kU2gNLAVjRS16n70mKIlaj3BcKTkr2
1IpcbpO94Umc6f/whOmpdZ6ia9AaQF2hSe7rZiVpbpTrJYv9+fj1LXLWBszcMX97
NZlANJd8C636rK/ByPfGjdl7reov7mIkb6MBtXKK3xDyXAn5u9nX6yZ/TlxdoPlT
FMjgawhCqAhQb8A+lCm/jfcedCmDjKh5mejlh7rW0JLNRTHIUf5uuxsm7luZ4d2b
k1rCw8HrFiVMC+RZBlYMY77jsYMyNoxP4JxLt8IB7K7Ghahc1HuXTKAHjllRT5X1
f47/19/QIo7epKJ653LWFAqXt256iKoufwysnpx/r8Xzcicpg2m31oB7qW/cipI/
vTdIfuxnMUulUy9SpDvj1uKe/NG5WsuXeADSD6L0VxqwhySY9dqcJpKpyiluivER
Bx+oR6D2PRgtHlg7zN3iUCY24iOTy8CC5xOCCni0FLcM/c+LtPitrGPWw9vXMseB
BRZM2Sm2PboLb6pobvLvtjCXWKJnu/xCkI5QDWgBAkKfg/ONEo527OwntiHRntFX
94O0Q/R8gkucMX/WqfetEZFw0KyZi+PjtMNAnSWqUlfHXDbdilB8VKEv3IS55Fo1
9kMHep7v6YLG9A7Tv5x5bLIt26BGnq1yTQMNSa3prF1QzgQMK05xNPRmd6lZ6yhQ
/aavXteT/o9kUE/SZpMaFmapCtGOaerLwtM3fbiNQx6aNtygQaQTNG9QVDRQcuqE
H5iU2y8+Y/x4k63W1cWV9nsc868/DRSytHZxJ5rc8lubZ9IMijKaaAEP+KAPaRB2
MqbyJFRB3NJAE0J8g4AxNNl90Zd43OuXzYEjycqentXFCuG1GRAbyyvLv+Cpu31P
wDGembjgYfNGd/ykaLbyQWXexqXuo5OhwwEs8+95CHeuHpth+diEhO+Sn2pTa4W2
5tGfEqHmRX0b58Rfo5B14IKTrVUcFCQgS1qBh7OeCPR1JWLsjp+iFloiJPYE5JCu
5vNnNZVRhFwBqSfA934APkGI0fHoyPbNGW7ImoXR5+94wM3W77IWGoJIOvh2i7s4
oti0ks2ewgYD/HsC6MWNtVaUmoP82ob1DHlHCZnfgl5rAjcFG0/FMIhIthQg6ecB
hRFftr2+orLc+TGKAPZRnu405z8Wiy7+LYFBRY/ZBXTb4pr6cpEr8ehfvyE5bcna
LwZ2xUW88or6MYQ/T3b7htwz3HYyO/8JX4o77cQYoZDqqBB0ZNHWFQ5z+4b3g0r2
smyb96GQheBFtNFWyRR+9cf0WvQKEMDEF3aPznGGhgvHy04g0Tqo67iNBSMn/NNO
7qSXe/4khSMD+VuHBrUB+OGi+U8kP5Z7HOe0/2MSi2Ngynl4y03idKkalBgftdQV
18bPfoyaqKCJvpOB9bg9+nwM1zg9zYudLTru2hJEt8DVDodSYvDjdmUHZtJHd112
8h+BqLzoBLAlJyJXIVEuiqgDFuszfgAXluorlOfY3VZQkQSPRlNrd10CPYhcJY4B
L+VROpcT8r0WMl+iV/8xTO2mmqobTDJ+6VoPngarGNiK9E1oaOnZCTwi1Q3lkWs8
za+o40ox/gfjbxaTs8csqxjeeKbx52fvzlXzof6mL83W8h6DLcAJbMkdXcaFtBEO
99wvd5PKtbE/PIgQwP+cINeESPnvtw/afmpE8RasHnktaEczSbkkpb6m66Yvqn8C
U3pO+8nk+j4QvM7bKsokkl89zqop0jht9j5gaokDikyi6FbqgBDsbkPEWnU3wYVJ
rSHlMmYVOuS8/IGoeusmqfcRXJ0Vfz6V6k/ecvVo/vUQGFNU21rwgX41VjaxJs1h
5xGf6DFB1qJWSjV216dIDkwXBAibFcYrqxpti6UMLXhraSaMVSk96dmUk6IoSRC/
MspH+JAn/6W5/61aJynNrVV7hT1pJD8s+gBWfvuQzoUf6wWhi4I8wVlK9YeY96sC
U/WRW33TK4ChKxMtep2kZzFBNyWpV6OL566o0XvGsfMzO3jidBmDMb2n0aCIs8z4
5usPRckkF0rIXYeMtw9oU5exDkIkwbYJbxEwD4nTtnZmM+lafqp+YRA6ZHWPxsOC
ODmKaNbnpBDNDS5xwm5AP77RfWVp8ph8GE63E6SEvBk5QpzFi1Y343zw03BK1YoI
BVvbk1UnbK6MJiqTxrRPy9scODjFEecWCV5f0Wx1LQjRLbT7FPAOLkKGxvbvJLHE
AKdBrFD0l4Cz2srncLuW0NVo40Imb56ROL/ap7k/Ui5IvarG5XSjkTeDST48616+
dZ9Fx/QNzagD1qlC/w93Tbyw62crOk5cPYqlP2AjMYX8ltSfVr60K16TbfGpkPNw
25/H0zzxgs+nyjDBhMUQSXaXv0hmq/zV01Xx7HH5sGhyHpvNPDGXEtXHvJyKBJQI
VWYmXOO6yBGXZQP5T1mJA++C+UGlj+KqqRRtMK46ImmXBUTLyN9wyjSc+0JXp8Ww
7XH3oGK+r+WKlBMrmZyF7KsgusFfgQU0y9ReXk13wQgkEpmuNW6/gLg29i0WrKJB
aA/T4hOSpCFM2a3y5PRxMKgBdVzrRdi5qM6i7tGOYjyiUl+lL+uZOA2E1/r5DX4m
KN14VBlYCpPUlooUqb52hfOQKdQx4t1VZV7fhNHpiv9SBlKfI72D9XjXpLJu1FM5
I0Q2xZGre8iY07z3oQ4/66O2tuP+I5qbAotuvdwavLrjAFZ49D7L7CcQLFDownBZ
QqLqCjwTAk03NchOLVdQ/5/Jlxf7p8noW82L40vgrPkytQJy3N5GII2QX2+/oDBK
edF5NFw+RU6cDXHzshedm/zfrdzDWnzrA3BjKSbHHqXpsKlLuBtxNSZ+kdXVutoZ
SpjvHXcse2J7RYzOpdAHPLCsiwPDZOdwvEcVOV59aA+2TVOVfZ4+ytWLihGcu5+W
4YMTz9F9as2Ri+emGwtg+HTn6e4daF+f7scw9ukQePCvvwe8/nhRCnPuVFzUSaiI
jAChSpIgpii5d5CtC9cl8F+0v5diwYM8lDIQKkOfnDIb4KAmhE4I/fqAy9E3Kxfv
ZKWwcSIChIz09AU4EJPOLxxmF1D6g4r8eC02dItM2mTjHZG+kC+dvMpBfWDreBx4
ZHVhjHoLYo9JMrlYjLfFQDUaYujeeuHmRhNpexmvLleUlwVWwR7QjUCxUiaNOdAZ
9plMT2Z6zexHCNwmX49V+JZGT19imCk+Dd92xrE6N4Q8U2V0PK5GTLT3vqpd7/ec
IhhQxIVt6X2xRkSURZBwU4hXmxuFekQk3jLoLvq1vc4upCVEeSnqR9ySO8RG6l+c
kv0+j8+kld3DEFc4Anv9zUcfEwv9iZdK4uMM52iSEl9oc3gAo18SeWaPbYO3NcDU
QBGReFLMZbCerteQq/EbyvmGgU6/Py2i0kD9Y7mAGbmH4IyHsPqwJC3XD8dSM8P2
cujl9DRLBw67XaIJ5d8njGc58c4mF+Vppk2XaWAhpDpr9C0yKS+4LCtBOzdF9fHo
IeHy7aZ+kcqbTm44a+tAw9rnOstoc7gqg+XMyjGnSbURZgVsR8q27+g8JqozLu6F
ZoWDCZYMFC79GPuxg+MOTbrgQ6CSOXUNTNA9OnyJ7h9DAwyKWP68FYW5du5W6rsP
hXzD/Y6yPlQ0i7bnNo9MvIrGZTWkJmzmHzKVRcBkwXyINGwxppQXB7TlaAfITRJE
3UPpF+JpuWcEK3iX6+n9o5rUw7GcqHki3be1Yv32BLAeiJLT7MNwbio0PwyyhtP+
YDc5lY5Jw2dZ4cQeAIodjVNm4aKgXHzora+P2r1XBoxJGNYwtImp0qQnOd8B0rF6
7c6xrZlefZjFQW4WbsysGsnMlcVU2gC8JPuAzkTOZyfI8Rr+3RCcuDzUy4cDfwRJ
1g+P0cg6Ki/DslKJBm89TKMiOmvceY6dgIq1BfgoZIRomo48v0lon+oiMFyGPTO/
jWaIZ4NkXtE6/3a4EFI82bn1krndAK9x+aZC7cghuyRlqe6FiT+THpkiAyVykl8E
5XhSSuYHODAWD/qoAiDOu/9E69BcnQL6etab4PQzp1PQcWQ+gJMVcnMlE6+KTzhK
ZY0QepFCtNS0Z0AcaoDEmvyOauZKkIB8xngG+OtyQNV+fKLhTQ0kkjPEIH2+HZoL
5ykzT1lADdO/shHoaV7oQsS1o2/3G5sOaO+MqzqjoBxkQ3AmoCtKMvwUVGSF7Ycw
EvsdkFdOzl+kO9psRbBi1tFQBqtLxyUykwvMV9EXbUdkK07IccibozZmZ9UehwDf
7B55t6B5OtTSq3i6aFU37MrFhArpLMb2/hysU02++Lq5zQLiJ/TDugSV+3QwTY4w
oRkfF3bn1nV+OglUWuKtp1eWsZsk45tvkFWkMti2lJHLyRIy8LGHe6fmo9q4+f3O
iRNYqgrTvS8wN9z/ekP1ffOO7uNCPmGl3YH7J7ujTnh/gm/Cu0Sbjxdq6BRtW+YC
q2jOk5yvKlTc4d+iBSC1OVQMnLrBmOkaLIx4AnK7Rtu/FaZx/QDEnfOf19QOu921
QDyFu0JQh7Q+I9BszZ8LKB4UnEk+Qhjru0XtPgSzNpQzCqzp3Jut2PZro6IuzSp+
/tkSHTExt/SWfqcigQHb3DuND5CIkD4kq/YD+kTglKDwoCgX8L4OnkzRRAykmU6M
MWzD0mhlGKEsABkOJhZ4ol3y6rejI5/Ahlld6biXkODVGdC2426ZWzrOkCGRkV4r
W9YKqKReR8+RHk1ufX/ZzmYlNFhaAUBCT5wUT5pd4nSoYmLsVZNjAp2JhuRi+BBZ
cyqnlY1iX7aXdq3xlMAXCPWX5FvLKs+JnRJBneIk0f0DNxrihG/EUxQ1N1MSPrH4
h66uATmCUkLJ6Hflc4AIfSEa8hC3kKsonTUMNotqoqxwFAC0W4LPDByq3NxCRy3M
qAGYPE4tni0UiuTP6almSgrSXWn7bo+QHGOcH+49WtIulzpffHvK/u4gzDrkESRb
OHUCRp8BrSrpsT4qDjTteOu/QCHIZLFAO35YcqQXficjfntWtm0QEaRTNQiHU1gG
T9POEHdNR7MHcVS+vg2WRZ9/bdzt6k/vjDn8srUEJ7Li+vHBLeCnl9S2CXLw3f1A
v8jo08zNnsI3PQjgctd2Por0PDOWE7KoYdIE+Pc77jq+Njciv6uTF1P3ust+uAPI
NY7X+EHixlK6fjPZk9/hqqbeQkH4NcTznmNNkcz+k+5SnJpValPd1dPbfQ4ehuFn
eK2qbtsrzZ8GjBwkcAV3WwBCLvGdDYEmt5wLneilrp0DGjFKVOYa171W2tn7vIux
WH9lhsJzL7RhwI9hq6yo/GWOm1wJqftVGsPfQoH80puv+RW4WmY6xq0ogdOee+Bi
I3zQDXnA1bqigKt5n+6D0YkRDQmvF77g/wKgDSIjVQW0UDoHM+BmISEBdaG6CtH3
T/T/v91fPlL0YgSPv3QgbAXMPRR1v8hLqT182nCdH7IsH6+5Wy+tEdXYNSBSnh8k
FM2xkd1Jb9lwp//ZZA2bPcTGnv/p6XFacOQwWvgWjgHBrvgr1mGtpjiYyCdcK7Qq
42BwfXa2l6vO7OJQ9pa/B14cy5LEe+9BRoJRbUilQ7ikS0B0Q7cnYnmtmdgyjm12
S3fFpbpmhUut+BubViDATB1+h/EpgGkpdgkJsLYRYRGrn8obuxJu89txU7gD64+r
05o2eEo4hV43E8K8eDSL5YwA9ZYQ6f5+jJmSqeGL6/1j72+oLbhcK2qrydMmY8Ud
U7rKleyMavlgiV+b70FsXSM6fTh7zwdrUraJ4IbFIRSFyLwShhvek913yIOEYA5F
NfOD85eiLXuLMkfhjLuuWmZTnsIQCJ4fSDo0r/x+N/CoDhB/x+b6jha2n5yfm1DC
RsDV3lKYtoxFtJp8s0NJ0CF5ioFBX8i8WKnNp11lHU8H78i3MgNnP91m7Wuy69gw
kVLtA/8YL3C/lvIQ0dMPnX+HMwVHJTpJjh7Pll66UNmEggkB3C9dQ5UbbHzRb/sl
KbjJzLLWApkjrDyytrgmTTnHb+UjWDlMuaa8LW5AeEfZDFWhMITwmQsEPA+M99xm
nQUUskln9pnTyngca31vypHwXbUfuHiv6hkX+xs43W7MImRtwz+ZnMujY4HnEkGT
xNFhOejNOlNj81UnvXl/qeFdeEfDlAw5GlvO2H+D9THoq9JX4t/4aMaQLMvco/yb
x9mOm9dwX4VM6DhlETRJ8dkU8bocTAb1v05nLUKFUfvbOi/EnDq1bGOeYlroZ3nj
elj6ju8Npkp10BXB1KOMHGZefppO5FFEAGLyCxW9p2vXpQIw0MtTvenXSQLcKidU
IDVgNy/nZx78L+6Gp5bHvGuWJzP8AoixVlPeGYTdHZLM4olsG0FUcNdesg0qJ4Th
lM1CenZBRqmIGUax0F4k5iPTRqoYOhBaoOYltuY/m7MsFJNtjx99mKy1FVXzpXIt
hyF2Y/7QwNRD030xCLpNCL5UdFbZKMQ8FGeHRFI89GTtPd424jl4nLe3dzEIr7xO
wsWjX0mh4IdlBwfpa2KnEg93BKnzDN9LV9M8Lq6km3jvSiCwd3kOjq0916mh0Lru
zcQzgS+UEqCVwm3/bNjfzbRUilHe6zYRJOFaDk3RO1JBGJXKaYUXKSqPrSXIPDZ+
i1caYj46DE1YqdesoOXMADi8W626fZA6VazxeUykoebRe7qes7nRsyDJzs9LZHQE
WDsOXouo98Byp1f8Sp1Tw0RyXTyjkE8+kmgQTdxEK2u9btoHOOVydJCsdTdlLivE
NLhFB81HPpzOlf+qo4b8ELXSSXLIVDQ8WjXMmEnpMy63ZlboxLwNJTcMSLNoQv74
ZHnmqETNeOE8tDNLuDtq43Wtpzrfm4UYnB1v0/D4J+BTWoNeUgN2zrDbsP/pJRbH
XqppLzh0JmR5URmJdCSxVTTmcOkDQafwxvDRKJErh7OSPP9PHE6dCHyNzk9qdlmj
czZ1a5pLU8nDF+QS8bH9U8h9M6/MIPGGtsoIB4xhtPraaD6vdFWYA6jkDjHYKrwu
VR3QbDZfh4HBDyGnFyJidLQZwiP8e0V2C7JMqHUR1dsQcvTIIc5heePF6Hp/iQMd
kWmmJCuNcOwWc3LXhQWIVwArbnwjJpNa4jp8pBlSlLeLN2faZUjh3115/Y1AWVZS
jLLTWonYKUjcyuldL+1SFS/GFa+uPJ/baktQOjbPSQDwXxbaiZqtZVpcpEWl04HY
KFAWK8FCJr59UlWBHTzbYEzAq9NnjlmCRBSi7b7hwqobPT+fAaH23ceSLYVI1aN2
C3ct0eRBERFKEHu/W40CY0/ovdgVqemnVOuB24k+IJcMvP+JSULIQ16WC6dWflNt
MObz8PiOdFUamlnxR5kQUuiQbMUZaRm9uKmM/9Y/usheNP8thExX3qEYhAgsFdCE
bXDdFQDQ0Qt+EG1jFkWnBZo8+Y7jclNLl2mBJCXeq6piCZ3qyuaIk7xEc2CIV9on
UlnWicdAf0Q22Yf+VmSkpLWaYF0GGHnHgL1PUlpyWVBNO862gkFPsipA0G12eaVM
eOgAXKcA9YhMAngK3V2mFSQ2htJctycXw7uJ71FSPgh01TyFc4vzZ3gP5YQ01pFl
zXSyzVutZE5i6C5KhyF5wU8BAY/mQPPS+iz3uKgdnGngQBjCVpO0uwAuj9xmDtBJ
/iS3m1JGANegl0rrf4mJnJhoRdvkzUOv8IlftrNS3SoZLXZfZKFLlDot6DNX/2nv
KaICwi8xinEW+uEE5xfiZCbsbb91yQ72EhOjqP/rEPl4ADmtym4WCOSxeC/M9NR9
wcSA0YajUqLH98xMz9KNUSOWtrDib+rXaWK4PYPk1+IGthyg3mxWMMwY1CypIBiL
vS1YVuW3tJEpntJbcAAL5rKj3bXPa82mArTS6cnIWDec9g4Bbzrlywc2wj1Ab4T5
vauGC2w6L3gR+U7atu/7Nu91IkNg7yAPLtM2l8SW8A1OyrzByF+RnFG/KUYJFWYv
v9n3JHDgMu9OHngBeqmBb6amcHzqeYco2VpUxqCJlvmX0HnSgizRSfXD/zVn1vpA
wLwFAMn/UbMhfOXG1B1hLXfWpcQNtFc8VZHhO0LqmQIrI1c1/HdHmYeI6FPSTI0k
6+/XG93XyZwpezD6lX8ZjKX4Fvn49MbU0jmFM4zwZbAfYkCtHvWSRTmoVdq6sirN
jb1Jcvmyze4A69qiUMr11e+eivJKrDoIccPFP1aMgQp/+70RhMoZZynGomR/kpNW
EcEwYW5MJFCvyL8Mj6+BE7p9/xNjnaq/sk+n4eoYw8k/FntDiLshq2xBULZHCeWN
iZbQ480NOuUz2+Pw5AIQCHkIpIoPDUi5uz5RV7jf+KQ+On31EgWiTWsT4kllKWzR
ziv6MEPAiztm7d72oKjkOBQWhHP85Q6K7Llw3MXHJ0qdzHHFc4uGbOwUlQhzEBzO
Elp9sQ3foAkqthFmVXbtT4993X59Gy7Z8ybl2EPKxnwmqU/Uoit9tvVqJUZL0py7
QkHG9YvZE4fncinwBgQKbwiPj8LBSRV05LxYl3vM1qjaLWgGg97vzjjeYrRXclxd
b94f1ebtx+RrQQN8HOZPtWD6tVdks8A/gopWpVWgYrh+HmvHvoRSyxZr73WAxQd0
hhFJ4E/mr/mD+lEvOq+CTI/pb/ObAVNrMrn4/GgkjjI2eUXb6LcXH5GumhDAcfRE
qB92Wz87UXLPUmyv05cncRL2jSt+Te9+svSecG8z6zb+A8dnkWRKgEpgt7oYzUZR
bY5DrIyWPQXC0Pa+aZd9Ua4elzhb/y+lpT38NHRYO8xH//JPovzop+1FgjNkyjsE
0lb1+TxmYKmVHEU4rqlqmeFHUUwREw0GM5ZyT9Lo2uDjIKyF6m1DV7EORwBTiOXO
E+xWQ5DmFJKN+ZFmiCDt4J591jh0YdNWmtT4wj1cTCGZJUeeEi4EkG95pB2SkvVy
/olJOVIqkMTYf9CYZuYK9fmf9lqEHncJxG0MEJyB72D3zSpJQAjYEFerlEky51u3
ta9wLKkDeCQKJjUALcQnuCmeyztPoQSeW72H5ddq46c+y1vCzgIUiueZYLNych0U
IPsxb0DUGZdnS56NMb+0rCGgy9LLT+OrOwJqvZTyicSodqlwQvDIrY1Dzjqwh/M5
oFQ8S0ZX1sdCKtsY1Yj5ffVNbQ4KB9+IP5kh1O2aqpFHIaQZSrzo1dgEDAFoJm8n
r1HGdevyEAGMgLGAepGL5AIEdlpSY3EXEQ4bruEvfu3ftMO+O7mzSmOruTuLuX8d
ZDnGvM4DcIVmPCFWmKvkrMpH7InhoZTUgbpUETAaEQ70biuAfeWsEui5Yb1lwTz5
Y1vhiTtWbU2LQA8kyQsw5HoUpFJEWaHYtxCnMXNbUmoKH8vXTzx3NcZRCV5bcklc
doKQS16sVldVlWIYqxKnCYhAk5H6ib+lTH8W+w2QFHQRf/eIpOVSHpmik12CA3ew
yZPu0Oy9JXgH62effaAfncqjkq4WYk1903YrHhbpoCzmzQ8pEqAN3kyudG6gwpvY
8ooIgRGI2qxGUPBJ7G2ZUKzBLaxyLjHF74cpbku4wkpeDY6uZOEzKW/Z+7RyvIJb
zRBFriZzP0jU+5QALKj0bSuylFPRLXpeKD4Wqn9pVjAg3y3APoa4CHLthCToBHQs
90BEr+mg0O4TTdYsG8br5Ap9A9Xqxpw3J68KfjFKFdmP0zafkiqN0rq7okN2ZKsC
FGQo2n3t224mEw2J8eyhuabwFE8FVjvpTzzFXNzVGyWQt20K0+Xd75CNo891G0mA
eZff0h6+lDDB3Z7zNnqy9iX1jCsOCJLigE3Lv+fJkWsr+7p+vF7kZsQB3HCqwpff
jhZak6ymiz7QnlsoAuWgR0TTY7faqmxZr1Q6HPHz0Hv5dzAKe0mQJmSG/eRZ/GMp
WNpA1Ko3AaEbgYiUd5rqhqONdX6gPidT8SOMs13LGZTgw+vHRlSnRPBgcBYAEVcQ
XNft5MGCpzUZXNyejtOevNWDVMBnL4OxVHuSf/CwcdE6OevlSh+Nitc6diHFxIRy
P5eZHRdp5SMv5SKVLYfeiHYAS365/Yao4cK8ZM2EYmt2Fax1QGJ9nPw0xTkiATKU
Y/jQhVmEN6mFLnY++rQKC3Gnn6xs8+wGLwUBCVjBZjSdRK0HqEyOJgM1FiYHwTcx
kInz/gvF8B/swHT56GJH5m7gw8xAMKHIwb8Jp7taI3EFXX7vtlT9azEoPUg1o1zv
z4hPcwFbbSnQE5N7hN8Ki/1MpdTFgQ0v5gT9OVyO5OztAQwUbFbcWUNq+Vca+Qn9
YHfB1texeSFpJQQeMDJZ8xbJ87vS2mE68Qh+gIiSeYXXDfl30qffowJ5mHR0xbOG
Av/4tY+6YnztHAySmf4Ey9EOnYj3HSQnmtcctdEwNdWOz39zgw7x6Lei8NGnBHqW
naLZssHhPKEZL43ThCI+gP2KiY9C+jOM3XkbMdsMUkur+V+zpV1GmyJd1yXAsAU+
7H9AdYbEmIR8YrgJr7GV/sCKpuervg6zuTu27OO8zFKT8VpUNu3MfN5e5TLrDbqj
KcNoI/3RuF46cbY7plHp8OVa8BqeWZTCyKHGQ6JLGW/Jsr6TX+zBcGAgL56LMU1T
s7zFwQUzKHUYaaGp/BnMdbd9fndVEEHd0SKaHD3wv2+f9HY2vNZAmsFCNyJWCFjo
PA+JSZTRrrate8YKU6q9HtCa3L8R1cGGyBb4WORmLRkshdEufouyGrDZKhlxFKXZ
DPXQ4Re9Sl0F6fsb3TbPvCLBKHWMgLuuzQ2or+VxKWE6ZFLm5O+tiDgoFTbwAUGP
DvIk/0F8SrKvKB5hIomHnv+EjquhOst9wzxAdAA98oMnhpI8GPY4z9AvETvmS58w
ueqHgl9gBxJ03k/dFpl/lyuh3/h8uzN5/Lt6xCv/GMiqm+fE2yZue3DJvhSLkWZ1
JO8EAMtPnrBpTvNwouIp/UsqaUm6dZ/jFM66SpnIQ+xmujkEITI0re4+G53Astf+
Sy58ltfWU1fHmOgwXE7RGibAEQh9jTI1L9cknOG0lNL01Vtq7Txumm+X6N4GJ6sU
T8/EV4dPCsvCz5lp2Rcl1sSXXCVbVgo8lH7eJf2qEYsiK0wEEjP03B2IlV8uainb
gM8bO9a/Gngb+X8SUIjmcG9NOppaYCKSNALT9KwUiN6CUZxQUS2yQIoskyQ8lCVe
VvXqsk4Nxdi+f8cs3sNN80HAQc9BV4kQARLFTzg5UUsxEmMXyXp8kYRymVMNlmYm
gOb6aDAprPpDWgNFc74wDl+CswpQYIPT8Ok6JCl62qvDvyDOnGBmnFsrIBm+9VQ9
LdYgU/FO1p/4bM1CQNrWOpza4cy1UZGa568nPeUFDNykCBK8QAsT3mF8CAmDPmp8
QgK3djhSkLPgh0O6nzZSOgcD4Y9kd1YbJQt41Eer5pYHo6McoKxxAmU33oMgEldP
L1OShqf/BxXviHclQBUZ6LrvjFuzkc3LXav4khsTjcu3p+DmaEnF4cBuAq6nDxNC
pTWjSsQIJX8zgGP1DV7NXak/sGoNnEyH7cTQukBfnAyiiXDJFPJbJ9NJQCqwVPJU
G1BWbKPuzUMMbXb5y98VJbYb94/HFNnN9a2VeVC4bBYNTL+a8lQQhudWWDn9hTnl
4C25VrHTdoae7aJyl/2Br1JmQbUuHXCFG068+7XzFN/OS5kxs9qoVRCePfzBi50z
D/6wF4njazSXYUhvWsT+xKxSLgLy3RNQCcxnP2iW02kC4jPPCIEV3nwG6W6//As3
U2Of4uzo18vWBmKlEh5A4dLB94gkvPTaI4SODfHJLEqaJM/LsxRkEnayi96ki0J0
lPLMFXchyNY86HJPp5ghT7JOXdyWqv/svCaHizaIShnoOrSdxldstapU+R+2mv8X
gjkfoPWrLzRlaNvo0KmTfmEFVRnVpmbMKuDxWkR9RmXVDUjlZObQR1pIamz/I/tL
g6kHKQ4PKs5eL1Vw3fJiio2APETq8meOtfgl/ZEcH7XaTWJcmUw0YgDUPXqJ3Eke
86q9kTOtEbO4hn2SQ9wBzIZDZoj80dLgDUmYxOMPm6toK+qgSUnjxniuqAg8hEmt
QR8J+qyPrL0JsrTpR+SYp+cERDfzjevAxaPGqT2N2ZEe/SKk2O4mvJJ33ksnr7ov
y+gCaidsBY5DGfrZZR0+vUnsNRY7rfBfhA34Z7f6PSo5iNq7cZV27IZ7UxxfGc3N
j8RNiSvZq4/z91HxwpyaOSyL2BmB/5wMJNA0AIeilwv0S7yBeaHiqN2gHMCCsSz5
E5U0Qm7zDitF7CoyxpS1hmwfV5Lsfw8V3yGR/1J3RWx7NGFqB4X6rfDpLp6s3yTh
BnZ+Uepsadw546vZ9GVMMrOwAkkJvKtuy+v/bldAxy9d+bqj118Uv0iF8/lKHy5k
MLgJzXS5cyqhDPSwS+q/eDB6YUS+sM58dVIAlXq/qGBLqNxK/WbEtzy/Qz80rGTD
cl5l0QAEy1OKInLf4InwlQXDv6L5xX3Ca6AJPh4D9DhfE6LWthil60aC3xttgfMT
YV5L9VRSXf1KMkmJ5PFJdRFYi29Ex6sFSDMJbB3HK74pCXQ1mKwxit53hTVRehkM
5dp1PXRq41fSDqmqr/n8i6Y5vlHcuuOABB4liUWb0GLeV8CNBWnC8PK9MAuuw1T4
6E/iYvo7ORVXwk5l3fXD6p9SYWT7NWgtld0KizvkhzYd82HFjnUK93GmO9E3Ib4T
F+cxWKK+lX8XF2CnaDgSOb6Q8aU3JMl0oqzx36JEI9k/8KN2yUyeW/DnuhVrD8Xn
mRXZofyEPWPQfMnCLB1C4UvVX02jO6DvXYDufLHMT8gGWYj6d++ag0Xt6nWjg+en
g4el0bW8BJo8hEjPavyFrA/HJZH8H+0cfw/C4wEYd86RA5N+peYCQ0qMTlklHyAn
eazNt9o99Gxri0wtvmd/01lqVVM9CrEXmP1D2MquqGz67v2rEzjRqkLSGOQSs3fU
N32JrDkCZWwFTspZtlNc2U6K53OjvUWFmQUmuA0lsPvs7fU/leMUCf0k+nh9oI9U
8hMVqIIOPr22I2Nmr8JlMhj/x3jahgS30IrpMo55JFBBDsO+3tq27Mj1l5R5+3O0
CVz2mhMDjpdOB6HUhwt7YU3s2eU2js/o3kYx88N5aMtQ1y3wDBUDxVkOov8fmeFX
Y6jYzWFXBm4KntWQJvtaAw7X+rFU52iw4NKPNbil2+S5qR7u/kcxwcrizjX26fjV
1pJDrei+R72+mGfCPaeApgFZchbvLM/8B7GXqAbOaoMGzPSgc0rTO7xArORZPrlh
eri3DY85Zt1rip2uKMVg09olwOjyj4k1NjJ+rY0CKvVnPpVg8jtEdZhXkTazsoxe
q7KtHxnWpoL+yar88ZQCjg8ImvT7jyBhqr/oLFU/pJK4497lvppum2KsK9du6+w1
i0cNd4QXIqYOq746Nff6UuSAvXss586mklN0RmjfINpohwKWUn4sDbKbAvFxNOkD
Iv9GVUnVjz4Pxe3LmDwvqyCsIJZZQ++3blbR2qj+CMCrPCNTwyH3AV6mNTlXTeaD
x7MLH6WrQ92Of37gLB6fryDYjZ7mbFqgC5tWlhK3Fqyauhy2bhMVGbe9APprF9L7
KWiufuX5S4eux1sNbeysl8fUNw8GrYixL+v30ZKPjJ5TvmV2scg6t47XLTWt053X
S41ZM9iGK4xw4FUheZc/myf20g9q0vEVQhBzgpAzkEFyRPGrXr29N3IaK4rwddop
nmKW107KKzzEAFCN8uStpWdg4oR/qVUhv0Bbz14u0KXiI9liEhVe1Csgob2IKEXG
kYCZHuyEeMXZYiV+Fm3B8K4yKhEtYJQ1fVTZLYO8J5T+nN7/VSIBboCL4Bn9NlB6
gdoDIj4hCyTgC/cvEbUP4x3/uuWopcc9b/Qw+mgDdRSMRO2hmfopKV0/kBuBLRFx
OPlW3cxY6W7XuBqm4D8rXh3WkLnWgJweMlQ/T5rwEM0UtZF45hvyVUlgpi6Rq1xm
gab+dMefc2oIt03gGWmTKv2wPZEBGBba8h8zN5y87GuLHyn/Byx4bNqxP384x467
+i5MFOIOkJ5Wp2EA3O8Kldes3eK5sawJzhad1UhPRC5qzyyNKLUcxZydkjUTOUbJ
2E7XZ+XtumJrP/jXqvP2FX9nbCa6mlN430x0Vrtf7vduMC9RG3+1fNRMSo60Cll3
VauNnQLuEZXfgQyblRzYqU3gGTSMXml0Xv+z49T+JSa5ron5fStjDXS0I0n2VPII
4k/Muj/7DS/InLfRLHto0WdGuGHPjgSVuZTtOXJ6GXiyomjynhwsheHq+9qU/E1L
lFGiDe9fleaBb2f1uwBNdcHQVav9p/3LnXqs2Xs21GplIKfvKYdTBQOO9hwCy1Os
4R/QiQLdkOt7ZIGxnMly9ViyofYFJmQnedsMIAm7r8mfNU7c/6I5eszjjpWtN1uw
qhuG7P0pRdTj5oWfS+MCti1VDzrZXZmOQI8oyjgSEhQhNL5BL0IsFGm0BjAYNsTB
8qapvzzjs5pYlqVWu3LHPMtSitG7NRGRL8l62lkxsdd7q8+wy3cwWLY2DmSCMMWZ
ytzGt5bOprZZz8cI0bxy1QxgvR5OdRd9zGHAOb3C3bnGxxzQ0gFHz7MSC8C+c91r
4zTBrK9Nkmt6mtVES8UYvIRmUcPCty+vufv/9H+3UEEtZb4yspTqj7FMbzhX9zZS
RSsTj8LDw763V8FPLXq0f1oCwDMQeUVZ/sbN6BVFwRmBQyoKAkjIrG9MlhVSj79y
43YCHjM7HHB1ExUk9vSZXYcpxMOOYrKHyjO5sHFQzKdkg04fTvBDnyzFpmEncgeM
pP6az15SiPf6EQ26VjBp859znpcNvFX8fB2ZFfB6eTo4U4ZLoAKBX/XrZpugfx2a
rYYqAbLHyt5/Un1bKT0/Pd2GvmnMDQmhtnn/KZ5Ltc6INMRt076nzuuiNHq1etbL
vWDO1xndJqDGxFwTuorGGsBbfxq3t45fUSu8p3XuRvmUn3ONKv7km2NFMnd7F5rl
6hMmXgGxgqlsZC6H4v6o5mRGyv2x495ebkrhavecOup715KSrqoWA3ps+gRFTvnS
u7TkII7AeppFHDnBVsLN+jX+5ez32kW6HQlOlUG1Gj97cNFBo/ATC9qT/kxUdJaC
YGmjtgk0ePZC4VHu80C1xs69M+m3I3JFcx9VTX3gH0S99pamJFoaAKGGYjA5m2by
Wl24e95H1mS8ZpKD0URmPFm+bXoQrQHpHx02szC+ebNZe8d2svMUOEeOcYxshYs3
CFRjtbUciRNyQ/aqWMcD9njS1EWCKpKwMUdNm3csij4gM8Paxxai00rQk4Yovz9U
3hc0elUpGJH3wnCkFBca8TxvThRsXzIuKF+J+RtMMk5jpTNb39A9IYw9M0U0aBmi
bRql2WMzW6PeGEhmO2O0ORDxS7sbb1G/g8HoNOeulH51xSBWTalk1S8mF4kpqHTU
LCiEsFsgCSBxctg0+xkPhQa2YnZB1eYh7mqWY47Nysjj+MENUvDLiTkEhUC1FrKA
5I2g3mqk7NhLwwB88heP9HJ6IKwgWFf7/7i4+eCQrQLdHlubaHLF7Iwp/y+mvn/C
IC/LWpi7z5Q4wvh94DGOo3NcSWLAm5FgsVpupq1KurDedjNL+Ej/cDOtlSlmDAhi
1ZP79SHjlCgc2Ou9aCQZa7GgktC8x+rYDkBEXApkuWhWs4xFEKibp+OLkGtdPfX2
v0DxxTEi6cV5wxoGUZA6G1a6uVCjNKQNXwZNTX4vtF5+IBuHmHPDe1smIw6aXNeB
ESovmdsbVEyM04A7UNgqEjCopAEUtTRAv+6M/Gv+YsK3z0uzqCYjfF+7Ss2vfSQN
Bv/LTGl382K0X5cqLo0dA8WOO26t2400QuHMcGe398oBV4QhGQ6CtLxob1UYgqQ7
xHtp1CbrUx/a4zGczFB7y0fZVDsWJ/1lYyPutI6zB5KzweIwMcgh8VOt0Mg5WF/5
9L3QbTdqcn6b6Sgip74RUX4L9NyHnoF644D1nWWAjDo35qBvt1yiCrrflfulKkvc
JsiGunVrTcwCHL40y4Xm1GDid0R8lB6lva2WFYh/k6N/ODx2qGkpPnHis8hXZPuo
xap2m2GlP2n+uBvlT7esEMELod9gm1Gg8niwy6+sD8jAzJb4CiPoUCsmt/Dz3ilr
ajfTMLohxVh2B3MN5oWclM+oBAgUyfS3jblDPKDz3OKH2f7TIi2IVKeFHTGhwMNX
KXLHS7JWVDT2i/VuZNHURBl2I0qE7E6OIH0cTU9r5CmkMOd4fIrvIlfa2XY8hAFV
xfNaCcJhg9yw4wLFJfmHea716zf3gSdiyD/XYQHH9P3CBKRGxhYi69X+nK3b3cmO
tdyi91BGvU1iRw7sGixWHvEs99aoXUd+fVDxeHi9yhsMmrt6rEdKtAE1XfUF3f7c
Ko6ZPMJJF97NAmungqGAfUHkVsEu6/9vmvaXkEI8/dMnSltfUpTG1VRCyX115di5
tnZ/sIMZYcOG1ZsItwOlcLnOCc4kzcLIBDX0i198qAzkaYV329s3vv+0nEzl9X8j
Gy9n3Allyk4XMcGZ3I2ja1BUvyhy0k6zJF1+cb3k/gDUpXTO2Oay80QRGOQDlh9K
JpHYXaGLVrZLm/fc1DCM4ERjFr6flzMMXRRtriMN1ZvIKQZENVbFfYOSUwHxRUxZ
fDPmpF1BMdY7wgqYpTXnUUixwJYZa2ytSW/5JS1NzMZ+cLYgVv3czN8WP7u7Mk0j
26iHw+/sbwupzsHpLy6EkevQjShuj2oA/NJplaN4SWiUqhQ4Ys1ZRSUrOp3taHlQ
TQ5/7CQgPhEvIMVuVw4z+NavZR8SMUs7pYjk4nkIVQ3zVb2JG4GyhzqPyERbGtRC
poQKluq1JkdwoZ83brdeiFqkee6MpVlTGKEm/eHzso9SAzN7SuOEfbZLZ57n2o3i
ysducA59HnwEkrbKiUY9oRvaVjwJKg9vOIBg4Ct/KSMHWRPZ+t7O1xlySQrhSO6U
37DFvaM+T0s4sBe0jfWM56UR4B6bHq/+YSzJk6GZo8a7/mkV9q/mI2kd8ahQdsOU
wjiiQMy4obz5bHNXkTeYshjYFrnhJ9Y11jlBmTu+t1dq7Hqv0awlaImHB5qzgz3u
SPFZ5LeZa2dowwWoVAb83aAYBgyCw6mdDgonpPFjgGqr4z3F/YNrrILKVYS6mv9D
Swwrgg/aPqWHPld7lU65oFnXL36Bj7mpTag4vZrFpw/TtKcHG4rVkQ6ACg15yWrF
J+qkQ/3BNfxY5KzKiHycGNmBHfWrF62MEJipnR4pKVGh2qkH9OD89atOJMO1/X18
zlgpoI82v0veGZ/f0H3cCWc9OwNKXPtPGX9ia4CZFoTwEn+Zn36l1cUMHfgJRjSy
l2GoZkyVsxclBTLNgz7yifRjQZn7bGWo2AG3EeN1LKM2I0oT7WJpVn6cpBOmPrxP
vC5OpB98xpxyh2icwIkJEotui/G3r8SvG46SXBSATAAg97YUReIiLuQ6msWVV5xB
HuemjE03U09/SCoihy9JTgobTJLVX9RLhUifXwRZT2BfpqF7aJoo1crHHfX1vm65
1C9BhmY6Uy1XpvptaEfEcJ3hZXdKN8V1magtbCc4ZpU4bypKVqA4Bf9UiZTH29sV
5nD88e11gYueO8eMw+AOrQM4LkQFIbx1MIwz3air0CDDUCGAX95KWvU3/2r56na0
qMRWoo+zdytccTOdgshxuJLMnXrJQfiDfHZDsBYvyBi+oFwa7hMDf0nqwNwzH18D
0Skc342RHrTP8tsgIlbUV7cxefSkDvS8RsVIcc/bgPNGbepoYQ5gyNcJ2oV0tKd/
E8ACQQvGE6wg3JnTgCBJ4adg4ic28epZ7j61C5Rim8ThcsnQwMKVs3nPKH1MCqL5
WKaH/2g1if78KDryJKTSmZD82wrR+a6zO1bGdNsbOj+zU/xlkD8lpShD9UYFZX4n
s34eEfCr71DRs/IW9R2No/2DsxgrbTEl307twcQVxREHORZVmv+07DRxU7XKa+O5
SqMcZ+bx//CsqIbCuWoBbPoU5OWx5t7ceHDsa0Jwcp8ZdJ4QWdh0IyOTMHa1I7/t
i0iuHbU5asCCUAdtY2vOWSqWGRMp1a4grtkW8vNV8Gpkjqws30HX5ZvZ1VQk493c
InW7hV+/BBjHDjmxjbsEYzRvWryFSBuQVrQlXmc2l9bpZrTbfold21ND4hKDawdD
xYuOZRK/OiUSlodFeT5eKJ37R+rAfLVp4qY4+Zp+2Vr+VUy0fCHZSo9/lFlkC53j
Hy8GrEc+3dGQfa+p3bon4U4WIeg0eWns7hTQAXfylQSNc19kvR7g+fZTIDlzDFKv
ebY1KRkMAFs03HTx7K+6valI/Fz3tkoE5yY1zseccjw04eOVP7uRtnua64s0KqgW
5+IxiYQzUI1AI3KfQ6FdLqmsHJVqJcFtj9g4trb4TJIV1g4IeL7uAOWO8DXRokek
yWJ0pvshiMZjV8JoU7aYFQotfHnXuuLbcMx3S8pZGGfCZUagffU9af1BbUl92VE0
ujNwDP9ih4HZl2LZ7K4R/eY0VLe0fKCcVO/Z0QIIzL0UqeXapP7MXfBcSdpsL31h
rsme3fBJLKVC0qZjmiGdgrZrkRjNMb38VFr18YiKHAP2CaTSM3Ri7QWh/Kc9ajGK
oj2HJAmpwtuDS149Wp2hvWD0fE6+JkFfxRlrPs79cTATpx4X4MVKfwPJ52HjO5nZ
UaNgUKbCFVRuFQUwK3ESWWAu+Fj7Hols3mW/SWvRh5XFsvkkYlwnVCPiTJVL9sYg
9JiweoiIUW7+QVNZsu6UvEQLHH7cxaMdaBYgcvbUn5Y3GFiOZUIkiFWa8q278ZR/
DpeuGyLyhOW9aXOi+CIISaFfUdanSpJ+XdIjRrCHYQdm8sAVw19dC6q3NhIVHor+
iAqvwyEfK6pCXCxkoR/wFL/HCE0xkS5N8Ov5f97nRLblR3pZc2hss24ECM/YYUIN
/UwWHK+o9T0PGfexDSkXP4P42nKdxlfNJ6WG8tnNReXt34Yk757GvqILa/VjdFqd
kkqq8NhnRfC3pF3Gzex6Dxs9Mz43R+v13oREjV2Ii3LP9c8zrJRsHW6Qk7a7SYd5
pc06zV8LajdEOtfrSz1ZnmR0woeS0i9ZG85AELGoLAsd0JKfPkTvEV1A/9lGenx4
9iTm+U47F7IdkpRSKMThxlHy69h1lO0atwQU0kl7SClGtWhiFca01mF0Pmq0Vi0x
JhEMm75+2HD2i1CuXQeVEpzs+1WEDl7w+Py/67R07XecfVn12OEEgy6nCP5Qq1lN
gVLUWG+5DIjqTEFHwLJ6ExQeLi+38Xst9hWZpfdAjSzYYa+QY0HwJNVWeVxGmzBV
91uGCRuGb9oEfmjiCTAsiU1cE2Kp25PUwa43VRzC0TEQteoRggHQMXHVL/DaYvWU
X080WoS01EtzHsoAqMwY3Y4aNSPhrKm6Vzq+4JbWYmwuy2HmN+FLlEvcpUDJB+UY
2QgACaTadqvalFsykN0LPUgaBxuo60BsLZw9wFkmbSvyQ3pQF4dJZAnDXRuoesib
5AGaLG/fm2xrMjz+qF+XYpheYC7UwG4bL/nS1UCgd68F6wmc/gIVBaxoZhEaV8YF
Y5jyAVdTnQKupBmsENGMFqFU415iA7IKX8ciVfZD0/wiPZl41X1lsd5jvTXamoo7
mGSo7Vk6kfnrAaoe92dDNJifnSFnJ0KScsHh5dB6JDI6tDYuhUWEYGZedLWIGd/B
8V6x+/0kz/P3ptTStgX4Ne316gP0wioWfgG08zTn64SKMszrCjpddSdf0IjlAUC2
o4oEpRfvvLNlvvFUw9rZD5FdQeiqIUvTqzS/GlwSPyAqHMH0oFNUn90VMrECNSYX
3DecPON5KztroNJllern6OJpzX8teHEZduJv0uvVDBPFNXWFCWuYfU7d/XkENq1y
wzDKsLBshdhSSSu7pG1rx52cJsxdoDNPmU0VJLszeMCF/CV+NBWBt8GEhzObUmzi
IEu6kdaFKP7Vsgw07hMKqs0wrx/9TAZVUd6bdtu5+Mr0nbkFHBH6b+Be1/pP/3uD
lBBW/1/FEPK/tVFZASU/WkXt9DSJS5KBe3lFvQtrEF3TmOtd5qqIyVWTmzxcUqzW
8ofSu8KNJjZmjSHwdvy7/I8/7ShRUG6xbeVs4ZE1LGK10joHgjCgOD41bzpuOYWW
MzMnnQgx+CiJFQgRLpqdNR+Ff4wP6Sm1zFbXfdhjmuhohDihjs3eHuhTe1yac1MK
PtvnFrG+5/haPS0LHoMuawFMZtfHbR7Ct+bkQL0z5LEzNfXFjABRrsTevzJUhh0+
I1chwKMgrP2y6A6MsYk07ZQeb0F9f/xdyF2eRIxriP2Z+wDmUzA8ir5Az0KkAJ13
4MOyupmvgFhwUaBfxcXtd+txN3m/9tZkPCR79aUqME5b8Av0M1casUp/djZmmUWA
SgvjfYqmQ5yQIvGIwtvFIcQbuytlGMYwWzrRbbDK8sA8hUIQAYlhoIA8mZA9YEkL
3W7E6zfK+CE3L662prAqb4PuoNtiaR22buBgD7MyzlOmCw4EyAg6upE8S+/qjM/W
eTh/6epP6IqqJcLE7siONSd9za+mGLANiLXBivt5HBbZDJhdmDqiMXuFlLtv0Dva
4TDo/r41u1UqGQLB/48WU5aQN+KNCyFPlVfpR9GKXpvtxbNU1m563NPkh2t/NH6J
nhozqQw7hxwpsiLz1wlpZKfOCsMtwh38W+/kj1Tenlco/pRLZdeyWDZqsEPIJ9Rk
ssVHKbnZt5D3i7+s8ZEN+wtIKtbxpZYHZ2ZjTvFnwJwA5JUQY6arGCvbc1GgMLNL
WdgHpQi4l1ON4z7QmPDQ/IrdM1u6WGUqMxqY6phmR5sdKTQ47aaR44NqsLrpBOje
bC7BMEiV8GSev8U/hJX6u0L+8YnXVBbW7Gb+p17vscTszh/SLIW3U5C/s+Qom8vm
s5hv5mPr026kphtGJ8nbXR0pnXyiX2DTGA8IMPEarmMLYFSYOJvwrRwPfeWnyiUM
5xrw1dMuVWJeS4Howol0ICb2WmkBtM+tMJCvA45/ceFlv4ExjhVCgDtQW45g14We
bxK5AmsSduhtr+lkb6RTIqGFyETFG+/f9ReZe3jgD/RkAW5ZNGBXUPZbrGr4DiMJ
PWYpHtIub1QLzZFidId9CHexIwxcuP0bZ7F1cablPGG4NQEWhgUPSPou9o6prGOQ
4nzN/D5Qh11nUhKvUR27Y0uwW3xfJJIMylCXKt8TutWYHg+r7MnSGa9LRxT0aPCz
rdq6t7MCA8fg1xLtDKfVuJZFqXP0wNRHqxDZY8igOixjKpfTh6xAPke7Pce3vDeR
YHx2TdqOoyhVLpUjCbpdyRvJK0/ZeQefda46FVv1QMc12089vjWUEO1Dnaj1i13F
tnbizgVU1pCh5dW1ZGFotjWQ4Ap3rHL3DFaW8/WiH1++heaSw8WS4PExI8TAftCX
Uv8zfX+tsGVNDQXqGcf1eZvLiEHyj63sQh7/z9rQWv1ERQeU531Rlq6Vak00thzB
VK6COBBhWKyCy3HsbAZ0ULXZ1UOJplxj/puQaMDEHKV4M6rJ17M7V540wfoLYY2U
B3O3Xnt0oXfJ0f++F1X4XTUVShrCg1iVgygL+XfyEIntOLU6DtmuZfFzbYsw2C+N
Bkrbx6jTR+EdZgD4FlBiwgG6xTVg3ErLQNubKZxbak+vVJEteJa/UyhFYV7f6NUS
1HMsTTmt46uZd1W+snplJJHxVc1l11tczUORzR1qzqnxBhMmAJg9O/zjwqHP1ut0
69FsycuCXtgCB3biHN39s4qV5/FdrnZ2BpiJIzZJPLlFaF+tjF19ApUUxZ2xmw1V
rQpHBBvBwlblNThnuH0qNl7Y/pkc/qjqVcuqUb7u5mycvDWxrXuA6knmZSCxN2W+
Jp4JfvEGmmBV7dmtiXR9T6882U3OKAxPN6oPdMUyFj/SeJd85bZWbW5YHh/nUQd2
Sn0AHtyJ70EpRsyHdCGRlvyDhyOztNjmdu/uGEytkuJOmm07qC/VWItf8gxheE99
LrQi7JJUSOBgnVdEXw4+GpQr199W4GyGU/NdSYFGCvbXXBkQ+jNkCHlIndMPkBSg
ZYg1zZ141azcl3aUkkXPkaqXr1CJcpR7rL5uDhEJkxDGvGSRFGYiz2gUZ9r4UxvX
k30AcAEZZyyOpTbeggVimZzi2+RnxXuBkYy/0EgS/tk9GxI4Vtx79Vpk/4ZXXSrA
pyGOwTpcX0ad12j4vtg7HxpHPT++p+JTSe+IMoTYWnDycVWKgpx5We9fQT6nPIzi
/pHFkWK+mMXHPlEZkiVYla4jUEDpGxbiZV94iZuYciBT6eTPh3q0jNV43xtZf5ok
Qoz9K/WAxKC0zqtEU4gCDcDbhtbtpNi9xdqQ3Lh8rt/Uf9NaEprQy0xDaoUC5IHO
g6JN4QElENf5K6z8xbRlegav2FGcSUqx38km6kBqCzSlce+PEVWAbfeRpLGQtAVW
pL171UFGe4U66ZLAHtXSheqnk6k8qUiaLDVnTcJq5cmM0YOBzskSsW8ZrgLBfpY1
L76SVg3yFAb76HNjGenKozP9n9kwT4x6uGosrMN2FDwPqepl+NVf9Xi1SZY9HWUi
ytpGpago6n9Rlnsj5/jKPLyJkhFCZDLysP/bm5zK7+GoqR17scejTrBSccNpPLhF
J6VumBDtRFkO+8R5ZasH6TqUTHWQKhf/Y9DVscWohgWNP0LeETpqMs8c6MfsuHO4
qcoE7qAru5L9v6257x7Shi+zGE/1WqGUpssVQpi2JGwDKqKIJfBrQ1Ww4DBW259e
`pragma protect end_protected

// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
bhSmlFN2r7uqGOLtUFQBK/0fFNJR+cVzrwftpEFbAbbFg7xbc0IZyfzf9OgZ6Vmxdy8w7U8VKhlu
aBAnzLsS1x/mWwznRTtKMh/R+7VUD0c1MXO9RQZUUABTG+JwLkRrmXPfsGNec/vrWzrizPGSEyyd
MXVLRSthflhzu5+5dWrrvZ5Th1w2+4U4ZfGd0UERaZBFD1x1vVrABSz4KGU36aOOqAlN3d/tGRcH
ZfGwvcU1v/ZHF7YlgKR/BpAjxHqExjJuTqUNNl+o4cGhm0QeytvmTVqxnAuWRiCx7jaQutTL0Oir
pq7iuGo681w02ab7/88PCpWc6ayurmcvqJm2Aw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
qZGA5Hrw/m4BpvtFgiaLQ6s9iCsTwK08Ste1NmrKi9l1ADFdDihDFGRkQlUXgPQLX8eB3awUKDGZ
bsMoj0pZLEZ4E/H+SsrxHmyqnzZJZkODNwxOsXGni9ZcaIPY2iqG9bLSjGCdcZ5Te1jdo+tD+pAV
GqXCEedZqM7S1YjAphwo+uekSOsJ0vVlMk2fQzEH87groDaMajQFQhvlohBpWx6H7b4kGG+u0cvg
jpTi3lo+FjJ1ZiREGqBnC9tRA7/pgmAafxCAca67kXqeopHjNIzIT+GlQm0h2wCbll/9LzWP4xPp
UbLj2fsEVjVZ33Gi7r2aMR920fXJv+C0KEgzWAE5LOB2tLWm1YmKKTDBbSBFlQN4HT2stC0NPEir
JuyFBC78V9sqEGj+Sphrd9iFIVNvEzSDMu6BvuEHTS0QHfhqLBakQtmCsG9dFbNExQMthmKFA0pq
2MSi2nfIjvDkn93DVozZP3uzVPBEahH3MQB97F+U5KIlyR3Ddb4Z7FjAYH3UdAp3AobSBk6ylyDj
yR0iY0eXreNVgb79TMM+kMqRwWmbHEoDlsxnbZnucOgm1Dl35nFcCX+69bLpF9vpW5NkywKdxXyi
60i9BSQvd/IuT0sKvHcIfn9jRWMrQB8wliJxgeqpxaWsND41G6vsj+vQd6PYP9EP2xJPKY9QopvG
sKq39uw+2FNgcFF/xStLYkwX5AAGFq4OOZwmU/zYXg8D5HBGM60MFE3r7wOoTYLoXcSteOGjk5aL
4cwhLUZhVpGiUBqMF0LRQt7esmBHIbXYYxhPM7Dlt+qaO+Sk5k+vA+FTG2M8EX6G/YcnwOlQoJ7/
LV13yL6vmV0syPnjVjdbNpMoZynA+M1N7q1+TxHucVOppA1x9nZTZ0P9YZPzF35uq5xcuMN2bFxy
/koV1WWCIl6b9CseqYoguj3LCV2LlFPSP00iLmBBpdk9uWw9ljFcCkRyN8/4ZwYFp3Msyu6wJP4M
q/dSWl6TuvqT3WO2medFIGlQTZM6iQC8qw3aU9nrlTMCvSFyvxagsUDMsUYLHEEYaTJkhbJ/RING
jn+WOBbIeq/UoofuSfriLAS3mVduIQaney8eqe7fm8Kf5OAWW//KrDg/q63bS67CzPqxEdFNJZpq
hT8HX74y58OwLWUANDc2/Nhhyg5VK0DxHdWouHAtd6RnR6xPSnTpynWo7ozBKH0a1/O5veVDPn3j
zP2+g6W4qCxyjXFNJlLRSkt12FAVDXrv5I3AzG1SA+mwEE1RT76MFQ80SyiLjJvpGadnFtJcZG3w
qFql6v7utyKEmj/HWXUmh0xzQIG5DoIpZ0dru4gSJVx7Byo6m4udmqxz6GqLRyOrXMwlAy+Hz+Y5
nbouLR1b4MjKZm+Rq3yPCdA36ddnayUZN9QRjTivE+rz7W42oVkQ6q4rSYk85Qrl0LQ2frgC06Ws
xNcaYBQjGkmo6Pumi9kFLYHT2aIMBmwcF8uuWZ9WwION+/AXHcn+lAd0HOZMbtDKggeaI+y7I2DL
dadD7O+79juinffzjFAkrIrBhDyuX3x+g2YJO2TOKtHDX/0u6RWF0Bx8pq5V492bNiJdsjsJp2tr
R5DxFbr00Gn0USjOJbyM+Y37R3GdjLakhR1lIQ4u/T+TkPu4CMIm4HXfVoXItPOYu3SEpTC6gEWS
4xtxrK/vo8Ep6Tzfd8bxTa9XGhBXrzqK3vIlEW+oIvZE4s3SYO/1uveziEbt6nSdPzQUeRn//hsX
fSh3JLBY2PQU7uJ8aWdGV203TJqo0ZjEG/GM2r8foU2zDUAP6bXM8jGzN4KZWhyk3sqaLS4hG7NE
uEs8LdIdWxKPCbdEqnNiHgEvSH6qgxG3qKRjWkreqr+5Hc+f1OV+2jAga61ZOzrxnVHP31ZQxIbY
/QGllcyQIte6YGQ7V5LnSeaGev1rnAwMpYcUQTAfbgtyGS2ZhyjytYC0H+5GB3BxozhU7ch2Q7Ym
oBiUgjXccljHdcr0YfWvYyKAz4paZjBtJj5w2XfLbwfttNrE/g6tR9W8nXfdxwza6Ri17IDyB593
RavAxKbjN6eE+lHG9GbAEEwVkmztAwaphMF9e9cMKXQpOsbC0If+OqD1Ukci4Xy0yM9MlAzGwAlU
VFNNVTXYjOtyYqTRCbb/1gCNe6qSa/GMuMPkmnCRB1DiiQ5rCYJ8I16bpbihACXu9uhLRv6bDqPu
zwJ2RF2T0ZsNUr7VMt0WCefkDp7irh2EUkKCFhXZ9HhdQXNrihhCn0SnK/XVovJ3tAXkel4xeQiE
OC4NXnAQA/jH2S1AIVuUoIkAobXhsi2z4FWPPJvbJeSZD9U69bnejFDOCYVV4PIgo1okTr/7gsFG
xw1rPnkMp+1dJymDzygTHsY24qBRtJ8cgHbndKVN4e9DXYqg34jL52SdRevW549PH9B2sLYWGaq0
LVfYtdjcA4HBpUTpk0aEc0NLfGdWAozVp4fGDWGpiuDlAOPKSt2nAcHTAOsqo9mtQ/ViQ40RihMx
0nLBuxyYfzmjz4BKPoVNqxSZ3zHkovfT2aaGobnicVkVLWdXM2JTlnKXC67mp7AXG7G+aYrhoX3m
bauhyXRb/UW0hLslnUXEv5pxs+6O8RMDFFiPzJlGDpQaT5ZyTDMbslepreF4bzUl6aVoBsolYBDx
UjSdnP7nRtnYFtdN+/yX/It9WHwtlKafcLcQYLMDOF5BCnqv3uT3PL0mO1JoSPa5VdMYPa7rGuEF
upktl6UDgopKFoTpv7i66SyXVUVEosJIzk27Y6+G6LObdyEMzc1DFk1iIjFAM8KTQOl2uULiymbQ
drj4/DmH/7P0A3GqPOwPJ6RZVgAXmhsUmHQVehq6mJo4P2yA8n4hHT4EOj0XnG4Fd7e88bxSND7J
I2cJEgPNltCd9WQq6Ic64EgGtMk7Ix8JeSYBVQM4o7GgkIkV7KvrIaljBdwu4QJ27m9Pfplp6TYK
is8F69VcdID9vn5gbWTWZ0nlwGB5IFiVo2v1+WvbGGGZPJzMArAYlJ/PUjOl9pv3p3Mx2bzCmeyO
qTYymnAB99MHvY41Z3HrfsIftcRLnM3Yo2+bdNTrcvgFTnJ8cHsaXHLECnr9/IJeHBA3ysJbK8PA
xFM/w8UqOnZYEEq6drozyHqpzzRqWYonZg7oRtnYTiYUhvWWs3YNSvRbMsflE1dnCecx92UkSvw7
lj5OdPZuP107vneGNFLJ8BP5WavMY8zTZVFI1BwpfG3bxNV1Hh83A6Fw8VKW4acPmnwRatngk9JB
WGmkkRckaGvArXJOUOewx21hUjEk1rJW+SUQhDFJ2tSgKpw3ivPX/+swyRTpYBCpMIT5ihosP4it
K3viV95CRynPbQb+ZR6sVDyqcro1AHV7+daCbn9wHzF+SQaVCpiPBCGk3UaNWk6Iu8fY5eMHQ2tq
O+Y+7cVPAx8DXSAmnNexEtQpwHh1MhiVfdidsBYbwVn86ahja8Ht5gZVa15CmOQ9fR6uYSve6yRW
EItf5CLiy/U0iQfHXYfB7jtlaIn/vauX41iDJO2UocANo2wCPt0BFv/MzrKKiW29ryw9jp+Czj5N
N3MikpbLoIDQ8ZQ9dljbvwWooD3f5cEP1XPjhyYG7e57RD+b4l4BUJSESrqeuFr9lcUFambX9IEI
uSWg5evFZGlgj4226V7Ct7V7sRsQyNSu38gkyycuQbmDPC3bZNPyn8z1HJQeeLTYltT+89bHulz2
Oo3ORafBx0WGczk4nCH+BBB5vcyQGEjWZeHgiEVpXwMOMXJ/52zVsVhuGmrZx3/YffEYmaeSFBeb
aYIST9q3IzQMYEVN6KqrYXWzp+a1NThQqVjZlfVVWkK32hEexDESFcCrz0afz3U/Xy0VWdEzR8cd
Nx+nj0v79g5y3Xto9LINUTAQWtLfMxZ+b8DnfgPnh5xLapySkaajKD+ZeBvDPIKDNP6QRs3x35eH
9n5KcJaMh30rTU06mA/YyQo1PyxSo0uyGORMvYu59LP9fUhThVQs2+U8SdkjPBEvxfBbhDYfQZBZ
+hbzAF0q+Rbl6BSs70FKT+BIhRf2Kj5oNdFuLm/6mKDLeJ2J7/qmtUqYv3FKZVr2msod2kZnB5gK
GP7V+oLAVbnfOZBXPq4J+nDiPx6q2I6QGMokV5MTgn52C1BAFnBxXPJgcbFR1g79qNWXqDNDLeqT
ZphVdix93I+kwjmCfupCId/1QCPERGCrs/8uFw0TbRAP6I3kJ3+UFpLSn82IOfQpgRpNAibmKzg0
+yWiKDxATX2rDVtMiQSoX9Yp5nZAwh4e+BudBV6eJCvLxNeBqgJo/gadm/c6NMCJj223c2dQOGsq
nCqbKZrVZ7rpcbQIlxSHRslwYnytrTEVAUzKadvmdnZ5SeibeblmfmAqjmC1KLjnWHHRLW1ysnUH
b4bAa/ts/6yqSW1+HWiE65MLm7ykJJY0ylhT2637cVPqFw99lOsVxLSSE6vIZWlJW39FxFSBpiPs
9GcfwmsFq6NqOpBvn3gllDfs4oQfbADQhAPytRqP3Az0PUdgwSmHFBlE4bJOGCW1hlzuJ91DT+YT
pyks7ZVEtvA7eVkA84k5fBxTmXDOpLJcobo/TnxWkSqPYZDaqO1PAQSQGp1l7ova1Azv/EEdwIja
1u55yX6rqp7VF5CQ547k28XjH/cDC8r+kCDeEyFOPzVj+xqcdWvPGMbhR2RRZdG/i13MT674coJR
8jUSUNfAMvvdOl0w1kRA3kqlWjbQsY4BB/a5OZJ54S8wn9ylA7AojTRJlTX7QxTpkVCYvpalJXZr
doBV3j4NFQ8fwIl3Ru0iYHTh56gF9a0zI8nCTkb4OvDfPklAiZE8l465b2S1L6u7ri351nw3KrKj
fA557sqMLCOruUSUZP3JGNjI2HIfrJHStfcgWmJWJve3O+m6+FPsbd1CNh4o/sr0w4bYC1295QHQ
1kdqF/WB5a1ZORxNBwngq3382cUaCSdOsL/Rb7FzTyrrgM40RfJnK0gVtw7xNGvOJDTmhV1PF7nJ
epTxdJSwSfCQPerlostDDlNyG8KBgx+isaYt2uvegf7nHPk8lsuRsscAnKq6nv1pGyVuG2w7uhVW
GY2kk2muCdanrmR16/oAVG+OzqtW9Xy17uXcdl7rs3O4Uv+0DldmlDwz9ppOyr7tsjWernKT6Brw
+S/nyA+95rRHPhabhaUxWx1JZ1OXBsAFtpEzlFOEYabcFL2u6K/Pvgs9aptC4ESyfV8xTCIsVS06
ss2oppnk+0JXYMjjz8X9CG1uSUtTvKBp/vx4o/G/W0NtdEomrx7VuuKefvhLaoaZGmS0shA/taPy
dWnJXCqR8Okdf2kU6aTFwTfbO1rWnkkSzz4TYIdm37yXxlLpwhDgoMngci9et5z/kwXJPP6rZjEV
UonDRRXYJY4eTimdKKDm3nP0LJKpyKI4TtrK7FOSUV13tqzev/EithW+UYn01WCNTdNss9cY8OOo
4RmAhtlePSCp9iXUYsQOVAvyTtDnv5OICVRtKo0sQsfggDitlPZ9iB4+H111Ivh6GtVKx2AC24mQ
aNtCEwuPTvGJwJHeoQOzONVLG1TGW0/gPaHsMIGWmfKqfm8bwsXyFf7IAVHs9POUpb3aFb6otjH2
9LBGBTPiHoc96IlYsKvX5RWn5HDAmCWZc9q042iHtRrcHUXKPkhhkxwr4HyXGDFoeuoqYkvoWRjg
GJFhuaaxH9Y2KWchIIi5OXs+G/BJUs8Pd4odjnzEru+M4HJiZcaIPQEDBHSldyyYFLWkxD14oQFo
YjTsqNFmpU7oQ5vMsB8YT6yxZ61d+Lhw+d0AAuAqEEGX6dJLOMsCibReXjrK6czb3/3TDEFOJoyk
PIXNMPb7+m8dHp/AjJy9sEFSNsJ3bV492RcVs3gkLLYvRJj+dN4zuhYtmnjp8tuIVNjWCrAzI1YV
U1JyGIHHqeLOkqG78b1T8+S8uYt2PC03GbjQqRIVa5mNek9VFx3WbRMnL9iAUNQY1vRnHz4fNbER
mi+46oSxMZ5Ij7QfhiSnfl3jB4mQ9sfcnFpMnbH8fPOXIkhfHaq31lak363rI+su1jdGhv7xpMWk
DMAXGbh56+j1MpVz8pPdAO1OfC2Fi/cg+ecN6z4Vr+J/aHFxG7xeXxnDkaIyK/QbtqbZ5Q8sW/qj
1ens9PU4x7ZqkFVPEC9uQAe3Fvcg3kNoLnZks3iNpMLnGmLrKQ2CIbKmdV4gStXF9k70rVoBx+My
CNidVeqnWRWgF8d6hrfTEc6izWWrp9QV8LTNy0Gm/uz3+osVxragNRitUVx1KQJBh4Xuns/i+KJp
39b2hiTvTFlsGFmFQXZIIxC9JkQ4oVZG0QvJoxLYBuPQ2ibWerZ5bMvM9wCFrF5h4phez6NEVj+S
1m1TEwbacnv7RS/1bc5uY5RuVQvf//TNthyTOnUkKLZUh3sm2GrLo9nmv7X+bI7PDeDm5XF5tZt7
n6taauM9+I1Bk+EjrXy9296bYAhcKquMH7Ckko853QFrjVkKkomqzOcM1Hp4RALK0kcVgKhrBZmD
RKbZ4wCYlnpojE2ZpU/48krY2ejvQFA79DFF3Eb34r/mLMI5yC3QcCcwVtwRKHfawBk9RbKXjghR
fL8juqIGuS4LeKQCrykIH+y3z/0qk7tCMgO2xWk6MecAIqftmhuoAtQgpjJYDp/Ng1kmj/Ywm0fb
f2oLwuqz/EGJns/U09pSVNy3XeXWUdrPxg8jDrRGUQY5pG930LgEI6hajytBk3Asc9ITzf3mxLCz
k7u6/MK6+iEADJTFbb0KnaX82hui9nPwB0YsVCsolreuxbN9bZBAr+ruqX2a8P8bCz2OJZ9Ufqjp
aE+n1yMAR1e/PbJzEPEBUve6eOLwjxkCpd3SJz1LYsP2xMzUZdrSxTiEgN8RAnadjMEm+3JXW8ez
7wQYkImQlXeEt4HP6gtpbba1B9mac/fKj9rmmRoVKWJ89n4f8Jwoydc86IP5SuNZJGy17nrXEFrg
gCzCiz7EBhKUU3ENLYL3/nJvG9zVJvriZPJyvJ72B743gQy/IyW9SYoZx0yfDp3wXAt4DdenVcyz
ytk0EjGnbUP2cicIgxeNVLdPzyXbKdfF+oSrk6wchgK3o7nq3MC9VOTSZXUETaZJ6FxWKmY8/HCS
WF6cIio0tf+4r3izXiwpXWAUgUOhP6H4kzfZSpaOEXa3dioKL55lgIQOCLJxXJJoKF3Y9ADzM828
VZ0TDdAJOlojXUlWzorDzrZOt7I8PNxvXqd7YVhybMdca53Q6fdyHQJRVUmZZMUIghGePQbJXjk/
3ek45AM5lTjRbqUUe+tvyrQKXqF9Lm/8xGFDd2SmTDvHQGWQ4A6uMT162EYE46RbvuvL8F99J1dd
OQaTnZiEBsKgrAR2xRtOY5907xYDfOTTRHD6CZ3VkYlrIFMN294HHlM8EkwKhT9zcJLtv7Cb7Qp7
h9axzPF0P+VpMSyFPhmoUgxMEASrA9nDufUlzm39EWGX3J9kOIDHDo7uTej4x93gO9g0BSyl76OD
Pi5C2P3C8FpuH6gwk3q5Glzh5uWbVudT0vY70khqzRG5Utbb8fr+GxIxIjp9xaucdVs2BG/EVDol
6t3t3bkqQj7vft0uD93oTonOJcbk6gbmHlybodrPCGqr2PwRkOcOM5F3Ftt7zWg/zbDjuPAKcmXf
45RWpy5Js5dHQZUzeT8WBmQJpB3YCp678aCEmA+14WGKkiJoL8WY21+BJFGQDHSsmQ8lKo3udikB
Im/ywjE2u+CSbE5sVUSxKUKTnb1TD+4HwKuCmGtaZe+Vyat8wvcc2oxvUaKGNE6NvSSVVwM4wdRg
X0lIm93ARG79N2YhC8OfvmX+Vi6RT1UuY560GrgUT7YiSUOg0oGrROaEwnmqgZxlniMjEvavwRL1
rx9NbxWF2e92+oveTZQGh81mq1+9reDzS3UbDkq7pWP18VwgTovGfM/gdfqUuqTnejdfwyHqmEoq
YLi0hTzjM9tUs4wyunKeWSuDTveDESIt1NCV4WOG5SEZ3lfaMj59jpluFsfsRNplgV2uT6N75GY9
eO1rzehCz/hGkMM2qUATMyISzXhhzxQgeDyAjL82l5XuloWdDnRpsLpZqhZJ0YDQ0zGRtHVK1TvU
pht8sX7Z4CFJKcze3BroAvhBqY2n4ZfODut0pWlX3/o8K6MWVKr6OdmghNqRrwm50V9h+8YJSH3T
nru2qkJSUoy/g9KLItKq2pVxYw6cxE3LQxf9x2xzj6h9dS981aj5YICzSe8Ps2SNu1nXNfEfpDgN
QFxlYrReqbgCvOcpL4BQZQ8r7Iq/cWcqau4l+o2+9O0DxjPvohqZVHlHU7GA4HCSLzWI+Wu4Pl2o
/0Gr0kOuJk/3VcjvZOh1WYn54Z/9ra/tGuHMc4I8fj7EcpvQIBCP5Uin4SV9Awf1g/ki2iCfTJ1S
p4jCC9hFl8D4fFMXAhvzhj5rGvfBY1/lQsyXSG+bJfveUBr4ibsiKuiUhll3SsM62uZ9DiEYZ4+r
s4npZ8O+dKrqSX7XjDo03sgPI7boVvo3FSAQMNAUk55qeGjX9SuNj3QSDd+YF9MzCx+2r6QcUY1Z
6Slbgd7r5rbIZpcIxCmV/1XtTLf5SBKBt/p/XVRmdDBsTUPCjrY5QLc/hOHZXVPFyg1SCKFAjpl4
jN/LLa0XnTgR68jaTYX6OrDvcNjNNnI/y67LxpJvwCtWQ+YKxkXVmNMCxJEavM1uI0jvQcI44YbZ
nP1V7Os6EQxAT2KSL4YvgHxKYkRxGddf3nYG5lHiSQ5tCujW4aDTH1SJitGNabfVcjxoTnLV6C1A
pJAQlOleOqoqnLy1c1zrvQ6cwH1AaYXkLpm1YuahjwO7NFL56f/3NQYPxwoGXYf8B2p0IJYC2DLT
AKcKnTd5xRZ6aZtRfsmmP72xvGtY2IRS6zpHd93SMEKid/kInSnHFWki6ZyrGUQ31IggsVsvAfmi
D6bgqG73M9yznBf0dsOcvgvy3EvcqYOQWk6Y0QkNLSOEkt9dwKjuO8HWkI9wOZjvwd/ot0m+Pitr
eFgb9g9EIfRATVDasTwihRX25MYQiKpmswioIwpf5Bm7LA8eRvA/YSgFCrLy+KXkryAftkC/gtyU
A0kareAOImMbJ4mDR6x6tkeJYBSBnEjeKPk9hy53qQEN1ixRgd+AJ/thX3RJs7cHEnxkRS2fGftG
qOFroiX6XD/BPOHRUPZF30sb2IpqE8QBwyWjandobV96Q0aHIbR11ikBIWT02LdWnIYeavDTwaND
y01bJeOR0JD9XLC5AKRVAMp7UqEdR78uZSIGVL4we3hfWV+R0cHGIQEIl+3gY3tD63ODWFjkxPlQ
ediya4x6kSyLf7nzNzUW94k8gPi1zqCUjHWKfUA7MMPjdJnuok5Mvr4f0rqzJNbE3r7/j4SdZ0sc
6bjEmLY/IEO7upOwzfGNsll+MwZsr7pTGnB2mJJlJAG8KLsR+zsQFi4Nj8fT77TOWfHMCokYJYYd
iPFQLfwqUmmmkLbKXRg3rKE5PK/T6vduZNNiaX6jZt1X1f1jXWJCACMOy4ynCopdkoRaqsIUIAxV
/LnYLHYmOZtP1Ux6Mom5PuYp8yK9O2n36AoljeaYJF8bUxi9h/RgF5iHXm0gysWVsiB2WE2ySs6z
jnlteu+NfPUxxbXnI7lCvfUEbRwD1IJX4tLuj+7bMT2FT9oclxePDgbJIxj/cR/ixEdO14kjHyuz
hKQXvcPlRWcfjiPKs5VW+z5acY+CIKdBjaX8mFGpwLEzGA+2S1EDBoSZ4EXLVDuMs3VuavIbWSn4
jTE8ZYgT5TWveUje6z01ITPD8jThxLt3R8LFPaY0FkG6eDvko+JMYiIdHvBVx2tijat+ahkr1suS
4jTKEDwPoKfpZPLWRUJMbjXB38CENDKASOj2HXr8+kZiWZ71i/aZqzVUTi+e6HmLyP9JsshDbIJ8
qq2pCfxVb96jGxIujtb92bDQyQK6J7yee+qHPfevAUnjjrN1SvS5WMmG4AOcy2CDX3HsfueU05SQ
PhgepmvHb96CU1k74YgwlRtS+O9VDaS1DWyvy/aB/wLdpJ1azclojIvQsX3lcc8x8B8CtoBPnB9V
35hie/5XWWWXGP07bIDDWxV8c0KpvX85s2Q1ewRdlfYbTFaNimI03ZNRDWVk0eSNtFCTEHILakWK
uHgZAl8wTVEs+TxI6beJSF6FF7aMWDBs3K4vOnw2D+e0wPPF6Aoe9d+Wv6aJcEpqPnhWZGL2spCI
/smlVZDDcP9jJOhLXon110TnsGyM4umfbt+lCICzsPXg7TNPzOy/3uxBM63S0V12mj0MpPPTvjfD
P3rnYxhVT5VgFYd0nqY4RAZ0oN7YpG/t6CHFQCjoGaawtC70GzA/7K//+Z6ukx/mQgUrypmuLnoN
jjQikk/n6sQJlV0o5dr8e7xzRVQkwgACK2e2Dw3GM8ksEnVL8mCsadekwNhw5EXW4WmL83dFG9xL
lsIkljEyU76de9VB4MZSf+tFaP8YQuNwMxrg36lWRqSKDuTvmYSOPBonpAujhz2yVTXp2miCmDMC
QAsHR4mW1nhQ/WsWHrg3OHW2BNz+gUkHpb+XercaPc4jz3wTW1YMp48jcucRWd7KGN6+8cIo49Bb
weS68Snlxzlix2oCDQ7I2d/sMu8htfMdgCupde3S8J0N8zkInpzSvOHbD1cnmPzLhzbmzT4T6fXW
AlI7QJJ9jxVPxdWQrlPBo3R80lf/022mDGb9ZijWzJrkrv+d3GK3jwhUh0+o0WqeaaGcD2fnCsO3
FwURNInVEcpXuD1p8V/yUvSCbNEX96sQ9eygCrEgyJ6ZFFdfyCF1I6YsNysEWJaTJIDZ/vhSFxYy
daz6Hv4qC7t2xLCFl2mz4w+OTy6/XVWrBhii2wf3O05elNNIkHtaB2sb+VIl2lkbY7ZjRx26mY+Q
YRX20KKdHztjKR4MidJ2JwlblMcT1IVL4IT17wX6SIVIQeG2ir4hD0raZSOIBntJd4I1Am0mW/dR
mHzpctUu+VShajEk8UX9BX9MyB0Rq1jxTvGQ6rvRPBE0VpbFgFp5KuFmybU7N9KejbtVIvP+vyAv
mpNyEiQ9mSLNVi567b/AFrfMLFaJXk6QTTiFwoP0oZ5CXAKGv6O+3RHyeUJhDX49MJtaHLBzniUf
x8tEFnvkwft/FsQRNdw3bVjRM38NmgQOpZXiVAbYzm1/AGp9WkPs9urA4vISDiWKBo8ELmWKvn0R
jHlQvLtvP7yMYhfo/1soZ7vb/F5sYyURJKPuub9yGfWrk3H5X+tS23KYs21yETR14FdQiLfyl5Oq
+Umt8p02oWsQwo0MVnSEb6tvJ/ozINTfCArNJnuSmBuDM1Rft1nOtzvVDA8bTweXaQYH43O9sWb+
wpMs/wc5gjDU5bcqeN0kYSOQl41sckS8I2X7v5WXNO1EcrsE66Si0u5GAUzYv5Uk3vcWQId7XAXs
DLs5PwdWmsH2yAqDsefmDdm1bjYEPgOhbrfFpc5HqgOfx1/nblbTt7qXfcnO+CeEokgOu3QZTIcK
QErKs7F3KOpLI/ptntOyubUIa0/RUCPHKBpKU5RxIQGmIj9hyXsBP7au+grCc03GE3R2LMSypJhA
WzJx9LU5gpsVgaAv+EFsMPP5sXXtMZu/dp0s45y033PrN7qQuemnY2umAk3m+A2YdxZCMBnsyLZG
qIgPTpz+2BoN++4G2SLlPTww2N7AWz9vaiMAgUAdN9iDFYXmfxg7JB6sfa8KzVMnLfV9ZWipTJ0U
xKS6zKANtf0cHjh1chyZfb8nVtAHTXoeUcS5Tk+DP/VZ/CrSff8/J97o+GHpDrLf57uN39BXgrLX
0PfbM1RAcy+ie6nt8gXpCbJndZxJmQ5sahAvVWRp1tsREzLvnKHGW77sKSTQ4t8M2Pm+zaiyX07C
Xa6qwm9ltIADkJfprjo9dBvTUw54O2c2VSH6LILEKE72unNuP9CMHmw/XGbae1BRJ71PSfH4Ut/f
b6XrsR5LR1EjU4rH9Zfa2wFtid6agIGT249lrwhA8oCfrLSlJ4EPzhNlWCYlo34kiY2IKN01PDtE
g5g+MI5jrH2IYTGUIhgUgun+WWkyRnj2LPPWbM7bBGMQUgAc1Nl9VoEDP7epnlyCH1knas4RJluG
COyrMnxxI78tSyEEUnd8XN8xjzOaSljfTP0b9Y2xHprTqa7xR+NtEMrxHfISQk5v5l7Sw8lJ+hOJ
4gtV0dXAsq3/LCje3x187ZwHldyNYQUkBHxNrWGFxM8M4B7k7iQiGyYugCrwOUvjI3+TfHPwSb96
QbUYSlfWLb7DeRkzGFl6j9+60OyFeIi+diamop2Zpy0UrLsukJCZfe52y63SELsU+siHNzn0i8Q2
wDA0hInMMZ66mnR8aHT884XWULmwEh7JyHQjQR5ewbwkScAA7/RMBuOksNktFh/0cBO9ZaoxJKqF
KfUZADwExntJAg+G4fsdL9qC0G9vQoBI6hvPnK9EjTExyDmTVXpVuy48mEQA7dtVd+zna81+2hC3
KZ51Yu5z+GmYgPveUdEWY4kBOqsL6+2POJFay93V7e+d2PEaF3VZnYupuYZgv51L7wgDJYq9bA3G
Td0xLeYMBcdk/a3wKTXXulqWlP43vOVdY6motcE+aPRi+8EkHXZx1QbUKTmgzWKAaKdbplbA1Sks
GdGZWmdy/AT1ug4IPAw2ZmhwAWZWqdAvmViNHxWKhbSyfbe3ZfkVAp0qsDg8bzusfV2zaKn/jQFP
Ugyc+2Tm0mv6ZKMkOLxLzSps7kj4zlrT9VktSXslC6t3TGAIVtYYvzYY/smUPkiuHLKXhWNArynR
EbMgjP/+J+62d6ZzqKBluCzCmgffP5DPoZSrbhK/d9ZjGWeDejsJ2wNRmzUMBJXDcEdbPY1VBhMT
vB7+99KpRNIhjYFYUH7NabkcgNGyUQlGw/vtWY8rBfzObO8G86HKW+3KXB8UKyI/jLIXPDNGRePg
0MppMsY8htIum/dU9uB7eXzHSRO34nACtM2Pi4zGhzGMY7adw7H0oT7ZdpgRUqjN+Tk+pNtOuJDB
Kzg8dlT/qktD+X/kTkyolKJeqjgGE0pK3DE0V4YKxRv5s06uPFqIH05ZnJW4fwvdqkb8n9eEdzHx
uywCAuK8JmP5/SKTDjcP/Mn4fvGMrhbyQb3o7k9qivFawt4wOomyxltbWLNQ6NM+0zc+n091g6Cz
o97tIwwmbhFamfB8hmerWh2pPtVJoy7BfFG42CHjpS7ZJuG95TRyjtWbI3tKDZ0TpqfdmOHvBYHR
81ekUdd7el24ueda1OQDp0lcoww0tWwHNpIwASu1owJ2TvrCuZac7PISx+kjahP8EnVlS13REQHV
XIRs3/4hTh5VHGDj/aQp+x9uxxL7c7wL1ygg4dYmZq29clHXkqDeqpG5ffbqTytFNkkpAWPRKkqf
XsEG/+JCykfB89C8n/os0fnUaR5m2WMwqu2WWL63vkVhDr5ZFXyv3Ak+qo5I4IJ9yXXYKjcwXEXC
V1Qo0gkouIh5xZXFUmJjnUC/TLIO/MOAllDJVxnPojzH5akWSsVgD2EaEBqZhgtfLiwiVwYvs4f+
y+4WTvYtzJopppEIeupEAnWLKzr0Rc5w5RsX4IpkKWPkad/8uXlHJJpRGUuHQREBDU0XJb47n8xG
32YEdqCLv0yihxfiJk9CqlBkoq8kMKyo6KG18ZbeGV2Wj+KGO4EEHxodOH7vvY54NKi1gZnKyyXf
X6sYaWfx5NbWTeCAyUgsFZ7NEUC3nxSWtYQZ/HH9ryD1HMicxwrN3YCLnOwWwlWzzQ0wzxHZATBA
AKoSLbWnnagw44icCMIhamYklP/sqBIepIf+Qv9DmElo2OO4VfeLES6uF7nHGlSr+5wEsvxMj+26
o78z0mTiZGokyjYrZGuWL1WFmBMXlCeJNyB0e1VmAuZwApLikHDnKjGb6Iyjt7t7E8iUuYzHCWYa
qbK+9qK89KUHv3x+2ABexcNPRAt93ZTlqvWxO7NHy3B/4EHKvTGz7fBTNmpDAI2USYilf1Fh7rq7
gYXLdh1S23UbNcxYHih5BeIQtw9r5yRJYhppCdwFAVxAvJ8dLnVFTQrwB/0o3dimDtEwhfN0K/Fn
XJQLglq23pqSR21Xzu6qZ8WcJCAiyt3N6C1DQLwYt3WlUXuhD6Dvt7NIrM8KloGR5iDw2IgK725c
zv7H2VPTuqVh6QdtEaViCqY4lcZNPPwRfJ1JkxLP9R2et8E56DrkL6uYVSaXOOwUAIEGje0PTwpM
1heuWzmdRMXWIVhQ6VJC81Mrfu4WR9NcoB75pvO8nfcnAJiN9F9VT3ZG59L+I3LyfSRGG06tQDKC
DATMp8EU56me4IgzfHegiJUBelfwj965htdqHqSiUIe3MG14lDM2x3vH+yPdgfzWpP5NkA/heBtq
5v1TMGvOVxvP2hoDmt5tiE9a5J4pPHSaFu3vQtTMPVSvD6mln1sBZWYiaHNQzdmyE817kYKINrFn
sgaOjevbzXoLHH/UqKbM3Sy0MWZiRnQLtf4E42Ug1PElUkauPnq4VjRPVUml4hSlC0m/1Di61hgN
eooJ68glIxHQ5fCptU/nZZaaQ/05BKlQlpZK/0dScn56LiZ9sb5Tfz3Q+gYI5i2JoBWXkQe7bTmK
yu2bpY+F/M4r2jxoezIeEk9RYlulIkNh7QQLJ18RSrYTfRsl5wHcqvlWcE20FE/raK6rddTE9BmS
IplIprFqkleCEnbtT/+jRlB8zZbsiOGoWnJhgyCjh6+/IsTxEZ4DSAuLWq0g3kNmDUCuIyDIHIL/
8HZX60jqB7ed/4Ru4L9+vNu0MAUKdz8QZOwxGlfH+zjS8+YE2GxwnP7HI+Cm78lCoDY49/1hlWlF
L/QGqFlU7n5ROebOPUCxd8ji5nPl246yinsZbtddifU3gx3JfKUEvTM5fBVaZMvXTVcsCKtb5FjN
6SgIY5LtVIytc8PGnXR9z+3Z1R0Hk7CdIEo3S2gWVC1bCBHx2xnFM4MGg6alxzmCDIXzg8Dhjfe5
mPpv9Y5vWi0U22oHlx1TDLGpx5RmQAOh/6tB4EMwzsI7sQ8R10/CHNb9GBSemmzIfSROTpzXiQ3k
x6j5ajpOwFw0b8X/AoONxJhaVWc8E/K9xz6JEJ0a1yuOWCfOheTTOpBCXuNSJfId1Dkpiujm4YD0
2lARzkGl1fa5DvbQjhl/Hmp/25eRFBMeQJfaMSEflYu9IpJgwp9RdS5WnOVnh3hE+VddsHzFhZ+R
82b+Yane03OcRwXph6OeWVP89SU0M/dCVCduuM9BAb08FGh/AgsQTC33OXbstDp1w8uLeHrQTneq
4UgnmkdO9i2yNBC034mrupoiOdFeELTalM+im+N1tyCekU9Xy/S+/Wjltmb4TlVjqAeL/Ko6EMXQ
z92KEusY6PHcVLAB26CI07jsjZYoweGoEGiaLVV1JXH07pewQs4kpdEuZqqS3kbAJuqQTMu7hplI
7sgqn86TwiUF7gojjOHB46XVxu2ScXei2Zxf/kG7aKg4+DkFPbNELlr2MzscQucG6MFQ0OGZLS8q
p8WyHsnFCCir1oHf7+EkkrqUU+a+N+ddeox6BijX2HbrAxbECI9Vzm9l3BmLsnqmBg2CeKklsfqU
h7LTvMKP4fPOo8wuqWBaTnXVYYNpFIVSfq+MmfcRA7rIQvr0EGsopFmD+k31mYyExB4V7dVOuCji
vpJhrOK+U6rvtlPEY0ZmpP8vRRw12QAdounKzoF6yoIOHRVsXx/pbGn/mMRRKyxxoETieyKcnxH5
EwWWCKPPIolLDgPcr1KWuLal0hdjOpSEgtijq3QTxqJDp0z1Yio7Ks7DXR6wc3VI3QUVi/csZCvr
UEO360PhlCnRENg+nk5/drcJgENiVPbBDa/Wy6sjDg5aqhfEK0BdSCWhtVuZejiVEdZhQKJcP50K
OFQ3Cli4zr+uYnaaE+HmHztZl8l9Ndu6dJQo4VMQZKSrLo+iTqS65TFOZe80+xqYZfACXPnx131g
8qMm3WFwMzREH1ZyHQK4lGuUkxFoSmctsfBZUlBxF0X6nsH0owejKz3ljq9SdkmU/zc1t0ndcIF3
OHisd9zwsRSYhP/kDkOMu3RCsRfBAMjiVon/SD6Nde2Tvv/XE/8/rZGAfgKCQodVPHsTe6XPWOac
sJjvyVuFSdK4pFPYx2+yjgsWbkPMkaLE49mIyUj69H1DW+UB3jdDq/UTZRGhaGlMAO3O17hyicpy
93o0z4pVWfJNnyr4K6sLZ+u4HrpV46UhWmB6UtFHyCy/NYNDCwpjDKixnllBHDvHpkMt/KxLiNVH
ZpqMwa3mebfvopow7PCkRr7CJjRmqxL2p63ZVC8HXIVWtOqIuaBXsYl8s5uJOl0hzktucQIEColN
7tF7+t3CAoFB4EmMuVsU5iCn6H0xBuA+ex9CphX9Er/8as5xykaadBRkoiLYmNLPiTbypqt+ouqc
YVtqzF6nDWDcmeaBebx693IpDKNrhLT4kqJAhDcZjSbsN5sWk02tuAT2m26s3xNAHXRc5YTxfyym
DShLeHBNOI3jEwm40SgKK9iIjR6NewRnPWCIvOMPbCNpmZWQSt+0PKMgsIE2UlBk4gnsyaL4WM/7
Mkl8Z1FuQ3jWVG7Qc02FxmrQrYunbyOzCUWk4Fs/z2v61HSUaHLEWrS5qpQKgao4guTp5G6+zs+h
VPcgAk8GEP7GIgrRwEKnwaUpG0LlETc/FwqS29MJOUrea7XQqF+tcZCDX/PH10DzfTfxyIbMtoIk
Xwo+F5Lyohtvu4J/xjVdmX5OE2uD0A9a2Te+zTqRRBLIacJTxYsgQG8jZ4KyVzsmHDGYhComAzg4
ES5tLg9KWgk+dxlN//MtC7hsCRf4tYn2VMefFuABSlkzTrSN9UwB8d0XFvBRwGA4FK2wpqDz27H5
H+VPCN8L4jh5DO77j32d88GjEq4Y3iuUFyHUdIkhJzDT51fftMs5X9043MucrbRpKJbHkI68J2dT
gUme81Ebnzhc41fcFCTIPceb93OOq+VN899VPtya5lSK7FbO8oimBG+BVw6KH7DQy6oT8O88uJMi
eA+fYEr3z+SeDg7u2VJ6n832U0lFCZPHvyJrtoOdcZlt/Fe+EZLU+KmcLABxsURO+qr3iOfptPYL
LEiQDQJ3OFCSv8w+/ZR5585g7KrPJe5OCrtVTLxXFmcsum4fieDe1NdZQMQS81PbXaXZuvGHpZdG
EG2CDVmkQLlFzcPw2znhURSIqBepbs6IYXfMDdMHyhyEAdo9VUuC0DzAI+BG8HHcCU10yo9i86lq
bA09eU53fHsga83o/X+NfK1tKVFb8J84XvlhXUPPYJQx3HTovG+FCoa9E5w4htThfCXUVY2Re+/K
4TDxScBtgJhB8WhMLsloDUVcqrAjjbjygwACfyaV93B3IeFriHfYOzaFSHmc6shjrXsHzN5PfSBo
bsOrwv4p3Z068PMnmY+Tw9HG+G19GkDXmOtZxHcJaiUR3m/ZqSAPKlALzYpHL012861Add8gAwZR
RMbNilqNIMFZLDWy+HyYw4ywfNTfy3j+MoghoCpSV84fFUuV4U76aNiNFZ51YaRviGYsAVbEwG0b
glRrjAOn1nn5Wk5jUNa1LMwB2m0raR+IZLPphjbdsK8wKOg+RvESzmfMdxlqIWeTj9mRy1ZEZfaj
//nn9SaatZfgjtLB8RoHdqtAbgPGkz0MYXYg8mvJlYm4vv9edyE9wcUOUNJ+sm6tTbsKkRRI1iO8
uV1iJpigrwYchXV4mNArTicJthEP1CKnVixXUwbgBgOxXmA171X34xl8IjZFWGRylQodNsv+wJcd
KMX74tCiK1D0ZluDg5ZO3+AnkLtvmq5BKHskU+/6j27PA/jxAqUy6+11GkkznfqA+r9XMy9GHhpc
AbQ3Cy8YRuPo3E7ve/fAGr5vZg3Ow8beoHB7X11KLMRSahyvYyZUILeIIaSBtoQYyOVpGDJ1ZIvS
t0Q3btuv3byutnBe7yJuHuUkohmSFc6x/QyCxaAqtSgoLKrLChrlR1I7gZ9c+sQuiI0qsyfyoHvG
2F/GPK9FRRmeafCxNtPr5L33QNPqhhEROZ1dhB73IMcUm93NS/hPWkTrTdXfwTR+1zkZ2IskSaa7
RQ/vZ/4HZ23azEU/r8fox46Ta/tl6ImzjWlbWDPmw7wcXG+QEzm1IRSQe55j5QhYDDijCLyzqnD6
Qa3C9a5y/BLTd/PcZc0IMFVbXne0zwDRtQXRcGkFd54f1nAciySbAFUMZp3h06FozgeJnjkx8TTM
GUjGEVqMP8W0YVNJjNrOJYtA7TSW36s+xzjajrEU9LGZt1+RZGimPdLFRwGuAM0xxuvqU+LIlpG8
1S7b0JDL4rsWPhGZbPj/12Qp6KInn3+ND2P3nXCkfEPefNwA0n8omPzKANOEjhYlnNXfCIq8y5/q
BUZrAwyp6spQIDhaIXcerAch5pb3DseHwPQioVYq7TYZ7IjS/ZeVh7uSixGnazXxbrL7SNm7XOhn
7dA7N7+kfHddSiwpIxp0I/gLw4ZxTRGxu8lhqcXI9puCFynoGrVOLgehUBZjp7GArq0XIytg6SPR
zDZyutTU2K1R8n+pDISAp5V1/pjR9IECF6bVfl9n5Qw3WlfrunZaWeA7JuhDRlcgfVFMPW01xE47
o2XRj5WVTDXpLLjRL+my7RpuFP7QcxkUaOXV7r3ha0q6VQobQmtyqw+ymNFD+2hivWgrUU31i1Ej
MAAc5iZh1nVbdVeXpcM/rg5n0KSSDwPifkI0ORPCM9KIKjWoZ1VtpbE0eYVQWcnbU2A0se/uNXBx
YLjl9kuswS4jcCYMBiaz22uJTj/2YDmtRkx+B4QOWGCrfTmIFA/xs9eYkeSFwsaKk8Mm7STKRjPk
qPGs2yeP5ypRZq6KjHnZSdwjpXDDVneO14jyLghaq6uF3cmWsrKzOy/dBXAirV7YAPWNn+IBqTxe
dlyrGWOEtkyrXBqquQ2jrsSp+cCe9Jee+eUF+maXDyiufSW8rGFlp/Ro019ZW0VpuoLLKLdjBJkZ
Ul0W5Cu5qprZHgMr53e16Yg+xkqvW9OvC6I5Ej6d98NfAUz2dnoGSCaCtJgpGGgIGEtkJa8YP/nM
eOv1ujsk0p8ZuOgzeRfMnV4dT1NkLuMNs1/xWWOOn/zFtnZduW0fP6gICH2XDdzuNHaU/ANEV+WI
FBGiefe/SLglzy7eaEKxAdIjKAp1C8IE6aPaOXa2N+roUc3ufdaFh6AgjbDDxTT/IpfY7Ar7A9n8
fJBGTi3aqx0X+7iYvCBa3wPa/FSVQFMqiJ3yiuOx94Y5alvIZiyy/nenwKbX2y7ENGAJP6jjNWY8
CPXziKxNwzwYV/mU+ZhGs75st9tqJc4OV/MpbiQglHH948leMU9VFmqKk+n13nfqO9DPmW0dO9RX
3XMUAuQRvIhxXns1c1T6xoR08n6pdpirmNvioTawnqeAEhLGPkg6i8LFpbQfid6Lanaz0gOYexEg
wHhmwOqpyUKvOAetEJZHLhbCe5zUe698vPVzVlgJmKR+lv6fEHYEXQ1paO/vzbvLIZ2dbZHWTjqr
1pnIonTd9MvvqYxa63aS8HS1/Iv7Mb/Px7nKxMd+zN+wsAuzmCw7VXGUS5yfXHTWYEqMrutb44vm
TIEbwdVbpO2NjrWtSXiaC3AYFSLPGXaivYf2uFYroLOJU2mgvQ19qL14YrE8STBLV+60KLwCJa5T
AQEn3JQnHt/kRd9FW03c4IGkVufbYaJDCyx3MvBRGf24o2JS3ZTfbgSaIcdLR0aZsK6DEvnFJzpU
wRRBtmCUXY3ewkwvR9m+5VkntWXMeBBKkTsIp66Bn3KPSCXmGhZC8i4nqeKCOtN/EJ7EN6cjXrAn
8lW5O5DxrFdF3qV9qbqUJd1ycDDGtn1qTE+b9v2ID0uUgi5d3LW94bT0l6QHHffkXJUwA69bJWH9
mHcTIqUbtuLBXhCRCWhjGi7BFxcEg2D2HmARKEvU1DCcwQTvhMYTrxF1E9P8to7yMjxAM0mSQPzk
Q57QmN5NgRxqPG6nRcPCflMSiFe3FzQMqjEKe5zyagxIW8TS+FSTBqSrESAF3hZ+8wSrJ3IZzEqs
uM6eEjDOb5g+Mkw/fDaAPmOGpSLUmmAfbCYfrd/lN26q8F2mbu9QeUOddkiC/kspHwBeYYbzgJYW
ECHLWLRq9dim7ZMDlN80RHkmktEutFfzbzAoRPp9hNnkcHAE/nAPIOjwMCwodPNtNoggtKPK3FPD
KiBb6y9xdmlmB4QoePvA59YjkxcHkjTOM8wN60iWgIJn9HkjOSKQRW4ZPw4psSORYDkZgWHrhGtq
TdpqNLU7HaesMCgwk8rhKm9SFw/7kyufnRQTvKS91TTQYKYOXlRf/izU8s5ESWhSawENgAgP7KkZ
lQQCS+LcOYXk5Os2/lG8U7NSmq1yCB/Tl+8oAIuyC/WTfLGXZ9c27sy+qjrAQvx1HF4Rh+Y+1y7F
eNBOLzsoqjRI9TBerg7cdxgBHIR6ScA+tNY+upUS/miNTOCxSd06VLmDzHe6XWmk3vYzOkMTA53t
v/08BJeMZ9MWJBSKjNMhoyOwu+13RLRqal/mRxgKMVAmuTy6BfBNRToQQoRWUMAllmw+tIzzhXHf
65bU8ZyribzvpRdXlhurPG1b5qGj4Q3NZwg74fY4EIr1bTcQn8xKwmw0cwBj0FlXqDvoL+Kf582O
0iqj2KZwMVQoycx7tQ14rL0e1nmGmkgrsNnOLq0aIe9QgiwXd8ktve3z4irDyhRNPCCDu3M1RQCv
zfHucnmXwtWCHCAcn9yR0bvEBLEapQuMvCKdDf6pn31EIV+7q6PrRTUtoR+pBlZ2zHUld8L5qaPr
bNV4qAvLeYccs6CRX4DViqwLI3/nzRkGcNE1R5zfb9utGYgq4SSJEWMrPPxr9kGwX0CIDx5It0ba
iCml/bMT64yWSbb6T2vazgGLOb0ObSHZK3tu8XGAQ2OFxsdR/F+alqZh/kRflvajfJMx76ATRuPX
JEv4Iw6mtXkHtiXWgb9BU1b1t46IVX26qaB/6fl2HOM+qesnR7EE4IAjPucFOGz8p421udWkVhv0
oeqmEfh7j1OR+5yQLUiE1pHVBFvwv88cWYujfKBFfiA9akdm3Q9KdFFKbJhxoPOjGTl2gp+pJ7KF
UKJlV7kSVSX80W8XkO+z89OzVsMV9Ntm+O2wU2WqGNiJYqxCv5x1j3m4wI+RrC3XFFqMJyzKAKxa
xYFA14A9lsluQmh8vIorvs/vajfNgrE08fAi/sx5hRUcS3DkZHs4iV7O8lx07VVQBlVFSxtO4neW
vUKnIjJdtkA2BWawL4AKh3J1z2s6T752kE3CpWaD3XkENvRV046Hus6hBGgL+6xpLL8vXYOOeC5/
5n+mln8cuKV+gh0ZJ3XkI+I1nLhBDUErI5h5XNczV7KZR2ugQf9cZPL6MQCQSFifVTWghS1zZCjN
28fbGZYk6Cb3+krjY5yQ8qKIBs2nP2Y66s414MqV9n0iDw/64ewzcyJ2vjOKpZVm+d+XaSxkr52U
NgBK5K15ZmFO3fH0usRCUeZfb9xcGn2ChkZRDzKqHUwQzMKQKq9zMwrwo0oySZICK9leRQysFLJj
j8nRLVeiB82gDaoZ4M4nAMeiHjhXppsyXjXxUQP4913kSWOYJO4Ow2CngHAI3xMmVawBAjN60LWz
KnRnzjhDrrmVRxFzm+XjAdfAfbhogNAKVBoso1iyjbeSoAmN6ugtGdQ0n3Wui02Hodel6qDGokQA
WCs7Q/FKj4nkCFTUnzrjgb6JRdai2LWe80KGlIRUbBIJSXTetreVuwNTh8qRKpeATmWfHuhPbc5P
dj+KniGdDwOwM2fJ6MFaDx+YZJw9aAfYj8X5Jxqv9+yvjkaBmvdm7ckNKKI3aq5FZJ1pfJmt0nfY
3U2obPaxm5alXxzRrW4SrbjS7CtyaQadkVGgc3I6d29rChCweVNvp3kG6t7lY+3/LmiHkEQCun7J
8h2Fl5SqZQCSUUdW8e9NFkc67NEA1GaKqghWnlNEol86wuuW0OqOmpQ9dmjf4JXK1WqOFXtrWV1O
3mxfxwG5O5je79isarGNDjei+o145ObfuxHgpZ1mJzGmLh0WMm+T/tlrKcHwMM9GqpS4vVnuERWH
Vpa9sMmJ6jxB7eU6hrRGe5ec1IyInfBKyLUhbZFdXA3jtjc4F5hIzDdtR27DfdgRhAj//0KXFbHM
70PxPfbCiVaGd0HW3CvvberZWUnenCOtdOtAW8ygepOHSBG2ndvfUBo30qT20t/Gv111tWuzz3o9
kPtc/XRmrfmDcfCb6LH8ivppUXzQ5GiF+YXTRjoefjL9dzHDlt81/mrM+2AbR39xGHn7Nva3SUeo
JMPADAQo8YhrnuGI5ynd0ycD89cz2/Eo2QRUYRkjKE3l8aiR/WNfV/dJXQ6jtgSmOHvjNDSr+UnY
0VMDCdkE6WQziyOl7jr8wBk0WIZ0IOYldtYoUkrnIN9Ma/83uzvVyOf517mNQoyIdWSrYGDzispF
UKwq1Wccl3/lpCHMMqHyFC5AP9aywc8MhqhEYFTL9OCV8thFo3/5hN/2gvPD/TORwdnjrDRQpx9q
7GuFV3TcXgyNCbysGP+X1yA/z88POmHqKqnkYpjY4FxKx8uIbLDnGAGkEx61D+altz59qIJekv9w
U5/DU5fhn0uOdumftbC6j3VLAFQpzSV622S8m+hFcGcTmLTFTZbZ1PjCEiLWF9XMghgQPrfuoagm
NU3L0AYZwfAIzGn1Y/qwFiRtnNO/m2G4ihX8vom+TYohpaQBjbq2/QITgVBj/VZ5s1IPTu6uqRmp
zmWuQMo1zKKgScFb2VA+RcdwY0fHl4QbvymPuWfpJEBTAbfM9xRP5eND+BNz7UcTR8pm9xnVcW9N
fPIn8Rxke0QSR4EYAoPIsSb4UGn7gY/34TpfMS9VbscPftP9dO4Sf0kacMjr8x/ng5aIBoEGD+Sy
wFRk5QVCPbFbV3s0DRnl+1IJN5ahlnU0Ej0iNk3iMr3avg94gs/3pEXFMhJGxq1/ISvbzLJVa4gI
P99V0A2DZ1qI5TIF93DXtyYdMpUMYQwVoGAw711yUBU8tEJErI+bG5erwTJo5ChhJ08FC8XwjUJ3
zfMDz3V7IWBIWbROMhdyTufjRsgVduqBt0h7Q+tWVCrpgnSo2RDFw6evDFm54330M7o0JDwcTqdL
UmN1KwotepqYFvjtFDhPDOdvQSrh8pXV/Sd7YU7DpAULVchjC25XXs/Yqz8VUvzststSYnHUdWwT
BO9sIIFTiN8Z/IH41K5twNtO2nXUas45tkEPGlftW4n2tQ9jk7PQjGrZHEvyZxsry8TfE9/XC7y2
TI1L11xYjZ7fry3G/Kd2f9PkWxqE1MZKIOSOTWcZJfUHurPsTgLTRR+Kvl/9iHyh7m5woJolmo7l
t61NG7sUAdo72Zbbzt5HsLcBFUNLKeWBL207YQxyi7ZdCBRKGjqM3PLXuKkwg5C7w0SzlznpWKwt
ndTujy90bDgC6xBuip3WRBHXWc4VqWMrFhuPh+jBHmznZNBmu70OS1dElsOTq2/cAthFL+9bgXBa
mIdOI8DjpkU7BTlIexvbhAQV9UgrOKuDEUFP6eRI43nxHx8Eoc82OD7auH5Gle4bd3sPktslhfgc
bnho1sajAnY37Js0a6EHQ0BNox6v69oQzn+9xg6stoui9/VV0cag+3sMMtdr1pL5Q/ejzvkw/cdp
BB6p70IvcA4PPVbvPSLyUDlN+y/ocBjTV2LBh/lDyX49UN/qKCJnzbOITiIuM3oTZEKv5eARZO64
5q8EG7mK25i5SfpFc53as12LkV5Fi4LtJ5Z17MrT8tFAiz/i8h2/9oB+oyOIHsu8CQkJrc58CNLH
sAO559gVS5cfdQGzahoG35Lc31BxwCbN9FJpfmhJ5SdhAxWAGJ9PXRXqe06quye51wV7Cd2+IwCV
ld1z7sizuzzxyAoACdXxI287pqRS29TuHWnxWQXqKC6L/ych2nN3KWmaqNpvD7SYF4aR65W/voRT
6vI1mHjmG04roy5LP/QFPEyuWfZxjCmH5f/C5gX/j7ZvzAhF2TDgXc8p75QfX90E2o2vjU6xKvmN
6drXy0bu1vWQkQZgvt9npj7sRqo5/9BXNLSbmau2Ai/49FSdSYujk6AHcgCa6BSGAV5EbwUhI9yZ
Ylu887/sgb1EHFus6s4/AWYZ9UXMoGWebEUYI6wCLBZgrGNI+DIfF7nL1/ZlrpkM2a6GFJBhkNrz
4/DBep5uQAlkTh6FGvB1Ou6VIIpDsszCDoEz152E9rWVUti6JLp+rD4rsd21voF0Dyj5pAm6+Di9
TwO8QjQXW0qXPYrBQU0Ah5pmZ1u4x64cOnk++5BmpkmCVLg8qrt3jUC2bHVlinHYLQWAmdBnopEh
N3hNvwE/AtabFc1xNVZq3/O4LcEusHox1/s1f6YVIVyMotnxT90MtGfTYU+X0i4rLB6lP/xIU+Qa
AWKk39g5wKdzLbNQBL+XeuSKJMd8xsTNeRW4hgWPW1ZDZD9FVgRvciuXRgvN/nY7Ng7J6kF+eS5V
sWIK4UhnL61VZCUYmzQuWGwB3YzGCwMAzNr3UIM0r9/X+9TCH+5+Fn0rpnAEb54tnkYviI0TXFbT
plR2vfbv9WVhDv5cnm1j0BgBi2PPCpLPPOrWUor3xSOKWbJ2uUbdG/JOd0Z5VC+VHxM7fQnGuyEU
BjkUmRnjjHUupxFhrt/ppCxef+yFySfjJRUE2S0op97vvPksuemk2E8IegGGo0sTEmH9NdReQgEI
OhvkUGoyz3M3iJAAYB8+nWfbsdHKpcgpg5zaUKhGq5yITJ9j/JgxMELmjhgD4KKU7fZ2Xdx8ZB4Y
OPAKPAx8L26TVNu55ZtoG/XLfNcdhz70CG4WqjyWLDQ35R5NgqiBLlGek4tfxi4+3QaKLDUMYqrp
6PRZg02/Kf52oeD0U484qB0pe9+AAnDjAxov/vZkwLNJ2GGZV1GX8zSwDUy0f+z6hd0M7UvswipQ
Hu4zl19lRBjVAMEuRHf2x5CW//aJo8ptQtl4VSkKsTJnknj5VwwiTSP7YxcsyXFYKiqbfy3at9R/
t7b8jNExt4dqr0vHs4zESCddV+sXfuQV4GJgYQMuyh/0PCP8B/ERKzz1w6HEghfSV+b236tV3sma
oo2A/fB6BPQJsTyXV1Ali0yZkgELPNPo5ww0cOoOEwEvqgJOUsrp4hC7eCRRI4ym5TD1T98RBwVv
pN6eUxfvYYS9WcCRIQvqc6TT0ON0Mmsk+tWVfvMSl4aa78gvI5RSVv9NasuVo/LOO+3qQSCVcb/7
jkP2icQ4AWDXxYaFehVfSh9R5mhOYYcNWWefjDWggZ6dD694Dj6IUh3teLryk4iOmR7DRuhJpM0J
kQLZoIRsWWAGhSEeN3HcqBjtTmw47dPPO9DCtpRsJ8aaSkQeWxkNGYfJRjIpAI/4pT7swHPp1nWQ
U5sqrzb+yoHjiHWcFDkKsK1t0gv0HT3yM58xl0oDcc3vVcjsBQV4NWrOohcg+qBCi31cFGHbE2yK
JWyFbO6mo5LtEGcRCEATmMUCBqX3zlMeg4RPEhFD+3rijilINiqlJHSw8CEWh2LEP8hh2DQkP+hw
ioAqUXlnNSP/yan0bFzGmeVkzffIBNmRZCVNCTUuSMk/LEdQHblXu7da0GOqtWCdXcHerGqlCAgS
skoVa3cXjEbxLjZOT1br8tbURj5Pkc8xN+Xr4cBl7pb7471n8XJwOFxRv68oWGd7jSp3irucF7po
4xeMhqvjx7Dghb2V9B03sZZSXXjzSKNzanVimhNXEWjlrW3I+7/p0ptvYG1P6Wv5B2Cg/E9D8yzp
tEi37Gnoc7eugPGjlaAt3CZTMPrhS1tcMpk6sP0YaL3jAcCDVcxCEZXIz/XlCyOwQbyHlq6zWLyu
yB39xwiiJN/y5hEl9U0UyQfdkXzEUqTfhQZikVQ8GMzcdagRQ1ugphttnyrfbfiaHmnakpA2Picg
U5KKvlempv2TmEWdkHAbLlX5zUMychya++PBcS+aUUZby+hEG0eG466PLX1NrtpdqeRYhf6drDoD
fh5JCm/c8C2EsG2lRVchZ7mEVBlSZiprxAYX5rSqt02moo9d7bW1pC+Xz+6VnEzRSeDV7bh8OlPq
nPKLdTZX0CL9obKkt5PGyPXDcqAEnDzNdo14po1fuhAN3fh452DAfILhSjWBi3Jhje3IO2hMj834
UIKM84zDmgU57Pw6MHBuIh6pmQPWD8Gj4ZFqiOVT/cXeCh3b9j7Sds5Zb/DmbcBqLTE35t+Yn446
h5+1FpDnGSdvQxUQEeBHpLmNft++D/mKHtynuaJyVPe4StK0ecXUcKV8KY4kZP+ZwAeiO717DHpV
/0cAInwCUOSMHXr7SiT2Ti/v8THbNKBHdxJu8Q1xKB/3V3rf2QuBdrg8MAmA7umTLtn4HEo/oZ6u
8hrmqNhawh+HZRxRuZ/jpUcpYUNtGX4OeFNIEl3yb2v+4xSe6BmTFrOVK96XpSaerhGaeCKCNNHI
3jeHvYiXi2IbUu0w+DepYZMreeib+S6rtczDcqIgKsdaxJ35TXkx8rDyaoxcbs5qzcW0PzIdLIa3
BBTh9pjHS1RFNIQWBt1mhHvHawB7xvNXdGZTopxJgcOP77DyW4TOdki6DniezCTcuKoEZpo1OLTm
1OpF6LnkCVI0NqG5MnW6k4HhlhjHbOIj1qZlA+rJfyZymDmboJx3hjcRk+uvRebF/VX6f93Zba/Q
Wwh5ONoSiZbwkMffKmTa248ltC5O0jEqMFGR1gnCKCXbMBjiyThLZv+S7THiAGI+/4eLLpRPxkpt
VFRQtqtrEfFvZbeEeIByjmZ/Oa+eWlwXnTj33/bnbtNFwjhngAykzdg09xARRK2DEqCt9e2uPJbT
c7/4FO3ePD7e5OyTkPydoyVwzEWuRF67MsVww0dC/UKJgDIH9Qpvv0Zh0Qv1h5Al3QjCL2VnLSyC
nSuvOjKd6TjEiSpaWe7gucFElSc1esKkGipngPuA6na+kz8XID9BaEJCj4fr5rYtGLoALqyZEwkr
VJfsBJp3aOtCl6vQtougnL9+CZPs+wvna6G1zdm5w61m748P9RDoACgSbJuvn0nUFcpu1ulQATFE
u3M1URuEc+W61PzYebvL3+F3C+ifSWyDduR36SrxZEOJcP6722Aphu8neC6f6PG4L7QXwzLEAp0v
dZC3/5xBWjWZsgnwM9j2QQojWUo3X7KipSl3H6IW58BeB5/R5qDmqHIranycslHdyGIXmUE+basL
uktSCBy1A/VgeVaLDsL5hls+iZN34g5L7tgcjP6Rxspmgm0DlBci7NT0kgT15A2fAgzQhcSUiMj5
ToArl8uznJJkNU7wK16FO3NwJVKENzOOddT44YgTJOacVAWK37WosEZfM8v/RvRaz713CsKoIH4Z
Y1W92QpqryXQsLpNH7ybdUTeng64rK44FBlBcx+j5bRxb1nFqJEazmMYJ4FI1qVZULCPazyAVozT
4BROpy1CI13zGvI10nahX129XFADWak0SbZqHu4LcNdW1W5zJZi1rE/70KUb6VQt+XMlJcIqVJS2
Qtw0LPFXW1tXe4Mk08NqyYAdC1brUoeK9Ok8184kRiln2FfpXCMReDkJc6SCYU3h3QGJDNPDc1KN
EXo4GyMAD47+s/Cf5lB7unRjL8xvgmZPhFhl+qUFcaJdyq/ufO5ddpZ4mnVGg9dz9pj5zdIVigF9
0LQEYAG/ZOCF2sjZf2g7n5ev+O4En+W9QYX3nQCZhfULlbrqfZgchxA773DYjjbYuzUM1UQSa/Gl
VoaGPy+QX5l9gdw7fW+3r63swyI4fEbCggqj2ryPnj7QaTRaQK5rlA2Jl4oGXiwvN/F43fGJWZny
T2b5grkQRHJ3JjXbUbYwZCvNDnYF51p9gXEpK5mfvOmGyXKj2MpbZoegAZ80Np4I3rIOjyQdrveF
Pt/Sz0+jTxGP6oGxyXpOPXDx/o/+6GJmccrpfJndTh0YoEJ91F2qZLOzvvhqtZX462hBWfoEREcp
Zar0wtp46jNhP1XUGXDLw7V3C7MhRBzwZcdeSHmVrblsHoOOa8Jz0mP7zJlD7W4CmSfThYmuBWXa
OSDrmmslSIyhs11RjyGfuKlhdLQ/KU8ftvBBXYdXgGZq60K/vu9/49VcZPJkelyDwLbkh852XUOk
UZrDqb2YwZsBM0d5bz2OHd1wOeYZbrrSrDzskEbYS+mEUP9G8TkTED0r900nDgPRqJ+FzpzfL+tP
bCA+C9VyC7qxAvpRhZSLfDv8La8z1rr0sToI7O4sJ1swbxgiMJDclfXiJ0y3B0Jrlq+EIc3GYHiG
3OxsuBJR6STGmaWVNPERydG1Dv3vcRMo74Uc9wFdHQOSB8bd8fMD32YiQPAeD168NKSP/VQz3g7x
BVXNIc/GTXtqKIQrjNlxzFHhl1zSkDlpY54vWe4N/8+40X3uNxwUalM2NIR54A9V++IOA2UyUwMo
x9nGOKX29pknWWeRFjSke3VG3zuLbsW4LzGasc0J2lSoCuHb552ky67cZN8LZdiaa+751fyypN7/
hPsZcvQMGYrvLRIrBehlIreWh7tmv/Ayscw9w1eKP+LSn6+iKFg7HgI3Xh49GFmg9/FEL/f5MjCz
ychgjSFEDoWSoVRE0rlAZfjzgh3gfbvjkZwhNBhe1A0PDOnXy++ZfbEni11PfA19IyXkKKQQQoeH
xBPkF4D2+yDDnx0mIL4jidG9lSG0OwBWQm8YxhJ5JO7Tz0KokDm33kC8EnLSHw9z4WH283sG8SPV
NPECb5lhQRVZ7u6v+CoQYn8W9rV/9U3nyQjEsld7lCs6C128PeXqcXO1Sdr82IAmrqZ90NfcvulD
C6N6jL7Xuxaz1Lir3rxnhxo7W5BEtMUds/r8ipa5zWUmhN46Uzenn4qlHwUBNith/ghLTaQiqsrp
hJA3nLEbLZXE80n5z/U7HU0o0oezvN1CsJF3qAIiyBeBPjIYNmum9KlquyNyjGXIzT72eMl7CAsu
TJECLqDp8k1i3b6AP8Bbo+vO4xp8BCDK9kCafWfUFKiMYDH67WK8kS/bjdaGeFNCOKRhlwnzJaP/
IivglrM5YvlFzOI2IgHChD67WJ7szth5j5TfGdIfVHZMRKIQoBImDRk9ioJXchWm3CgIMk71Julh
5VFoURwdyvw8kthPU6shoK9I1mM3wST3yqqS0cRuIyCKKsJOq/94fdDuDLUZfFEU6rViXZMIhsl2
4cl/MYYblqyRT/Jy4NflIT6B9pLSvV2eiW8LdNGJDvFwcUcf06w4fdGoxPJCVp/Y0t/yW+dZMNG4
hxEA3Jr9yBixcUgGB6vMhe73T+d5+TUmVXs/qRkAXEwy3FcoxZXbrsZbZS8WIHU6Uv+FSuK8Qy3Z
ECxhgcQW5nYumNEeaJ/Ddj1L6rCCUg6NysGrN8BYN0eFK3PNvAAGHNgUT9LXsaMWv1DgmK0Aetem
ji5zP0vtYWzkXRC8wiK7x5wRxSrhgphZfJF9JhTVsRg+Jzftlm9I6A39jXbUi9vBVMHOG8rH1Dcp
TFL1QpHWQGQxSsFezRHmMHp+SxSv1DvQbhS7cI20Bd8wz1ClEs036pXXGAV4+zZKat69+kseN85k
KP9yGTj49fxpPxO69K8BwXSJeMqHLXJFiHsh6vPtIlK+KageIT2Qri+YQbBGh6wz369bzMamAa5L
JV7UGhDw1lsE8awF2PHustn2IuX0hOV96XKXaXCaD2BnQ/kASWpa88H75cpOO1x46IaXan6oGgBu
zPeam6x22stThCpuNpcP7z54Rb86w5UHM+ePt/gh5w1xU2LmJn09wG/7YVQTnc7zyU5IS/sD7UIr
/MVwvqeNsVKK32Ticvq/2P5ofPAZpKsSN3PxfBgTrakbNddSJYg763vdVVWGlF8jpE75wRcDTOSw
ARRyt9natFdrpyMEE7IbfmSYYI+OnlEWyf+ZMPf1IkUiKK7zZCOhPZAss/zYD2owMft9Oe/nLcYI
RSnEoqlfFP4dM2BX3Oe4lN0iSyotcljMPUjXASuXCb2B/Y5p3hhQg6ScWdQPYzEyibcLU37b//DZ
eqZNLYt5j9RDweaB1m7flJn64q4/SOK2xO52FPEDle/hzdD5zxrtaoXUg9sD/pNTaUrMO9+Bi658
T5yB61RHrqdu6mH8MklMlJnVBlYUY6No1fHmMNoqOvTEyZmRNmPQH5Ruz8zF/MOrNsdn7QBiplAL
wFLW/RPpmaJ0nZ9vlcXNRXHO3kgXbqdTVWGI69fcgjKiFJ+fkeZsQqul2B9JpQO1kdM9xEgHXf9x
cPGLR7SF6waxek27D5i3MC7gV9CMwSWd4Akv/H6jzmMSqrbQKb+Nst05KKhoSrAX8/9byAtdIZr3
5C2cRtI8wtjPricrq8+Kwke499yhhDU6E2qNRHrhEYqKqFLwiMJHD0bqZdUJ90Cid8QPY/MYO6Q7
USG4TSFHDvN1pGkQvusphhodznycjmJSN7KBstZpcERUH6zqYXNNNj6JNoecTEpPBf8G5HLiTSdA
n4Azr2ImNazzpII4ANZPaMPOmp6R9X6NapdMjrA+ao8cucIMgoaEVKtWnv0d+Bx0wKaU/jMNRLKa
IaOT4wFT1KnYw0ykxujjAIU8p6lXj3TTNfbW9/T1zS5rNXjl2D/pRYLx5KCbyRE4xuPqrmFgVZt7
bfeMgP8AElunb7iFKos2u+FM4ikyTCuhB7wwRHuRoObWdhw7KsSMmjQU+6HI1vEzrMvorzG/y3nZ
iqFAHmYcYr/9ANBNRFF2d/e5CBqPwucDx0/mk8DAgG35TOxFY56xMxfBc24pdfErba2fycFC/j+F
g+3HVsypQaJB+Sme8ZnBUsTw1ckxQijg22ENcHga6nOHTv1QK6R2LYNYuJMbC08bW3iV6+fvM+a1
U2eaZhf7XGIctJCFAUNeymlqsGn2FEAJUIv8B/zcdvYYS2aiCAfX7l5KpqwL6B4O2Vzi5m14Ws6i
GbdZFtFJ5zuVO42EJbuZFeWecQx5ehssCIkkFBzChi8lm6YnSN6r1u8jMuCD+HFr6QmvOSryfKbn
YkGIk9bkaKBnwA2mHEz2WK3KHcaR1CiDukduhMdAZZdmmko95crLhuaeNgnuvAjLQ4EeuWJc7qdZ
YUpuaYJMeANTqhwMUocse8yDntukNQqS/JOu7lFWzN4QtHkYsyUj8rJeXg7rlk1ez5bXiuBBBoQC
8Tzpy+TRCUTSBj8yDyp/IzACL5yxjVB9KBJn1PdkGfHxBSqCwgKKbwM/ol+GoKYJxJ1U/IMMqXfp
RaPhGgG/PpdRr3+Y5jqO4gxzvzibvMW2sziCGlz7ZzieEHPCqQVahjG/XaH7Bmqz/RinOCwRSs+q
bZUMCfco/YHJhsz0PVQd3TXOM2/q/QwD/tP8FDwSnnql9pjRCOt09RbVgmNYYQSwLFEyLqfkYrvR
bfZMGc9Ml29E/ymf6NlJjB6X3v6H8inDMEZYu40KYGiAWRKZUl/1fkMJERilqZNomc/gbmo2njuk
YGHiAOnz2yFXFJVJ381/+pO1AxY3h+zn4Z5dudAL2s90E83V0ivcBpPK8DxvdPFof6A43HhMFe6M
7R6TjFHZpibDLT7bBaz0tk7TL/VzrI23TV/pS7ZbnylgkPVvXzSqzi9JRa/4LxDtxUEM3GFf+I/+
OWrVOYltmodgU2fMN9ZkTlpGGm5JR/aftfkNqsoYRWagkpI5PxkwBPLuJyVW6UYhy5D8Yd5iKyoW
nNzVVqAcWGGUuRHiMsdzPsf+Zis7pU6qkIwvoFmueVh3VV/WFbU1oJNRYSuCH80WmiqeUernkHww
kMN1IpMBuq64D5O6X3p8IW4WWV+xxSA40q/mvpMl1oNHEtATGHIqKmyeq345kgSdQjvQDlZFK6s2
9gcg9JccF6J4ERTIUZtVmEwV9d+nt7k91wpnMULiGEa2nVQ9IKAsyzWPqQBz8Xr4mlM8C9bV34mu
D8bunFfr0PlPXIQFZJFko53+wypRuSjQoBKfw13uMf/3l4nJ1h9sS3XTBkqjlHPFW6fCqp+kyVkY
QZ4B/jAGURfZU4kA3KdADWIrAotbpWecaokgHUW0076IXZScjRZVqqs4oRiZSp8YqvkMUGapiEEB
AW9TkKunXuQqeWUKR+fBhvX0wpbJG4FcRBULFQ6yOcYW4RguaRMEhM/+9WkpzBFwahb8aBGk6nru
/SxSltaqxUQMIIFZ85Xr55gPK4GhJt9vGGZVXtOoLcI+cRXeIJm+ZSVQgQoymYMkqNhJWWJk5k8p
/IYJ9JuDnkXvCBXKl6wzjktMypwT2DZqUuUWz2Ewap0uuFQs74BfvYinS9YLyB1+ijx2jHZsX+cB
1MWgZs+5gHyugmtRDe/tg1GCFaWFco4ForCxO1GuqIxB0OtrCCt8rAeMOGyGAdqmTrbSqdC11eqo
usSopXC+TB9tmph20TrDSFpaU534NJQKXLc/zKSwPD2RVAkFMAeV4+k6mYgylpts4KyoydC70Hah
NA4l66/lzTJXzSnB/neH6AbzQVMLjIfHhJkcj6p0vZggUt5b37752zvCfZC4rjo4hv8zkuwODd2M
axe5y2SXeIgQ4cCBer9EsELKfv6ZYUXGzK6+p4WYryExyCaf99rXuWyzVNnXE5DEqJaS6VCxURt+
whVugUKR1uKgRZDRh6A1aN55py5ON27qdC4Re01YaoJu+y8Lc+oeRrSYW5QUo/h8pMtB2u+fgS/e
M8p1QvmTSol+Ye0bIqJSm76YBctrz2tfrFZxkeJODPCqARBEApxe1J302O1KQGfMM8mTzcIrl5WO
0ToOZyxXsW9mkWPD0c4aSrStMPZw4YWipIrzmKgw2TPXp3DVBMSkG2K0QTqY+K3xjHPxG2fJDDZN
0pkNiAv9aYdx+89KeUR/U9Dg88Vco/LBV2Ixt3y6r1m8AsZgGjbql86V7I/oxtWIT8sQesiiwj0y
+ITxDd7D9KCQDuFbCvOk41RfrHWWizIt0u33Oy7WNqoC4Posy1Wx28rrTKwE3DzUMev8d84Y6UGk
4UGlc1SdB7hv7YXHLlPak7PYivzJKSMQ5PkqvVINitSnIF3FwygWUG5O/fH3KBOpNEj1mg/c+IMw
5R7+asYtc8kMCG6W7roumF+4ejWCf6UtZl0Q9P34EmclNTn1cuk95Zr8OTkF2uq382wGnMSqU2Ir
rPRbUMGS6hcY344U/ut30InkL0gkwH+YJDqYN2HaBYL3XVxa+D5RHeJ2XDaaYnXRWqHcjVN0QSMJ
1hG3VuToQa1uKED/BJC4vvO5N3FR212uH+DhNgaup8gFZNRNggBikH5UWKn/gwyxf6y2ts3GEv09
lssyv3kvAQwcn5bB9kcS8XVcTP+QVZssOIW7/BLvSD0vLDYZ8SeIWLL/AWFY0kgeQJbRSMEKaOiV
5qVIJwa0YrOX1sxPvWH35T2Kslfa6b5dgBQtJ3L3kZFitdpWNG3Vth7LgOyTrE28D9hXd/vqDTd0
f+TCCafjFRvUL4n+VndbHiiRYfWAA7aaLnYF9S1qsgwdvD+tumFGi/To7G7SjNvkbCVdaJO7nhaE
BU8C48iE3dPBHdgP/IbHnZrgLi+ye6gHg1YV9BbmTnja42m3xs2cXqpsKLBBhOCS9Om5SpR/pzr/
ziHDoChxO5kYW0wBJyhUXl3qSb69SJPvkwM5r7BTc8YMrQjmnbQTcZ5WKqrYOxyhE5PemLyY8ewn
rPSkL5uluofoiNNZh8hO01WlW38ZIkSDeleCAjVhucf9nYP9sWdgXLU48q/A703V9Xx9MVz2Rz6I
kaWaZZ7ui30ZjP04EeRJ8C2uunGfA5t0kHpihzPxj4HfIbiaYj+rgaj0ZuHN/c4ENtYrTVQ8IRfd
qRUnwcEyYs13eh85DoRYHOYVKlO0c+CYpEiqU6InsmaHVod6e7nL+cKBMX0CCuNlh6f/wNQ4Wv8N
j8XmihXngJ2xct9Htu4E4dCcRbBzU9AAoUj6x98lrmHIPUrmxAinjSxs+VHGG6uikils4XTpoNEa
ruys8jg+cawfShY7wZ9divzgaIvNqCHM28+5oE0sec5YPVGBnMSn5OyJrDRapdWeIIQMcYE0Ekr3
q9dTRyh/MywrIwf1RH8u22CN9bb2+gbZr7/Zf/TVMJBYAieCpuLetXyRX8cRInX50kHVDWJDRa9O
aj+oet9U3rBtoDqoBWukCKVV70wqJA5Iyb8rv4SbPQXy6FfYDgtsuRr+SiiR5rWF8t29re1ZXNgQ
nzQrrBoM8MMSGnCrV/ZtpTI3Umm+P8I3ofA9o+wZrgpbKO8TCxbj/iuBVxJ0IM9YyHalGloyI3dr
6juaJ9b/HdOAeimvHyZIUxRcFXcNUNexZimpjdq0p1HmoKqRbnyZUW7PaClL/ARn1w/jy+fHXpgc
OOlbSDc8h8G9pv/tLu9Ov8MlD2vc1kg9f0YiIaY7U0a5NPPBKqxVzVSnxjxSkzu+J6H2JnuCf/Re
0w3fScRdOF/ioSlYYvdMbFhhZtcYDejwR5Ah8t1oS4PDoat6KB5vRqHNjCzvGsxgdk2KeN/M1dwS
Ql5TdhwkkUatAXRR2BtbmS6hJGeSQHvuMjpQqF8P4ZVpubgDV1kiV32V7n/tX69uaaQkbcwMRvuK
BsPftCivDYpIrSh0ffrF9UatvjDTfzq4anN+/oHmhLE29I+IxqC5pN0de5QTeHJ106hQSTTnEHlO
uJ1Ac5t0RR4bx05dbM8LiOrio5XEQxxvSsFGcPqdyAajC0QYcddtQmRoFgHTn6vkrhLcbgWREhuI
ui7pbyLTYBOrlo+5mgPW4I8NS7+YGUbIFd0NhsVu8ItGLp9gOqaf0bo4wi6JA7oyYbkhCj0YptzG
pQSkLEj2TGCTWire8d3qPd5Nqwvg1XPQqK5cHNqTsy2dujJlq7yQZzf4usZVWZ9mVp9OGQj80dIk
8KPmx7/HONmXE589f0LkaDS5G4loGNht12GH63y+lD7hhA+DR0/QPaQKU9ynOLlmednP9Lfw6HkT
K50/ZUeDqZ13A3nkJ2mBxN7S+4hc5Zhczn+1d5w0IpqVK/k3DsYQ82HEiBC7VaB7j1eIWL5uR3F3
WqSisGcnRVXRUNSt6WITge9LOrLyD80iyXQsL3eqmWPAGTh9DJF9ZdGuLk+dUrOQxJfDqPv2SQSp
BKlydXm6xgsRnoFRaeI4lyBBbDZ/nGf5RPr936ADJSvZU3qDc40Mzyc45P3ZD8JpTOa4qjNk+4JD
l0TVsADyq/Ju20pQcfn5bcaciBkciOXAK0R3HgDc8Sh6TQaWVUwUMeF8z1cT+wzHjX9PonN0W2Zg
gJ05qa7PobIeljMvh9Neiug+iAPR/iY1iHyHW7LVubV1cEKyZA7+sOQUfPiYKopsi9KV4gLbsckY
hSsGcKtLpaVledllx4pdu8Fe1s3KxpcPxInq3dnYnIUnZfUP/3pywFun/UInHra6Mhd2B6fw3BIr
7hfIjIYQfJANn4+gWACW+yxUi6fONiTMBLPizqkyNR0gl0i5c0UvVC2pt0oZSFDUW+Z+OlFGMWvZ
ZJE0VbWeKmXKQMZYZpVRHU87tazTA5EbspZe9PGqwwouZznL2e7iI2u20q6oRKrDiAfe9PIX35Br
zFfF2knHw+wqQtK4taEbH63z5LPJVLDjk/p/7mwDRfm1bGOAW/6aN4DwH1ELKtpHBkBCkaC6zrkU
1WJo3+31hdE+8YI0On2NjtqDiaPMqyJwoHwCyhHYmcYmjXyp5VLZvQ2VR1SV28+jG28muKFNjkp6
T/T72jKBXwtBKIwLk7FugIgVmDNyrGuuDq5/X04JMjOMwPzEA5ZfHl0l0gCHToqw6wg5TizVA4oX
ed22yV4ukZQh7t8qGQ1OGEw4uYPEze3LUGg/EMT3FrTjJDYJo8AxsOe3pRwMARvknGwDb1Hxqprk
ipseiCWnH6Q5/wUWaRQzFM/0c8UivjIqbKsUq1wJwL8BKFfyUqO8aGZJ/dnFGzDqq/KJ4hhIrl+h
zZzD8Pjl1nB+jY4CDwGW0zpwP9bJviK+oICYCE8tkF4r4YlHdqfU1njfdNR+Y8q4XcBl+ZXRLHWl
BorDYYbnwd+NWKH+SlmJRNLcX+3lCMnJS/ow5ElyCo3DAmlwvi3jmI2FDbTU4Hu50CsVOGbnMzBC
DXBQzfl2DV1nwePgO1T7xZ69eb/TG2DdPciD+Bo0G/xGrdfz2AFhijAFqZNhGip07KOqmlUsJmGX
EPKyX6llFuiejauxnnfVuLgPoR6xCIApxtA/Icy1bEdQo132JfxiU0gBvGYOp8Mxp9ckRE3dzuyg
TR+otO2S1J3g/3NefMFnYkUgzGNeQIzVYmor8TlBwDkzBcTU7vH4qWaL3imOQ8vGhnD/1r+AZZjm
GT23vkSEU7SkJJ4H9qI3HrAJOk4yFgA2I09xdscmHM0nSnZaOcqL/m91ooQ4zLCSxtEve9sNqltZ
4V4F1IiSTc/9n7aIj4I9BTQOO6Zc+Id1fAmR2tjQ6VIbS4jtljPoBlHBish1uqdcLQAwmmhWuTU+
FfOOXWTHutua3043yCGM7lb6qSrgLlTt1hKRbLObJLmCXae/EJAwh5aoMpyfBfv0j20CJ25J1mBq
rSeXqdO9YH3ZXvQ6JQMm6A0kwnEJQO+bZ+ErNvlEm1eTTW2Lb7TkbFvqFn/qwcuO9MQiyCQ6YwgL
YGfmhL2IFL2QSeHz3MjW3E5+GfuLSjP7BtKe41AoRH6JuyAvGcNiLVWqZjC3iOhteEW4qekKiWDu
w9e0YfvhE0gXl2qfjichf34cr7Mj6VyG9f2t2YKA/aKCPNao65yEeciYzloSjqdiUy5cd445IPTm
cymP/3IIaRB/8OiaNyXw13BfE/SyVEn0IjuvMMS8OezdumJK0kpWqFLGZWpVLMGSONExOCjqXf1R
rgKmfg+tqQ4cdnpld7Xis8FPRk7UpLMmFaZuMuLLLicYRG9xrrJCMIO7FadArHKEmzThlOoNHCSm
2c9lNawcHEEI7Wg7KhFC4uSYi0scEQkrR5jRaVvPdtH4rqqnByyamTLI9jI9CSZEG3Kyomau+Dnn
yccuh4UezdRLo4B8UXow3LkGjbpaHyyxkD5HwBmQWie7MSpWBQ3O/EPv0OxHjTaoJq2HWe6yxHGT
hp0DGzMYuOTuiA41fjLcWsq75HUlYxSaSzIOwoOZcSJtMISJZNHvmKGadyOl5/zDQ3u7qwZ8Fd1O
z0ZvU/7NCxfvJ6GqkBomhCXkkwM3KPyCMG9aHWldi9G02YcIsiiZIPlpSNIZ12b7/0ptBbrw/gew
hl4pfWiN/arJakD/M51ouo9NjsqFl1iTjyMo4z9o3g77eiaulhdSugNQsQWG0ORb9+qudBuRRxOt
pdsLt2ZQZdG2CjXf1K0FiI+5NMZneL6mJ4hqQ8/86zangwDM06qiBepoVqLei90DduQdwHGXK5Oj
NlPvIqvuJ5yW0bbM2MURc3g7xwF9Z33fslMUDoBqBwETBMJPvnNYVLsSAVsoXE1WKXKZwwz+qDPV
Fd1chC1iSEg75tCeMmXDOf8QWfoXCJg+zL3tvksEFzcdVDmwIRzidNPOxflCZqJFHMmYEaVX/qWb
AL8weJrc53Ve6qmHMsiFuz9JXNRJCbnbFWaxDDaZDFh2a7yUIdVNgrKPB6ZV7w4IUzxAgdb/8AHE
9NjnbEO4GVQd8B5KJ7wdZ8Je5QfS/XsOw0bi+Azaob5E1chxlPUX/v3I9ywEnv0C2496dJudzqmR
IBbvuuYVix8Bh+irR9r/U5D4xNvd8PSbsc9++JxVZ0a2raCEVUFSrHrjnPEEezPOoD4hlq7tC09h
bL6ZoPGz5x3blJ2+WjO2InHDwRh1gPQN7eREN4y5BckEmQL+mkmSIQdj2H9gZ7+r8YtyOZAu8hCz
PTOTzQO3HHSAAyi1Ss+BS7pjw0R3W/Y5/C9qxNdnouHo6s2jKjLfKSzyzQaZcPSUxJ8WxLCNcrh0
rR9pvgHCkrjQ29Ut8vMxKUHEKoHQ63ma/0xrHyLOpZUUtKIsAkhYLhhPAykD1A33yOhPLjCSNHRt
678vIYwAzTTLTlTlWjfPFun/OHaQikp5HSVTmoiS9z3UvoVTbF1RBPsFENOaBu1y751oPAEIdT2c
sEp9nRB9uI38pEMCPWFTPkwHauDO0a2HggTMi4XePkV+Qedienbbg+I/oukhdssdw1tODnT+ZxkC
LjdxHrsB2fgSXDnG+BasfcCG9fmePuqSE5MUjNhJnGxC82FuTIiRO2MamCg0FEQuzfyYpmVpUOO5
aEoAIlEcaIm48Bz/iGZBZtCaNTWsRdWbf4t013uERh++DWRHUKcT52RqEt7eEZg6AxwgfUi1f7RD
Rj3ZG2MHI0ZG88wXlSoXyektKqTJy0Sun1RlQna2tHwx3FCj2iowQzQHJfxOUSJB4MoTyNo7SfnS
pFpr43nAfK5b4/LOhuWGof2Yz+13498JDGanRJajuxdhKLeklTQd+9722jv8Ryyl8MEv9SIiBh/K
qq5uFiBZTQCX7X9+L7ROBlNeYLmf2zr3u01dDmIq5bSl8G1Cy922Fm7m4S0CEsoy/O/4+ANsBrTc
zec1urIz6h90zqIW5Kusouy+xgfnry9STG6bqc8/MkNnZNpFbL9/XMkmbamqe4p/zMY1iifcB4Gj
cb2FO6XUVtXVOPUtk++AY9QaxKwj2uiEKO48+q6TPPPpfuofQztH/NHUoe6GGU64JjX51Dc5d5tR
G1gPObY8w9cCB8e4u4/6/Q0ASCz3uuth3L5esrOjAdQDTZ9PmTX5fIkgxPjWyJp84+f4v8FKjEke
o1HikmDhPPke1RS83skiLT4kyvxMn7v9hqb3cKozAWdpb9AOjrJD8GzGnvGIdPMgTrE+HJxB7iG/
Wldk+sF9g8tBgZfr+kk+Xp8zySgPxDmqJ0WeBwelSxFjr8OQiOq+dm77n1JbI2kV+Un/D4FkTgct
9QKPQs/ooIzAFDk7nErsvKP7VzDV0ND1c22ULezPIlMgoHLq8pGWR++vzIuvacxkn6faUEQd7Wn+
LjcgmYnpwJBZxwE41tnVJqbueVwMhVDqHx7X8nL3XQ5LmAOXdFoHz73dE2XU+ytqXk8vtVcxqFts
i2YsZDp6kbe75TGWCzPESv5+UsWcK+QiQ0Ik6E3M56IJ2kM6cit9oAPZ/nud+e3IoCXwBnAehHA2
y/sIA34AriZhLB4xuf7qTTK3DLbx6N8zPLNhay0KLvw+ttLlKxm4CH1trvK5AtU5kfzNggtqC3A4
r6Y1sfmYeDN+QlzqiHxPJSbilcGUILAiQNPLZYAPHYYJwecuowtqMCJAfueahtCfYnU5FbIzJfDQ
vekDpuM9uKA+dbnjDF/aJnysjgDSktWZuPXyuOu6vJqwjHA5HZx4svJy2lCl4kOlQ1/RK/7YlECI
FJR9j2FsUOsESP8eP77Cq0mfWrWOVPPBol6jwwKzmKwXHwdIUKMTW82/Um0zRFnjAO8o9GVHJVce
TzQ/dtpz4oVJPtfWx55eTNkqqLd3eg6uL/5VT8lEvJLPD2tMlnVFEc4rYM9d0Fhko1mU0Jd9RtSE
kTDCSTyXOJkjgChnA35a+frpiPKJX4DK/qHRE9uYXgSfEpQ9GL6+2XXiHjvGT8qOepOjuzkyPW7Z
IylyU6x9c7n8wdUAjK35e5aKOwVTi19SLy3MRhdkj7SYEmsuJA2NWWc9S6pmj8YRsFb/wtsePh7p
q6ts9RThQknmEs+7fU+VyaB33a7zZNDywbr7sEHO2f2TDDkg3VjSFCYhs1xtQMRxjFO0cy3MaNyE
rUU5TOAPGZoj9uFSFNDUlg48nGTFgNOMhC1nllTZpWiqLddJNeh3K5k//p1KPjSub2BgOleI2o1N
syUeaYdXhkla1GiIr//CuHwrfCs4MosBdlEdSDH0PiYZxV57GXm292gSThUMYJVx6WinbJgHUJMG
Y7WXcs9nVbudI98o/ZB6GXemSHVbYtnZzIWiEgCy0v9HY39QW1vN1Ad5iN9fObUkiW4QVFOsMFY2
LW+LLFk2UhkW75346+EUW6U3EjcYV/TBvtIMKe2mVosiXrByGRmZvc+J6xgTwymxzom3NDiRrXcF
YR/r4tkkiPQDPTtlAA+cu9IS18xvac/0+T9HzNz3zXutuMMLCK1gVfmvdt0GiTny+uR0YDaI5Z0p
1D0VTBsaw/lqTM6taffJX5qh/zcnYWXQerDPf1wKBl9fFLAXed6DwUCBM8FKoBN2Tbu6AyTiYTaC
Fhn+0XoEMs1LyI7+tAJ807Mq2H3MCkxgYE1EdIq2Bup8JtIvvvk53VNhbHaDSd1ikHDWmGcnH5m+
46Y6eEoByDB670lRN7XRgbC+3pJfRb/j6t0KGqjzrx83LjDAFoceUOqNlVQLpY0+E6dd3oygbqMr
v1K8n0o44Vw5JvzBwE6DMEpAl3GNWOUSQTVW+VVo18bGi4pudrJHPDjJU7DVXyQeCykTypsYk+4E
9tFOjiXGAYuDMg9Q3zOPp4NTmyzmwADE1iHAH9gsIz/NH47C0htXHvB30VWcAxHGvbdCFvrYJewZ
YK6GqOVt94IfNG9nX7yt1hOAAajMiw1Abc4PMhRUZSA0KXJ007jTFGvzHKmG5/Gj9GALv+0r7CGA
Pj4bZbb8arVnuHkmb3H1ILomnvVTBYR5SDP0t0stQSwMDVGmmS2WX6oITimAB7ACiShGsdlwIVVS
s5+ZV6ow0MyVMHIa3gUHTfKm01aGKxE4EUSJQpmeOGhptL8d4Xtj1pS9+G+cAatkOHVvemRLHTeu
9e+lYrREsub8nQvJA/W3oEQQCc7fiZ/PA+Gf2EI7LgRc0wS9Vqt7sGJIi6BNdzPuIucN1MVXZGge
P9HMzIwncY1IzfWRDmKTHfKWD1kbl4vC7qJjqA8MCfs6HeyML+t9J4nSSAeRmoKoHvGhtp4uAsbt
vi8KZh4kgyTDZBUYIkxjqh7ZuEbQ5GrDqS3G8XY4UcX7PG0eY8Y+X+NTiJNAUTeeEY08cfBMSe8j
Mq7pXj7Dd79btvmEi3IKeGNvcJhTU3D1byPfHs+7+vjUcpXfsqhqoufaAGhvHiUg38DSMIw4hYd+
pWZV7QQ00HR4I9UWL7sQOzEgRxtraSYyH+i6HTT211uFRAwgXU5Fgpxl3vtQ81i4NS2E/JZYh2C+
horfwViAnQdffqLEgAMABcom6WAS3nMzahW0JMjpxPojZJ1q3B7/uvqCxzo0sZBeAMjKqov3YeuE
5CAQ2LggYaF4tMxDMbphoBzoh4Kj5mk5BogMen/i8djic8shsSkNwr1BGUzvedfTrqNNnYhet2UF
+rle7j+xX5UbETSU+vvp8HnUIvJ55DKo7ztrfFR4aYbiNAYbiW1b6Kd03/l9eO8/sa8qrhWFvzQp
5N2xVr+Pq4ms5YKD31WJAlSblGAhQZwuBPR9nAOdM8shXSM0EkcrGycIjh4yb2/9+EbXxXmZAwzW
z2RmegN5LWdGKZdZlxYm2kUi2+RhbE0vMWDBAaTZmavm42a+JyKPwiwg9RbEc/Bsfq5HCdJFgXVN
gLN2udHBMShLaKJBARb68VqSwVCqibU48mi5Nvl0/1q4A18F3BMdJc3hGq+NczJw9h8Ee1wcngDf
zvwEyNcg30s8BIJH1SjwJvDf7r8RHxb+tQcpiB7/sXG9SfwslPuf8kj+XnBCHyPA1NVcZImq1mC8
bosMtibzNkkziOMsp66hLj5Z0onFMK7cKIRWmC4M+nPurj1rDoTRCiz09eHOJF8DM8LRLIm/O+l5
gTeRi7aZmvaP30kj9ROsWzDsdLlonowywBY4l9mzdpmZFxnKtZYKexrBzGbFdnV8PViVsi3D/Yfw
wLUSRwFtPazarpq8kI7h1E7aGznfg8o3Rpk/8vIHeWlTHHYigrYdsz8MVCAfM/ntmFLvFmB2yG/E
Yd57Is8wQ1UiKyYFqPDmzHGqa06j8+/YdsvJ6rlvx5/SdK9Wypn658vhZQj56zy9Dp5WyuyGgUST
vfIdRYAZ2xr/qZjs3OwZsPEd/vNnx2tCiaI5oeq78kuX6T+TzG1gBlI/8jCJZbTDqiGWtoQjV5pv
zmTbwx5y5QTulWHHxLO7W6Kua9Z+NZCZv3Bvx2Nu2Tp18f/CeH3fG+2YCyPSQfwFu6I2WPlwd+Ca
SYIuj83REuZrbyChHd7hCmrUEqR5N+SmtSlsoybONuYI5VPOr8D9jtFSz02HqXst7fzK3zL01W/e
beskv81H2tpalzyUkQqLQHfKhHOcB3GcvQvE1EB3edrfue2WJVAawqfjDWUYw6tJ+FfGt9QHAc90
VjoyroCLp/RMD9LJ0qmjt47SpjuqGVOkpMqcDt9zMslp6SyAKc8cMxrH8P07AQtAn1Jt/VRHDiT5
K9ESeF6Wo4rl43kr9lr0ivKjYzI6cVhO2Sl9XNc4oP8CbwNeA5sN+TNSgrTWOKoZVLdUqdVWe9YQ
hkaYSJ+ukG2AZTZY03yJepe2XE/MzcMjzwaDuXXTq+d8WKMb2WZyNSt97nUgtBOh+FzU4LAnFs7T
3AkJ0/6lR9DYO0kyKJA51KKnsMeOf0xSRNzGyP7PiFk04TcwTdQyonde5bTTdDIU9dpvMmTQ6YAO
S/4+uZAp8/GNOj2gWaTM34JxNBTKEDONnePs4WLvMToELRA5WKtIyRIQ8iYRLPjAaKTFdq8zDhgR
8pdp1g+9UMxzWBiAVT3DMDqDduW+Pk93sTW1DD+vQINSseTAlBmtnC0LtB5QayaYAuRvaZ84dqBv
YS25Z3185HFI4Z4noNuxtqIdkLlSzbvmU4tpoYX0LjTrd7Kt0+ZzauyA2CHhztnklrl8LOs0ukPj
pGLUJ7GHQjlLn3Z/YuqGXKhiiw4Frff4tk/aFDSbcGhBnRzT6kTz1EU2CC1N2wK9kEkpR1IwAfiM
XnwtghlJC9K4I3tVVPe2l4ACZ5R8K9ATb0eD2Fo/pO1s5WuaSIY3xN3Lt8s7uyLMBvbACu6bDvcg
aVhfo7YAZMwE/JuKyez4uwnAF+GXCi6TsfqkN+VvTH7+dut8r0qPxVYzqMSY1dDKLHSoGtSa58Pk
FlcvfeG5il0+WkRuwBnXbRRcsLvrbww4trmWPzDSoG3dNDYyMPVn3EfjX+9gZNSPJvqXjwNrm3sO
Ggv/Vj0IGEu67YF/gYk1UoGqVxRAM7TMUmytD9hojPa6eF5Hwjv1mWLf4KxbIQTxwbSzIxryHao/
qER0n92PoIfYBQ/C/jjXioLb/30YH0pQm3ol/EcrolJF7v18PnG3c4qQtoP/OWzNpYF3zszstagT
lKmaPWtqUR09R41zZy+8gqawH4SEl7u2Dy0HzSvpGs5dOkXM24DOd1UPytDLCRO92jX2vLA1rCS9
7Lv9drnYWm1+WlmPxiRAUT32oDPslPRf0/oU/4u6q87LLhC+75hAH3DFUq/y8q8iOvo74Il3N2tl
qeqq0HfGxRGDnSkUG9gxCm/2T74GAG7RXD+8OlFWo4+FUOaFr7RTC1xH1fGWh+RqHpqOP52NjYXn
1voXvrTH14jH8DvCKOFJn4gXo/3JfKMLpV8+39deEAo9xQ+Fn8vF6vCkXDtDn8ga5k88hSqN/HSN
x3lFDlQ6UUZd3k+fwS/+sox6VwTIdvZCWcwid2PWPyUW0NaMnFnJlt0oJKrP2bqnENUf6WY0kj6G
4lNU9gT5D2sRFSKKmw9ekL4VmN3gpyOqhYh19VN8H6R7WHXC0/5tvRDyzGfa+ayqOn6x2TnldvfH
2RA22ZNB4oukp3Pwpccf0K1F6grJU5AsdpGM1Wg1o+2undDmEvMeo/RK3IeLpUhTQCSGG5/I4xV2
spny7T6TqBLgn1zP26EWRMwpqtz9MF9CuJVXkJR2j89j+hfaI6PtaEhbZehLZU4cy5SydlF5GdNu
gwgdER8VdZUdwym3gAVx7J6lZndDhPh54nxvX5PsR6Z5sFXD2gZa4Yg3wK/VtLwCVVgsb9xSy91/
FeuamY0pypz7z9MbhPqZPVE7BkNxjE+unAaD474e+3+8+ENmFQWzJbW8GFf8WfMoNf83aj01wCSh
WWBbT9F81t5uiDFIazc/loOG4KzrAEphf4NV9esSec5+FpvrdechievC8lLbw3I11Zo5/D6mNE/W
zlqJFbVeY+s7QHa8AJnsa96o3jLFkxj76DNz8mlLRKI6jQinfejYJprnCoY1+91c91Lvu/bmxfps
NdTemMiIwwJOmyCq+SVAMJeJJr1eeZc7aJApe3kPLLmxW7LAe1I0TECBA+5V1CKHjAGdz0xb9yao
C5KZuPAWulo3furR1RrtowLuqOvURcN7JOVI4KgKE/2UWzQePb/mt70w89imlFYR0Yc14gn9HzR2
+O17XLaub+1uhfIuqQ+XJIO+b/1WtaaajX1N7aNRzHpWCRFBA3DrGC9N4O15cNUvIA2JzGd/HV1/
no891705NHTATcWmHs94ye0xgoTRO95PWuzm5EMb4xd6PjEUBS38auRvCgWtm9iV0qGg9DlpgP/Y
F0f/jPe6kYOfWCp8NvzUAb1UI967lIARHAnoylRiysJF3mV0KTAJ2FSpctG5ozQjA7oAw4S5k3I7
n+5Y1QEQLr8uNVcMIShtgyrtnetS5gJ7wOSXOhuutk4E1nsh+eKPrCPLuXjMLfRlXCzMcmJMhFrC
jpdSyFlMvPQJPyBUpKYLTNI/hgMxORhnhJQTRy3b8NGAPEspAZQot9c3h81tcLmuRVec4I0ldmMD
8Yypo9YM6Z7D91OkY2rAeMM8Q3VV9nyzrOs1zYdRfDd28GsY04XXzH/5EBdETlFkL1w4rQY75rdi
aPg5SDELQqMxgodGzUcFloTcE+pnt8OQAdajZtwGgvH4qodP5aLiAk0hVNJauujIWGIeqcJnCxxw
nX+XTrb1HVUL68JJ85lqmm/to1wRBAH01g8yrhYgq3YUllH2I31ERKmDI6hrDBS6zCyO/iPHdbaR
5vZSVHREwgx4mKp06cBmPjquLAvqYbAXyMM38Q3cnoitC12n/mE7ZgarlRTUY/Z6JpH9ZR4YVxT5
a8YFysoyORMiP4J0VwgFrrFgDvth2WhbtOInVFVCrrd8TmIBhYpubLDiPAi4IxjPkwUfFJs6ZJUC
iECP0JU0QMBbqHfoG8Ay9eMsNKmWOuhtRiO9wshCtCreceBes4rQrBG2GLF6GUg0HWqQ5w8CR6II
nGpLxNizTJ0JVYaXNg5UFkH1DGcBKRp8uC+58DUxFdHiXwU5s3CLqiZhROGSsjlebpFcmhiNcDZO
2ZcF46BgjgkHrfczLd6XaSqQB6NQb/GENPqjSyl4A9GQQ0MK2HvpwFLVCr8WnCaQupgtNLaqSFHg
xZu8iSGOy1qHAfQpQuT/ebbNcDN9rIG4yQbnU6XOgv0cGUEGC3pLvD6hoGpNgBpek1WPVR7UpfrL
9tUevxOnp8pF1rQErAMSdoI51PVq1q1jU7JO69fcVVF3LDJO5t9cLWOHc7vk4PFXkaF9jAqx5HuK
rzKglm0T2VZemFB+xQPHdLLsUw4ZiC5EiWfkhYuikj+bi6M/gwjQMIJTbaJ1nQl6sFqVQjXf2Zr3
FB2uoruTBGypk0+LPX1ElZFMhMjdYN1HerGGaICiqUwBYaspff61JW2z34FbzXeMpNwrc3mEYNRn
ddLU9h4wHt88Z29f+p+NnrOwNKQ0TNswQK/bztQSs0VcRjv9dqX9v+mZLb0v+6vEHy+ezJVI4x0y
hmlaVho5uLZBK9cQzhBZxQdgDJaMf9w+u2aNMOkC5a23wPb6pkmG6YBmiBIyjNb1MhGqRFCI8qrl
1S30E4mItJCMAVNGldGLhJ20cBhUf8ZsT4v0Xm7WI4T77qFTsaz5n0ATjTXuJCLm7y4J0HdPYpw8
uMNeXYSb84qiU1rylGlQCJtGZotn5cd/czxpASf8q6tgwH2C28uhzgQDxWGsEu6xew4HA5/vobD+
E5QDNw7TERwrJMUyYkuX4G43HBKr9JghHMSal+JUQ1sbkyOWD3z+NXdHcYQyEz/5jqH6u7cwgyzB
pavn+ybEEvCoulNfnbcMHXJAaaxTVBvUwoz+UGJQ+9+gW4qhrTvq73prmOEeEFoJMe3CUz32ZAzV
Gn9PCXzjEKOtknk6qh9bhuo/7/nM26GnnYrk9t7QaA+Sm/IdfsaNsa1WSCNaNP33imxN6dsWzKZc
mzGd0Zh0iLqaHMH/uIeXF9wQX8LUDYStSMP+nE0m82FW3EGFL9LRIWHjuP+JIWUK3T/1Wlh4B3TP
6UpTiPZfmSAlLti32bOyXNCwPfOOlKBx7xAeuJ/w97ngg53jZ0EFRGDyPuJVxCyVnUAZctO3/bo/
h9Ky55BfdNXtnQW2wFYcqz5tTB9ZW1bTks58iV5oMtxnrdbsTIDWbT3+FI2WoJDo0D+WW2qwJ5IY
3Z+pdmTMjLvWUwTyuf+vfcfXVoAXTKpi6iTcLbeMsaffADhGxSADkSZ9gJel5GTdaRM2deSBuF1Z
QC6z37K8BhW8qJBAye2SHdc/UkJy7Im/CdzXv0hMkrpCpxLIDVz80Rex+VkTWD8FpjnWDvbLKHDf
7QW40wm2syR4tomwo4s9RFsGP5md0zRse49PwDqFvgpflaPKMnuFsBcmRgrVHidfc5G/AjxBUUgs
vwxw2MI3OR0wB2TdVvgldwbpH7PIom2Yebigl/eKUtK2OBP74IpvAMjirAnFyi+anMiREN8cjUsV
rgic1JOV1j9XQevIJLv+7PHkKbfnD0yDTlOvGErc6L7u4jq+fdMM+aA7srzLGwAUQwuUrH4L3sp2
gFCQylFiYr6v1cEAnskdA0yI2nG3SGLM/koAgTf8DAGS9TZvQTDXT6Y496ei8fGUzJTYX3z9n5WC
FDITHSCN+rHvSc5e9ohRrzfjMNC/D4exumC/limHDUukeQN7+oRrulNgfs9fzuXVPYVTSSkxVdIf
nzacLgjdKNmI3fPdsAAhrqWxQkkh/2Cfs6juUh7hweBv2u27VmNdGvnyT/3FFw7SuTf4DswCsjFo
fiP8MlGj8TLQQo6eCcFpyBP2lrcBQ4x2lCs44IaGttPFcke7NNop+VIX4xvEd0zaq3QppXdmRAaT
/p4U5HkFhKY7/cqWycRWDMYD2Dlpigr1yXcYJxfHlNE+swsvz7Nummj2tCfLnZbiNZk3TGQ2Ts1H
RgzaW1W+EomnLQBWH+1R9nvps7SAvDuAcRIl0XiQOGv6uWUliwiGOkasIqPGE4JOI+yWKfbdZ1pj
sYxpThVf17/LZ6EATFkgNy52xdd0pv2qUgI0sEf8WCoPmO7uT2sjhYW2mNqLvfhHvTcWLebGp4js
TzhHht1EWQ38ruE/Fqp4KbDrBHhKG9WUSN99nayWt1gNy+YLLtrixV+6nw1+eZUELFlIQiEORq3V
X2BjEfNJeMpfwN+1NMBzacrNI/ikqmVae13JS30bUzCVX60aZbgnWwNdHRYCOB28oOvKPNXvmjZ7
AhCJkpYZxOqhQ2bDYc+WO/wsX7R67nELHz2tFKiXije6kLY7xora2qdvpoSS8sh9zNz31CjULe9s
hGAQpuoyTpT1IKfwOWUH3f+tWAVV+79PWW1ryNDW9i3147QjQLLQYr6h3ODqnUB4kBIVY6P5tEhP
/ybiVsiIDh4lQFVcbs4Vn9j1rK9YO95JkFCPg5wDWlXT8aEUzwhPM87Reg9w9Hcwao8+DJRSlVUS
gObEFQkOX2q4572chhoRSKBk5DlV+X2T1Yy+keu1y1GPAFHVbQqtM0xmf/7JnPtVdtuhuRlD8Nup
58KUwi0I2uzrs/DHSZStwflYoTSN+NDWoiT35y9Kp9ULq+ds1PtB7sug+/Rsr2OtsrqGX97fqxP7
g/azf4QSGCYiykjIihw/5jXBcCU+jLcFG9zp2tkZvyZeowXBvzUfxxD2Sarg/InlrQrngGDAEEfV
c13aroJ7VmOJAAA2qGJrDv/QzthvNExGUaTS+t41b+ZYhz/lH/vDOADkaLMaBTi1S6cs91/3Lz/2
d9flQX4tq+hxEk23oKvyvMYd4aql0S+QGKUI0RrirkKGScYhYXzvLPvzr0txFrW1enHU1T7aigFE
/eoDjIvVvD1O04xp+eNa0IJqXT/XXgI5li9GGd2LgCFywvCXXEKjKIEprMeOXkznVoACjMy8+IGS
UP2mgPNBZ1zX5hd4eb0ap+/h+OXAjuqlT18NebTBsazNt8H4cxcUwDDc5GQEz/DbT584IbTJBHhZ
0FkWP3rP0zmDmdHScrx4U/xt9nPe40Wgxm+vwt3mzLO30WYbSoE/MIVdTie/CGPUUCGYYd0g1odN
mnkr4pe44T1+I2x9/b6CIhx253XjYkdGr0OTScwBM2wC+Mt3WxoxR6DqPKez6YbFu3HLbaEYf+lZ
jHZ6IENpqElftoIGD6ZCnjlHFmitlLkuj2UfGf/fdYxJ85WCTT5WRsP3veKJk1R4whEV3mccOMP/
UBVd21UHUF2StX2Lp21AxGJYLtysQu9mTN91W8fQcirIldDXoyuF8FXGMRydkwdWVK+6FHz+tynV
O7n48LIqEkm9rGJnhBs1Qna+o2dtwXWihhGRpWQnn782fQ/5WvFuPdOgJilPwq9k3CVILM+iKC92
XIQwy0sutBlWrK9L/ZlRggO7tvYB1L/HH+0SVWprMAJctBYwllA6UoTA4B4ETBGUKFXwlc9Y4jN0
Wbt/CLT81E0alRlEzSlIFoL2nJ7x9jLC3hT/mmaQUIZXjFK8ELFQMrzpMxCazxkGvGc2GUDXerlg
Wb6197txci0KmYFd+93x4mBYbM3iLbLDbWFKdNiZmEGYiZiVS75i9nU+9sHJNjTnEdwSJLhOHc5J
i//3GST2ZrHEkbfj0o8gDo97A6kDRIVJByYjB94LPZFoN/CqeNc+v1t/kNZLb3bcn+5ZjHteGGUp
nxjR9vuWabeDKYAPSF7fZAvJ6BxyOV7TpXxTqOghIgoh9YLHI4g/qonNEsOXQeY8MMjt7rEnlPie
ypak2TfpAQDSnCMZfHSOt37SeMRLnqv2tAAvk/A3SzHLMZJmTjWcRgOQgendxymo9yYtRE5X5Zmd
bMM9ZQlqIQnqtJwgvnrhO5NKVB2QNsnZOoKXadFv1sS02FKA0ItGsilQy2Zufbm3WzbMrKhqD0H8
i3KgOtFfE0ZNSEerb1JYw7M39Xvzhr1JCJlQREUqzhfI8diKyUJwKUjxXr3QUQg0t8B+EjpKvcun
5KBmi6Ln8ksP0yJMCJ62JjcO7RPUUqpHrv9UFQUSMkmEm1bIx7C6DpmX9Dx3egNNNF+QoQB/aWQF
MbobnYPCvXRFhIqofp2S5sagPVJ/oftmjSaMPhwa2N1rqCDmjP4IcWPxFD7mi+xiiP+Cfj0WFCG3
1GVH/MHm72MkAqY8GmrMdSkMNB+5+TlHkM3A/yyIJSnF+nuGw45zoRqlWctVeDrfUmdkwfqyLpmH
bQD77N5VThNG3/hcxXkAJMSzbvD2VTLZ2pd8C9mH023j0vTHgzbtx7GXZArPnY1sSH4IxtRT4DkL
wFbHAShUOv31H5OfqsZgd+77Rr3QsSW7i4J//a8tZflpz2uAznAiwB8wriAmRSh3J32tGPfcstrk
2/hE/2pDCxPGgAM2Vy+wqtQMM9ib1SEp5LtuYduFn2xv/SxgqAwNXRU4uTWgep4zcwcaiGXY/8eV
rwFII82itszMd+6kURijRtfxj8cAnDc18R/a9sbmNzMM0YDF46td2ZKnOgn8kUTqVf9HXWvrKYDm
tm3+voV/mtWKhZmgAnM8FZj2h6HbE2/0frTlOXcakwIaQp19u+3SH3D91Zwt4Roz9z0JS5f4oq33
Ok1cz3ocATUozH/51CZ4gmg00byzsuPv3oXYFb/xwXVVXoymJiAX9KKUB1yc3KGu6WN2xiz25qpy
J/1RyDNGA7bfr9SaWvN+Nxmz93Tf0G8MlIbBK3WU4Fj8js6Q9NDarJaZmGE9IimYrqU+jLOoeLkM
GuyR+xSPAOc6VngF933LboV8D+Z2ETWXSl4IBy7csLDVmdheBHtFAlWG93pN7ZmPyyVK3RsGE2cR
LFHMJWqHd3MW7/irJ2Q/SYs30SyDwAbbHaySjX+KbFy6+9NWF0Pz3KIwJo2vwjEntz+bC39DVnNc
ljaVc/++763z43GeKJXuLFAcFyiAgoGS0L8SJtTjiRk6vNPss5sswyZOqyXwyhzdtYmhbLenRfB/
rHmJnH1VSh1NR8CFgVNHjsuaqGjNFWbkX+EKhT9KrUMXG563khFW8hWrIjBWzSVNp2g4LFy6y/Y9
uwyuNs+2qHsWB+bgxGu/mpPg5syjHUzIHNX93QyWXg5Wfqh9R+rHN9OlBKOth7KwgusEobr6ZIiw
UOLqi1eNQqLp04uO0CeeaIjTFQYr+CQlgagf3sGYcGVS6AQHzMrcBQ4ouaMRAxGss8XYeNuPP/Z2
Yw41kAbvlC6ITzZkr6M5fOdUidjB6+AaVknWsb/avfBga8ZjQl0/E4DffgVGHdjMIXX8JLJ8tbXL
sLW54KNfXh1+zg4gSZBsddkQpoP/6u4JZJ1V/3p5Tz1H8pO5HnE8lwTCMXakCry8UcrgO8GdJEWY
fLXiHkAbs1r9YMXS9qun+YqWsaLnjEdibghRt+T2j8/GQXUE40OEoHKSEAAe8pjj1I9xOT4Dq9l1
/dN+TeQhwMtmysyoHrN77wC1bbvHT8enaiiwg+p3qrOQfYNVPit4HuPvpgnJLFawLG/O0i6isl1J
UgZ8nWsG0hldHI+gSXLuA01WpPvFjhwuICHfRmGP+bNXZHSRbGlrZ4pJft1YioHp2eAgCjE49rQ0
ip4+axfFUtnsq4D5jIeBuacMWxDgRx/lyzbg5E5pxu7UT97Sx18qDjLp6g99u2jeUhlSvg0zuUl+
Kiu2ZZUw44NXvvrLKvWNnOaBVEGNgXsa2qCMJiYIcg2S2PaJ4dwxhYPqwaOCcbp8ddaCjTLrruS1
X4s6kKPyGwrlFUQVt36xkME4rcxl/t52HodMwZIGlusK5nD3LTtA8VVTqsEgOn9girIC1i4nDhDm
X0c1K3MPPA3jvSs372aV7vxfIF5mskEY92tXX8tcbs6vP/EDgxqCiYId8xEPNJZwr6tJpOwsYRLF
1UowR2l+yOJUFsN0RJ8Tmyem48IjqmZ+tDPenNGziXId8+xXJWJbW8I70YUiuKQ7sz0Cwkm+TLph
jcIL2uCTfzVDspZWzwve81s2IgIZb5LMZz66HR/vz0bJ82OH1Y0V+GlwBqcSK3qYVaEi/hyVsKwL
8qO0AmSeZ8WbIMaCOr4i2qYQXGNJex/QhoPD6KRh94uHjKgXm/ODYGUaWJ4KijOtJCcTsEf+lSZK
dYkwRfu+S/ekEyiJ5diWMEsOo9z5+MIGPJRog6fzilqfXgy+M2hng9M61TPtgoyZTCo8tDZ08QPo
AvLo3YyWdxlGq2WfZf4hHOqA2ZniG6bpSlXrMewRUKXiOLTVZvb+RrGdtgSv7lDmH15zSuvH+BDi
ZLKCrBiXndBM6+FIuL/FMFdvIXbUnYaqr4abGz5MDdiyZY4lN9w74c5qd1AMSxDlWYsgWXYXgp/s
BIR0tUPDB2194DrPe+AmRhgrfpJIaJl9z/p1cdP6mNGHlUHIArv5qPT3ATu3G2n6pcCzdPk6rdrK
SA0Uh/L2RXn0nGwE+lyUQVMBkElLynIo3hTFyVITdsV+Qmrh5Pty6vDtFsxhfn+qgu1EPeWs7VLv
tLv1Uv4sZuOO8L1AwpkLaIwcxyVtv/Y3f1xn0JmhMsk7/odw/l/uc+W0XRyE+eHaRq8Sn28cU290
DyGx6BdcCxu++Yl3Fr2xQF/3ioD7nGuYtu+QYK4a/hfpWB2o/AwJ6USR08O4BUELZXEYSaLlJUd7
pnWgUmbUBd1m+feiH1EjMfTSn9Wu9cU7o8ye7krgsSpMRMMObfPcN8/XeioL0cadiOsDWRkj+mS/
8AtKHon0QCmvKqV0drp9bRi7cv+IxKXCLn2GD1C8fznTA+n5lQTvdUBRiGOBCrFAszUeRhyAlBaW
n3OEpDgx0lDSCMHD0//9QnvwblYfoRQt51oqS1fU+ax01OySBBqOuo0pHIkJVOrE2vDNE7M0lTXJ
tNcP56KCA87DVaiZ711pt+cowCTzGJxUDz8ADHUJP1xyPsXfb2mAWEmzqTf45WZv9ZjtVDUxkaHu
QQY+ZzkmZYSLJ9f14I4T2Tvy+PyrW/KQHqgLwxvqTQ5MeL+HzQpc6sDj4CYZsKFN9KKLSoXFaE+R
QIQjDFMZ+zdiSibPX+3RM3+g/t58XEVSw5+s0870ZEDMkWFYrR7bYyfw4s3LbyVkEX3P2PVLSJND
bhIb9CPbfDr65D7imdiWmfTlSTN1dVZU5LIVJqcObnZm8l2XJ0K/bjxZKUJIW2UBX/uSCsyf6N0c
aeJJp8TnxSU0JVtM/Hiid08fZkLSWIa7jS2DJo4TACuQTxacDE7DWVelyVTKlEShe7F4OiFzNqOE
ty5yhryIouAyFC1P+85mEQnpcqNi8R6O0ARcLzQFjpluR+yjDLx7ivObTH6WkTcwEIahF+HRIXR6
mL3lBJ78DnWsHgVFPI3fyskhOHC+96MWyhTcB7+YWqzIDkOW6zM+JkZQOBKp+yMdkcee/Ye1OQuh
IO1+dbG5G3RBGodqDT2GVlIYrVjYIqoM4cw5ciceX2so3OLKG9pn27PRfdAp/xKA/HmQ8/VMd8Zm
o8daFVIF35XGfZELBLITbPEgzNIlQHenO494xgJsapQO73kj1ULMC6KeEqEHdSozFGQtDWz+ukcG
Cs3esf0EgKyGWaejRRRtTCK6+g/JO8Lw5lSWNlD0T4kMGYqZzRvXYakE3LD+GUXaO/D5oNTHsHIO
EXlq3etWcamBZSW296ItZyv4b7xowXkOVubUtGH/oiPUZ4ySnj9B7FbWGinQVBCmetnpbf8gVnpq
1O7KVTHuXXH5OFiKuBY5X8MiYaEEd0iKNRqsjl1F9Tni7R4erXikW2LLA1uDCEUWJnprnwBvjkjb
qXE1/XDtt1QH4BLTb7tYSZXfgdriQodq51XPmAuCkCXuLurr3FaN8vAQod6aKP1y/Ku0mGTMG1WY
6qxFEPJ7nxpMyYRwA96m4rkE20teg4Mc4pmR9T/Oa/8PDrsM2tM6pAVPTdrEDlYAj3mhsMLHnUmW
STr9Onkbf4iz6hkZD8y/w87hZZcAK3eGpcwqo1IuX0nkoAhptDjXNYXlCXyhWADtZ9hxW24OjkZt
AvfkT9q/cv6zufMNEw2EJGz5SWcEo6rZyLi416KoYG0lOh0ayLbFe7k1IVOyAwjhXVOgIkw7fTvX
noNpKa5JfRrWfmGSC80a++HrnkVrcI47SrfPmigoBkdLDU/DKJpZPsjfRw+59vkb/4K6byVv8X1/
36DHv565idG3wQUVN5wuWDayq0fQisfN4g/wS9kalKtlfZoRiZMOxSU8liv56hEZQhcI87ghKoTB
2/KuS+WerFbFiiZMmW6C2YbHtORstlYFcCvCo8qcN5FauuMloFwygL+xyWyTysvJURc8oNM5MnKW
mhTsH3lS+UNGT6Hld9oy3AJlWhI7R65+JorRBnu0lDReHCqu8U08i5QU6+5z4noklkjIl2aSxhqR
RUlIQVvrFUENLlKkRCSNtq92mnKv1f1vxjslvAOcjBUqGjKsNQzHxT8wkxY9v+doz3pE4ULblvn/
adRRM0/JvlRiVtSrWicmN0zXXSsYqIrEjiy08Hsx0511wbERs2BBsIFt9Q0vp98oP5c/3+8EWQMy
5VhQMgImEU7CudaRyi2VY43wjdPJzaTotv385j9b6xcA7cThszrkeET10iS+awIExciVwGWSJV+n
CAfQ2TkD5C7JHq3A7YN3sVIaXoYI8Y5zS3g1y6nrMd+BFfCW3U9Vqv75ATmT8n/f7K3N6/WwozA/
+FVLQZlq3H9tn4LG4m1VjbWFzFukOkQRIenJ40mj0SCCAJWJCLFmBmaIBM5uoQf01+fMHtVrUYm7
hLb6iWCu37bD13V8LFArtJcS5WMwCL1smeF9FS/9UsZnK5FIW2vv9tQxG0k8E8AiA2VgYY1lU9Lq
uaYzFomF9qph3vCX1rWVL0ZWY19FXUxghz+7YpDZrA7+lsahx/b0/ZSHvM0xaB6gat9t2ylo11Qd
/SlT7wJ8Ks0iXCvSvuGQ7dUgg079hoyZzRV9jsK0vjhRJo5+4qEwgTNvLcN+TZBAhoAVzi7iDKSY
vNc8w8fiEqlP53PXOEztCueSs/anzQyoSifzp8PVQs9sqlJPWCO5WqYLeFYpzzidNVowXyUeWm9f
6E6ntfCt2BnDEMJh3C+A/XeS8tcTKURm9BN0rN6UE551JuGvKcKqMJZvmgNiPxvIWggEGAyo/fL0
IOyi5BfqwumUXfH6+ir48/DOveKXOKSC+nWXv6bo2BtM8QTBcjLrRcG1Cex8RzxGibnEd61Jnn63
RTIStf54oSZyVXNVEOLQZvY6rr70Fr9F5nR/NDiMqpRSSis7lJZpbPe/s2MxNsidfTgctiiy9Sou
rBfh+9djCPc+P0Kg9dhIBE39MFlrggr5W5F6ylSMcqp0Pk9EnTAWfWpVGR1DyGUm2aVcQqN4lEnb
StOrHdCsHhBAJlxqJzHF1vKN6xugb7pZaO2GYvMj3Olnf3ykj5I6ujiBFKYqQY/cuWxftx4cjnMD
USzztlfM1De7rexKGm/0LastTclWr9bYs5xIV2KS5U/9LIE3/Td1oDNXkGcD3LFniu4LzZNMm0p+
CSjdES0jZLCcwGyWz72JemsK4eJlIZCLAWvsr0Z48DZ+BA9nstFKDRoyOSrUTkimsC+rZ2PQu0FC
8r0/A+vesc+nv439McBwDnEamCTi/44WjYIg/zUi5UaaN6jEUBTvdahYrUD60kvZKF48sQS34qbe
/r/gd9TbkCJome854xN6n+4pc4IJX++ua2uVgdgby1Dgz8IywJf4wwrZkybWumKSBjCHjy5MHxEb
YpdzHG3qg34VHFup4l8bCgxxEmNMR6qGUnuqc16JJXQ2IX2DWkC0ujYKUuJEQD/KYF973I0i+2RP
TkmOOdePSIYNPKwSgGpEa1csApiBELGE6R6xVtECvtZ6QnT60Rtszeu3Pnw1HnLQ6Ykve9KrTTQY
qRA9al9yoWE53G1XkoVx4e/InR3eIUiRsf5lFM1PbgtlaXzBtx3zRk/IDOHgvEI0u1O8sjfXqWeN
oPfr4w7DQ7cmAywf/9BYTrWqqZY/E4IGHlyEJl+vrdq5Pt64fO2QMH5A+Q2IvyZbcH9QwtXH0ohX
SDR+HIq5CTwMjhQbD7cg1XsAsm5ta1hIG7zFZQB4r8qlH8AdLTYDiyLCR9ZBKGMsizpOMzj9piWy
ValpzTFSBO3eMZN7yG+cTMHeuQTZDKApcxb/3moNHd1+T8WEioq0BpLixXRP+uirdfmGLBqNETgl
2HrvBpZrnkc0s3BiDu/h3Do6wbJhBg8S6ly6QWl0VPfx6+597ct9SblMWdYK25WY2I4ac+WJfyZc
UEHIsJSRZhpp7qm3ISYBZ+kY+qG3uaBLGoleg6VRxsMz3YtRYCuwkpE3kiYYtffgbh7vi7ZabJQd
MMCu22PVSznF82sTiIGPbf3zXt6PR7m1+FhOmK+XTWW7LPe28idZS1AT3kf7RmABnCDa+p/mzcWY
dsWZSA1njSnWxUw0CRc/wHKSOeHVnDCGUgnDl2jaNPcrU6r0yQhfR3w5flgXIbZj2//9mFAE1vpX
6unNrvVz73ktpOKXEuG+1KDI940F4eb1HnfEPQde3LA7ZevLY4FLy//HFp12jNBfBOu505djEtOH
CB6+oSTdR6CTgfrzQLkluhuZyc8NuBaHj+L/hG+a0UFh63LFDa8rXqmnOKxH8bKT2pv1JGao7Q6q
IYrh4ECJPtrhs39OQTuQqXUOKFjxCDHuV5FSbqa5wOLPbNE1sayYv6ISJxvyOd7GEaLwaHoaDwBq
7S2saQg0LtRvGD8zhozbTwGliNQPwu1cUhIaF5fkrruByyKM7x4+DPuAYcmo6DtukK2OeuVytbWw
EGhWe+j9kWS4PQKeqt9UIvnNvhpEEAJtSVzoXNbFHfQbM+kx9Ml515ejceg9eAoK7UCUI26c9rOG
rmNsC8QKGEz+iWzL6EqTscX9ndLW9YaE/5drXi5yo5SzHp1O8rZcJ6cr9Ar58xpp65q8CtVhEhIf
xZtmR2uM2Yvpia6URtD2yYzGlNc+BypUnkON10Dx99mqo7gE+5p1COTlcGjaiCS4uAVtTbk3DWBY
QXPun4uLQTC+bxhAiOe0H+arMIcZ24jVdeBynjHObb8SNa4QVYjr83kld2iHI9OnTtTN811Farl4
HJlkuRrvCI53vtfUeDjKrZJOnP6cLEgLNrGhdibVe+bVSzFMazcHQtQuQSLE/5hfiWn5ICtNXRtn
+l7ukUBFbwSf0PXguGmCk63AIv7lP5EsAwq7Hq/69tw9niND99cUnYbZV1jQJbUuAbVV9+HA2XHJ
V5tqB+igUkqd6VqmqKxyv699Sdd+o7hjIfeyKhTT/OI8Bsbefp9U1lmehXhADHbJ3pQQ4JARLDPz
djU+HC7QJFGKzyuyz8q3+FfS66hvDYU1K3Vpe1bA9Rk8ebKbpbgwEAUWdOPC8sGxKbyDmb0Jq6Z9
S4VbBJxDfN+TwWm+FjNjMHtztFSxMjYd7m/ih42d8XqrltEb7MCj4kJ5v2H3XDx/SLoI1VPdjCKi
L4UW0EJ1yyxtnHfnmvsROPdj42Mfhyj3i64nOJwiWYzV2QcefyFnawh9HSuWprYnJ6ZpjJUaDzcw
5ebIxSwXNOPtL0UKv2rYQMuTAHXzXw09xY4HspOGoSBvr7hbbOR1hWpiQgt5VWgUnUXTDsI5R3HL
07g2Xv4n+4kvIVAZWKbNN8WOLontpe9hXFxAlda58W/p89fStY8dMzywPyL9+8DMDhJkRcHR9hjj
igTi7kO1kp/1LEI2mW9dgcHxX/kdnez+gKaO8ew9nUXY97bMqhlGqVVN4ujXEH6uo4PNJqvF2X9W
TyMqE9mRYVrXXnkvIMUJIBo+Z2NDwsfSgNRAvzhDtyPoZNnYy2UrKZDHEuDzW6dM6M7eCLpR5X0K
mb8nbYnGhLODGDQo6FP6J7zLueh2TBLxq62q9YQ1rwTta+mNoO/xD1wliWP62H6sx8GDodqR0C2x
riAOw4oJOe8oVHNrsHjtG/GiTWj+CaPotE90MlbCaMueombQuuFh6BL6R28/rhCf4XwV4gzNY+0H
qdt1WratBFO2zNY+46ffeKyQL3nua/9pt26SJiRQqC3UvIG9TPwN3v/1VIBOP/mAKlM9UAszH5Uf
z/ujlr6MnjqlLeiKurPkWtSvDxu9HmDbW4N+fheG1c2lBaYsxXH5mGP+MJVOzqf+28hruq+dckN3
YPSI82o64w0P/YuvXEzRidgYmFlA+fw/2nzI7Gqptpw+JEiA/Pok7InvlrCC+UI4u3DOy9QOWt5O
mj/wjwzY16Cc8KYDZZeGSl8vtlpBR2QXqIOrMf9gmj0w2gQqrqwvblw/tthswQ0dSVFGQuLZOgAf
Xd2U0/BBYL97ttb+xN/5fvsgws6zlq9HPAp4S2ck5jxA6j31JW1YSu+w/FfWUVI3diyL05pZZ4ir
PR1j1+AfTSEhtIe6NtM4cq+RICht6VWKC4kOF86cZZaoulNVgsiIFzRr3W4AhhpIhQUp7Bgw+RSe
Y5WW+H8Q0hpS0VGpSMuMTkCRnWVxQg3G9EaWJ30vAMM6KTnoN0D37gjCAGJ6LY9jfWki9kK8wmu1
P1ODziHImkvYwnl/d3/uSSWx9ASeuXIVLjo3oz4sq12lIGu+VsHd6shyF3QmYQ9a69iXVdd1HOUi
1s4m8qD+W7sx2UnACM7ifWOekvToi/VyE3v3kwErMNN5uKaovDRqebJ456nS3EdbWPJaesRZzhcE
gOUUELEG0mPcLn03gKao0UhtqZ52ykryGDy6NWJ/gTCry6tAik479rva/AKjqBxCKje5fu0lQep3
w5WCxY4uDCwBr2/W43fFqipInzvQWbJMA/nrrGS3DbRdNYg5FkwA0IYfyB7SVXagqZuFUs+UVPTV
vdLUSDcoNLQIjl9DQMBoXNTZnTCtaSEZqqIAg0aqu2jSX+xWKCETeTYGknMpI1SyrTdlX/62wuVV
VyzPD/sJYhnXa7GdBFPR9dTVHjb5Jtz7C5QjHkseRnmUZpgHKBv7RaA3DfpDzgwDteCUqZlCLgUa
x6guiOKPmY4xAZcVY4X+XJGADkLbd+QhdYeDzSSFPWxRhlfnATGc0DyXnMNBIPX4yQJQO1MCM7MY
14JddJGVgFmHFKNsoAV0c9zbnCyn7i9oPijxGJ3RAy6ATtbSXXpEVJ3/yV0dAYAimcLu8VWKJnRR
tujfALnLNs++czLCh5WZXAvit9TELgiYuSl3J1zrs/pJHKiaG2HL1qBo0T6mPCWXX95PhJ9y6G8K
AhyjMPUda5YdeoQdfSNSpPSRi3l64B1/jhGjRqZ1goT7QX+8KPY63BcnDfRBPb9zrPna3+vDNToW
mW+QrXXfC9iwxgfCmUy8PYiKQiQwij4QXTuZT2nl5mKnyMzYgDZ5zAyT6vc8ovI1qC6vGbxMTQtz
bQ3MD1ir9viPuvROohtmE3NseD7KzeKbcFqQcRnGhSIHJwpHbVuaTo0IPgj0hj9F+2f8LlzMZAwv
8OtJpz5UVxJWBWYUjRNFiHBXbfJA7AsYEJqiQowsrmS5jfzJAxYU5eIaa/6IJ62QCMjp9qR278ya
VoOBlatD67mgGi+fStXBZ+jrQKrBUZ+jOJjHzEniVyOjgE+oiRPX+SNNNQ3d58B9Qy49PvHJewWy
5GA2T28sdm7by7ZztbmNMGKh4joVVjcp2ZuP9eK7saBy6Ptp4KrAqkDj74NmvAdBfPINaG3pSYOA
sd36Kh2GgnD2OMCAePAFoj8izdYe90JS7SWaJXgKcl4TgIxEj4+OZvXdw1r4oTwTF00wiGKhBxqz
EjoxmxaUxcsRDEMr+2eVfeY8qOsJK3re7u7LgSFiR/pNbd1XiA4aSkiB6wjjPeb2nFVxouk+VWeE
TTQjk4KbTwWja0F7N40JCs2ADxOx+3Bkc6ZEHx2uQs7sV9MgDt8WlLjH63/y+c7T8Ic4BSbjPBwg
KLAyXmOTZyH7fbZcS8r6wUx8eTReRDIlwA8etsyfB8Or0fLs1kkYgK6j2onCPLAD24bLtBbxC+yh
550h3Rxm9FjLGGByG3d93KdRNBCaepsH4BTEsffnUAqNhyB4bGKABOBJjY7iMKLaVrlSUppKHsr+
YOGNj4wKJh7LqJOh8wyAAzEsFGFRz7rAHYYMiW2SCvXv49eGhbV/TK0plmB14fCk87cP5+PIo0UH
fUNP+cvoDv0aLmfnagS9JxSALBFQKCRFG8m7+hXHYNT3se8eoqnTllMSzue6Oh3L3RL0XKdWSKGS
fbH6WKFwvTdqCY6KnTBdLz9TemgdoaIQvix290IXMZOazrSFvJj8Cyq1CvuoHMJGFn8kTBly7VVR
GqZWrGbYtqCugQdG+xCCjKzCaBQVZyFjWqNJ+RCDhPvhyiDQBQDkiRu1zInNT6gd3QipzGB54Wsg
oPjbkOax85mjFUUqQajBJWTss1X6GazLC32XsQmeLxvbGofK3ucGpvCTyaQXxxSfzxalk3uNDzho
UD8UvPxQ0hWQNUgwCwZzOzdlfzA7FTCfCZ1ncU2q8L1MSlc8zi5EjMlUKhagFQam/0rnywqVq27r
5Jpy3qgfRPZY13Cl77aRCsAkPLnvSiJYOcvGWoGP6Jos7skJfgIIqGy7ix01/jVLPaRfDJJrfUBo
Jilw3TWcfCRYQ2iV6wHvzs/9lR8q6k7WbxfiCCKs5+Pe6bibt3gICkkPtzPR8Jd+wFwC29i4QQ4K
VwdDdIzuT1hPfZZtNePogDq9dQ1Gjca8EkN4jUZrJJMp1H+97IyWMzaqb6+SyJ7Yks260foXcI0/
bH2CXlgQwWIPd5ECHFawAP6eZS3pMYeSEeR7G+hMaOeDUsRrB44RmK9R+G7bQAGN6AqT2d+uu6eL
7fPDIiarFhjAn7TvkCj+ZOYOB2rRbEWewjx8ugJ+pm02Sg+yuhp4GE6qOo0cZe/bOeus+Awrcsgf
xaiXpz600dnO2zDy5TdwB3PUrPl/mAYFO5wjdZWWle3N66G+oyUcnHOn8tMMjCMceWJXIgsCvcGk
jGkhEfEUQkWb+AIV+Z8ChKB/PzVHaf5hqE0m8UmZys1DjMeSf+ojRzG2R/R7zenAmkrejzCwLx3T
p/3t6X5Jvh8KP3CVZpr/XDk0DAXViiznVtHnDup3FangrCHku6cGjPqy9S7oEz1LNqjdSf5sbdY7
70eoc+kfluXYoeLsfvKDlLkWopSeLqZ3+JjpqCDxdFabB0eIJvo0muVt1jCrioP+UjWwi1IoGO6c
9ZOKT4RqwHAo2NL2LlDkI4wy/DrQucZ+fzPZ/ocZi3i53lCaLAaqhMsbokqs17T5ASnfIg0z9Nei
JbUBZqeNyqvjYh7jxltnTzFpq464RUoAKcK/tE8XS37SqTo9aWH6qOw8EONMlZgbX2P4nwcoCbgV
STFJGdotEdiJgaHNkMAWt9z4dVhnKJgjsv35xGjNu+4rCDoGtXNz9MZnsY+0afyb/EwIGj18QkJC
tYS46ud/sckUXVG1TQxEY3fYrm+pSTy85tdIt0im7p5unFUXVEN+4aXr6yPcY+8oKB4n/TvnUVP7
FqTmztywh3oaQAh5bIhARx5MUJ+OvRnhx0eWyylKTvfvKle31JdK8XuD7HiAaWs6yZhtngqAHQas
QYoAt0J7kaATwfd5U40eoKp4tL3UkU76Ry1gfHKfZCp7KK8VOiGwPDdltN0Vh9YPbvqPrmi4xWC/
qz+4rYSbpkYwQelanGEXMNPeFXEZIFuxyV51LnvkB5PLh4cHx/10PX2F+RrYoQvG9uu+BQ2tBruz
JvS1uwRkel2LOUn1ASwgOi+99/M2gNtX1HtmCftCJWE/s9eV1YTw9nte+JrTi0AC96GdIELwixDE
Aha+OwSHpAtjb/mijRDST9aGLV9zNlJZLBa8S8Jp+kFhXdM9HmfVnt+Rgb/b7+am93qZjFzuN7Bg
49sPjzARKDMRZ+5NZoWTdoup0NHSDe9MBYAYq3EbA3W+MKy/0jftyVYZLMmNuxE9zeJuS+CC5mq3
AkknSECbWxhiqF9+2p9QOnU3Ah0K0wgZbYTC45Y+MstB+yYjtZsaCYJFI7tken2dM4ZwSkL+JdB4
cSaa8Xv6LZONN0/PGwihgDaHkQsBfSixZ0PmRKBBJZ4qA4bpsqBzfkyRkqMSj7KIvvv03gH3PR9y
taqqC0oohJYvw1WPoypskq22aPz9oS1aWZnPpA9diAEyh9UReuOxW6EvT11HUiGlU3COQZrjxKt4
LHproVnKvoQ1BCCovH/w9EUHglHTtoLxMrSs/u9XGzidZJYve2k7NS5q9ifSchzwHp+uL+Ek1xbM
0g/RvGMEi5WKi2UhXHg9XgyKI/x+/fhElgj3DIxClXQ8cqH0kJPQIadVal6AxtR9+VYgrbeT3VxH
YrlXfm/I+P5/ZC8G9Afc5vVBX32IxvsKS6H9AcuMs/pcwq3S92VyI0AqEUvBrhyWe1/9ujuNtXA/
HWliANMCOOH2vX6zqFXcYoqGLOblpT1kPo0LBP1tcB96+/s5lXjfCKxj1hkA+Sb1lrjTTSx5/z3n
s9XWxYRjWmVL+D+FtQpmtFDqXRTw9nkat22uuH+qNUaHmvElpeuf/2kYYF2AMlPWwm2bfrorBVlY
nj9p+YsHiX1YoFJ6NwlIA5wpuaLQx0g0gDUc3dFZ6uwFO8OZCjP3pTOJ0H4hTl8I4FS/B/jpFo4n
YidJkDK2Wjb87q1EdYTq7v7LdjNbHx6oCkYU7mdTBl9qQ7mCUsHCr5v9ncZhFRSmsY6KdrTC6Ks4
BM5BtjYNzdMWqNdxwa8RGOxZIb1emYbuvHfn8qQ8KJfd9j0xvtmmmBNbNXs8zNwl5sDYZxkQzDnc
svSla3JmyGBH0aNHH4oYXKFqgsa/tffkMKSyzD8NDGBDHNe0nELmxc4lJb0lxVTAKZZPKOoMY/xZ
rCgd2ZgN6nveIi24mH9hhnCrQ/zxYLBfihOLwobFL0M7ToOZDvpLUpb5rfOnnto3H+JRFyA08pN1
FOKcshEqocAuqv4CmAsA1VDHGYA3PxjUR15fPszl1gPvpbE87t2Q4nmVyzuLzpP9km35auhoyxwb
NSV7XFJE4OSFEtSSp7exatil5t416oYD1tntJqmPP+vCno6gZIvM4V8wIkFSqfBgKTKjR42pVBkN
8aVxaSgItQ/beh0lUD6Y73ChPyD7uZwOirojiQRdSGY8j27Udw7pX4qck7cnjb5n1+D0yjeGL4Pb
l/oGd1gKImJXIXOAhPAudqA6CL0S8+emFHVMzb9yc9fz7zBfCoMBB5Wh6Si7sk7NdWq3i0mekv4u
64O4OEmgJbPyU1T44clz+wyLdNBEIcf2t86/CaVBmriwHr9YJmpvpfzKeBwQobpi380/cN/Bt1Fu
iPUnEqfp+/MOeiEklugK8yEtINFAlMERZgsI69uCNbW9HQYtljkT8vKOBH/HpOySy/nrw8jrHadz
Q/ELgB+LhKo+6Wnex12Phppej8YDXAq6MDunxyfCSSkEcWgAgBwmNWcUSZ911RT4shMscp15IGpX
BPh6LNwdfJb4Itcg1pJTtZISM4ZvwHJfvBo3ASa5aAqsdR4mzs7pO6Z71Z0VaGEnpBNSzGlOft1I
rAHjW565S/GiUNvm+f7YwUfQ1KWIR/wbjY2GDc0ysjmm5AzKp1gDgcUxMo0kGyeKcNTB/u9gTzUC
6WT7i2PUry/WPBE+HsmXGXc3UwSk46Ni1Z11pYUwddkQxiZ3Hdbu4X/3Y/oUs6bK8RtlvEFK+V7e
l18NZP4eog1Mzp1+0VMeSGyX/x6ytGMmauyaZtF2yfktIBAi9fj8ppfMB/IgRZfqLqQfvFoQP1dt
FHJF/Wdqc6qcXjpslNLuChDL/UOml2vMN/EPgUDgJEPTjdA3Msibwv9dSIfFs0hZM2MKMPcABP0L
dOkbg6iTgSNke0YDsTB4EE88WK903fmMvr5hNZQnHip32329VeyHKuW96h+Tw6fZ2iEVBty5R0Nd
KP4ldzMz4QLIaK7oiyj8soQVruRMbT07POQwmmCWXIpNWPGhLaZsCWnf8bf1yV5jKYIdtEjMOmO4
OGFZetOLTcQ8nAK+06fNbO+5iOqptww0/oSZ5kOFf0l69qkIesp2eNzBhG6ijJT2Qvp9k/MnxhiJ
ElSUC2OrNanXJOilA7x+MGuWlxfGXMBoH/899bl80JViNOe9EhMVWQcvjpCCpOELFQgYazAozG8y
alFYE7SlvaV6ucRPcyALOqvRlqArbxchi7/7gvhuhsEXA2EKBl8sey+pZqaw8jATu5s8W4pghr+j
gcVjZumJL9bkmcw38FwcjCK/AD1soaJ+nP9Of5r9EbFScxEZOnKhHE0Hv0vMfbucTm1Q5xbcE4DI
crz+hQ0F0JJzeYOeIYi6Y3DgMs37Mv4ZoLXg6a+gAvYq6jxrc27lPVb3veJ0osDAf3W7p1iFfDLx
UEg1F2WjNxF5VeX/vXViKwoMmkqQZmPDnfdK9XnujuTSIAtdOWiZxBAe4mN8LLfN0y9Qt3d7MPuM
5WozcDSBg3cUCEaABpCsZWHbNz+HMWAmSwBm+lJj3mr/GQcKIu4MPYqWAjEnU/CSVWPk6rClf+w9
8g78Oti5vXyDL98wZOzZvQjM3LdbwuX90KFxGSdHSe2id9HghLZmWPuLbMOVbvEroyQXgK2ELA2O
n/I/KiPcgHVTulDOZkUVCRJVoMVys/4KTKWQEPDY7f3mkziA1yCXX5hCd54BqPKJu8YDzDoTLntE
8ghfQtZC0sCN8I1BP/QOEP0ewkuqtaLF+Kh7nP6OAnn06VfGSmarSsUgnTKJEdi+VJdc/8onjMEe
/kNayVtWRPo4ZYH99wnOxWSPg/KMvfCiXo+aPnLAaXmjPAxoxXCWwe8/FPa4amcwIWTS59l2kiRk
qbuZEvt6iPe7xSQGyEY6SL8T9HoAV4czg3NXntJ7JuwbmZFDmoKwdNb1lLI1KljJE4ISQCdQHzs7
sZnmyzMYfUHWNqESyNE9FCx2gkXTN9UJarsrau8eMOsaCqJVwD9FJPSnLT3YF/qUHjkHbZWEuyx4
08qPUVzI6jvISvDBzlz0azU16zzhcZFnxSS1t0jLML8EOUbL4nr6jaYuBFm3weccaVbSAmsHFx9o
wnu5CrN8AWsmUJ7DMAOJYmacTMLnlIy+FqHijY419KFuJ7kf51JEUBgfsr11izbLJpWrV00O5XW+
MCma0q5NOrmLmiVHh6FkukNcI+YTGE7xVno7sp+ntaRE4kMTFfwsPlDGx1kfCPaosGmtMRaCaDZx
by1WBwDcp/QxiHNEirPtQAFl9yEf/qrBTtewy7KG/+2F70UVTYYqSKeZZGnYd0lxtqNEIUyAqBpM
r4FsqFpy/C91Auy3ZKM0n8JVyTeCezwOpNth060JaXXXDyHVEc15rB/tpb6M4lRNKI08H8gkoWYQ
FS399huNhvMr4ADyR+jOmKrbzUnLWPhlcurqRJbrG3+xVK1YZDvAhIBwdhy1LXWrUsgfqx4ZeH/C
KyjgRk6hkCYpt4IG3rjj18UMoQdiOpuE7epLZone7+sUBA7NZWwsbQNnCEqRKX1lVJk58B6b4Ds1
p+ncECrPFtKd8n/tp4WkAkhZOANb0aP3Ajun8l48k/Ln/TY6yl5DMxhpCR1/Qq9PXAJJoxYnApYD
wWK2AGeUvVTqli/WDxrX/aHbrKV+kn0jeTATbCa+6inJMyTVzTNyF0PInEyMAv2M2GDZ04xNYZps
4X+8KK0GtLjOVey645Tgqj+sTazr0U0Y4jZ9ME1PqUxG0jYgMVbTdRpeEqG3S/mAouIe6MBSAvsd
vitIFHVKW389NagjV80uYDN9LTZ2BCUIIWdLqn4i+n4eaYn1c6iMaeSi3m1FsTE9vXh9Oyu/Co6D
pfXiZzoA2XhFQ11F2xc3Zl0wc9ZKwoTjjSFjUzO7GZ3AqSLWUcihHMi9r53YBlXsg+Qzxf+RSjGu
JtmwfLblrZzWePSFdhFJlb+dJkSjf9Uv9bNvHeg9utWEfddrfFLXrVIqPVZLNXv/9vPbpE9z+YOF
Eu67kFZDY+L+/IDAMni7KRCfleILCUdqb7L8Tt8hl8w+4hP6UXqRm/KQHFmGWpI4MfhHIkPkALvR
7jUD/DDIn4HZ3uMJYXacz7mYyIukv3BpnPLz2r9qEW0VKRGsJBJ1R18UnOEd2yq8FIurCHsFT+vE
+Hia+Jhaeg9wp1P16G88E9UTMyoR/c6A8rpfBOr8XAHIb/zH0h0t9ADiYHNBqFT7vDfUrsm01IIn
4YFP4neu+G3mDecioKbHhwuJNrbWxX4fuW33LGVh9Ut9aisVlaOKZOjqTr0Qv67SbpvcUs8CwmnT
mhlmNPylKgsXGMVGMvbpdn/ebqkUE8vT0KIhesIatWKJZcqWFmem6tflyVaS+WVIVX5iHySrDlW6
h/A3k1llMo39HqtE4H9ezH5c+5VLmjChm8J8f98V6vh0r/gSwrY0o7C2+gE9NU5TriSKr3QMg5SP
kAzgaa6rqoQYPwyZ2sCz1a5rJcHYThhhDjHXgCpVrb8uX6HRxrbxvnj8fh99QZ/sR/JCOdod3c5M
CKCtG+ZOLvQVQMCaH4XqEdf5nB68JwmHC81wvAzUOPZFQxgeGI2l9cYwqiQYLo6wzy4NeH0gTt7V
Kr6sCOBJYtvhw6Vqasx6w9F+RIsRc9TgrOpay0frebjzdr8t5OEgXgH+49/BlcvIAKy5ZYc8iQSQ
5IWTimkukyi6EHjuHZJat5FaQTdm92oQjol2YvcdoMy5XImWakZXHkFu2ji2huoiUJeKXMjsj9/O
pWotxEe4t5S8pH0SPaAVioclJ4mCWF8S+Qx8UvxS9pJoyBhDo7txwWat85m/eJZgasnb+DHMG5+U
mX0mXKojUCzG3hh5TzsQk1D4bXRc27+mG1eb1C2o7eb78YkPnI7rS4/y/dGV/F1WwKeai6cbfFna
bgX1nrbsRndFttNdBoqUSXTx4P6TSHgEZ6McyGvVydWGBCIfLtnlsjjzPp/v7vxIhbJTyNeAJ/6S
8xNJcllxwgX9rBcBEkJ1V5/8uEOYiBUVnG8P8uTqSeRzAn1yCZJK0FeXTaI19vlegJ/qWLqQgkZE
itYrEtmCz56BO4L7GhwcfWffgv3+CtUaQAEXHqgBaPTgHWuvQiQCS0fReIi687A6OQK7sOLVBvP6
zoxuvV9jBbSKsK+L/19i9W7/UcGFJSDT+SfxjZoBVBWsxexvf339nnZSQLQPNjMSMayNnp5O8GXN
g4Z4AyKms3U5cngydscxnGtVzckIPHmsZmx7SX2zp4cbTOvKzdQ9mH6WK2Pz0XVHnVfQ2TNRRCDS
U8HFZM4lp2d8zqS3bdJxr+kEHWc0F2B84p1tsAryABasztozBfzmB19qRb1WOFcoEVTn/nibuDSz
UNg6tYylQPchMMO0FGFbO4mrJYy9RWba/ndx+hlid0hurIh0eUk7P47CxzCd58sc8+r/R1pk2ZCd
eRt2ujix3a1lbamu/O2lGcbMIvlx012kBWER1Ke1s8HcTwlL+X3fLQ8pxIgV0LdxeE5oc4wt3mfL
849rWMULxn9EgcIHK4H+WbKTnFC+qIuSAFijUXaOWRDnEXPX29LJkdcGXLcyjptDP0tag5IpuAKV
iNUUHCd60rh6OYLaOQ+kgjVK5+neZFseHyv4B5/Tg9lR3e8cNPEWDjN+QK23xR/ysN6IHdAKnTSJ
RRQnHGHtYCZB9WQZB3SUuOXzFaYP55DUrLi/coAZRk4hAooqJNN+MEtTCuKKrLezo5J0sRrDMUb7
qqmiPqp4XrQ5vxKbCX8rFGx0GETGM4EfZy8WR3efMcyvt2UY9rHgkfJbd7EOZSVnmD6EMrn2qsiS
X0d0NfNtQ5/xb0rb0eb8UdxOzHG4y3SZTBxTLF0S8fkcZki0IGum4b0SDFqLw/xawkeFcb8bf2jM
Hz1Q0aa62uCOIV6O/zVumtIEVhrL1LEpUxgJs6EiEwuw4mXlUaRBee1+Glm5V/BbULwLI3Y9L+jV
/tT0rf/3Ccyzx6ONn63zRj7DBd5E2gD4E7nkrubbAshCY4t5uOu9hCk+k5Awsga9VxbR/OXc9atz
YlQpu7YOTHzepPXePZdYngpfrFovo3VjfBRsbmWnkSsPNqsjn3GOJIrWqAU5fB4OokboIcvL7pq/
wbGwpdXJhLBJHDUNYp7gpH2Fvjt96SO2YlwummBe9YQLoLMdMOLwbfnb8xk2knBan44O77RUWTmf
S6tUZB5qYxsr3pOkP9BvoCM90yEHXEoKfDeeDO/rzYrEF4cB0+xsfcnHIGog/3/pkf57GiH5LShC
7cZMJjqgXHPuOqboA8ELuzjJRQ1lmpS2akkKP0duiI2Eh+Sifes4355gnB3ByF+ypUol5Douuo82
LXDK/c8Dws9RnMp7dyoMXKuvWjlT5phGpVAA8EowLQqCkt3rboSMvGulh/FPGOhdWUACq/fSTHPP
abGmZ6bfDPDNeVjhwL24RU3iIqyaTPdXJIBV8KNQqbFcwp0TmkNCGC7NgS4b+864UjeSjfdvd6x4
hM8VqI4Ct5LQ4M2QTUM97dS4EWxL0MNnEHsMI7B9dB6D5E2xWvfuxpOTi4fWMO1a1PmoCsnpns8Z
a/8mpaBMVoARvvljyjXlXzKFe6KgCcBcwTRPnACfh761mu8E+yKh9vSyiFnRPpGu9m5R7rN//IUg
oBXLnveK4vEjPc+OkxV/iFvxeb/AoGuEMsPFL5M4gKx+tjK/UBirbagNV/w4KcaBbzNxar+70qcw
YwXJgNNuJJfpbS38erIgVeH2+NKXGOa9SHZqe7e0xsXslSUY7Wct9lFrPVhCdW0IOJfu5ZAnJvNu
lShUFz/K7z9Vqc9Ub6h/3dl3ayUk8gUPMzVPW9TNmpbdbO5FvBhSOwciz9A7deDYA2KowJQFb18O
VyFyTwXw/aG99vgK11/AIW2Ozf5xXtZDwsfTYxHsFn03p6l2M+a9JMVBaRdwFPjhCJsae2SEHhQz
u+U2p+HqgggXhLLCtKmgJSS66aLJWFd0nx7YLXcI73zprKvGkF7t0mNR3ccP04ZLwhd25TtEJRmZ
HX6OEz6DvRgKTPPhDZF39LGgO6qKLIzJlOlPa6I+YtRy7cNJQRg5gP4dn5U2lmxbOMiGjUeGIuHD
OWfsq159G9etZiAXVVCd6YGPZIGixW0mqiMnkJLLoXKNSkEd2mGdjJYZkL/spd87b42jfK1aBAm9
5LA8BM28BhAHdKFQno0Wq3JKxPYO0XN3ouWA1dZNdPQgy5hsSx5tb8phd5C1lzxMe5IwClIcoeAI
q5URTy7M1glBTJJSnmYQ27TbvCsWKU2/bPTgP8nBF6IN6koDKbOXp/WiLznD/bQIbGsj5dZvPc5+
vFd3ZWGgSwwPG8eIz6ILP+SRz72BEeZTFmbxbmiMQjSSWSsoNNPjdt2fYJ6rSc164F6bIXjnvEBR
lFy5tYo7IzecNMLLBTZDVwQw/ugYe0wpd5PiLSZe5QzEQ62EhX7GJ4XPLt7CS2HY0QATMmk/XQq3
nWzxXJRO6lZvNOjVs8vcPrpiRpsUpgt7fQUV4LkJUEhCsTWPoqB/QN25s9wMNE2J4jm0Z/EXF02O
dafxumQdtSdRWFzi2uIE6d4Q4ecGgMeVTK3xcxzQkStL66K8rr3W+yW373tVXA0k6BZa8TM9Kx+y
BId7XmbjYeJdyKryUCdIaUnsgUcI6H3q+7pZ5Flpj9qqOM3FYdCU7+YOjYNqa5Cy6jKHRh92PN+x
ttmYH3iiddkv2T7OfbRZGtMuIlE8TVLZhE+UMVLMkIzM4wPTMUhEU26Yyz6uh1P7YLLUAnClwYnn
O9Ag9/38hPXxt2HzcecMwPuUPgXMNE9jvjbSUOu5ZGREhgSRnNrKfzlTnL14fw93Te4uXRrJtwJ5
imiKwWa/Ka/b5qhs/B6+MiW4TwXfQPoux6Ql/j5VfXuXBg9scxTKG/wVmIyGNgmu4RfTCeC5pYco
q88FIdiCMWSUG6lxtUE414cCceRKT11gn/syzGdL/0HBvqAMIVT9RQKHgCdR1xEayueO5f8lqckz
4ftBs/ySA6G0wYxQaIOsHLupgiCYmG/QUDmZjNejrB5ljP2qoUpLqD3L/3uW+whYlb2KdJKdrlWK
qNOSwrCXdJONLtHjb7yGalhG/2eEgR6fvWi4huNX/1lJ5bPNGhZOwl7X7VETi49gt/ssGWLZmsk8
cc0BElDtDBWO5pyXNZ0vtiDjfoVkqF6CEOu7rbjxpvM9UFe6ThD88Y3ASdyk2S25xiJOoMq7yoOL
DYgQg9sNNpgMu0piSdglT3TbDiUhGOEuYNBXPPkcJ95RZ93pgr/8rID/bMwgheSQhSn1jQgPv3UR
7ogJWx7P9ZmfEy7Ddt8E/vpIcYsgKuPcnT/TL7ylYedoi3kTKXjGHo4BAaEq/HcPGmVZe2+bV1Ld
CGbquTmiZrUYhHyx9ETY0lInQCuONSAoIUbJUwBCY/lmrGraQfIXxqr4f3b5ZXNPeD3Qk8sldVJj
o2zkUqrhoePOI3QHNxdWDPelviz23iaqJ7H/HRKNZmuy7aKnnzah6PLZH+hrEFc1nm0SWnZMdZEG
uotFKY3oQpIK8GF6vAVjjSLrjMCBRc/iQg4ZbHZ5iTMDG7YrtkThEfB/maVFHxj0MC2SShcR+NAn
7HthwSkKhheuyDbYk8TwMVGq+GbIq9E516EniO/a4mfaRAVApFQSB4Hrm9y+fVz1o7bQNvHq2JMe
Sb4qjYYuzxeTj5zFQMQipVlgq2+M/yiKXxs4N5KUdv5ahLW/RGBuAtkZormztM4fI4xqog6QumTr
E6PyOe2Z4rMuuzCA0cm7UH7Ru2lq/bXjYP49rw8eHT5tKXLcpswiiAtG3BCK1NJiQiH2FCAC+FXJ
2RhlZh4z8sLSeYJv4ThroPPJxudlzD/mwA5pbiHXIDj1lVk2cNFCCBifHhhBhkXTTNjN+Ld84bIS
/FfXhNF3g4z5Ij6WCc+YhIqxX1ckvH/qIuaKPR+mjZRLRL2rfpAWj0zaJuZxaK4MyzBUwSl2cKJ5
7GET/0WmRIAV6LKl7do7x+FSuNUgQ6rPv81IeS0E8hL7Ih7ODg9/2k5KGHBIQKVJIPcBU6LfzaCF
U67mYo4wSnn9CAzo5S6LIRSZ1s/MXEGc8jYbc+O7r8kX7oKLaDn6L9u3c7zVvJYZ53i8KSfnj9qk
i8sBEPV8nwSPWBOlxs8MigpebGhOl1FIfXOi/Xrc6F0vKgWJh5X0fCNZG/DgJLRZHd7EtEeThnrW
RJZAOQIn9sIuQydPEZlWFre6VKIPCRW0acYSnm0HWiIXh2MKdh1Sne1LFHcqqlbk1G7gxzMaCBfH
Cq3iygTIix5f+PNe8kzstxWX9RfIe46yt5SCWj+QWIEDYrDLxNM0a/ymExyuIssBHojkbS7Oz8yB
Z0cBZkqLzprQxeAi9kAswFoBPt5hKrxqihG38s8a0p4Cr+tRS5udR8znKVtpYwcMqsnfJovoEHfE
+L2IEVsYigQiTOVAP4sN/4/6NqKPgv0Viw2gVNgdFVcqrWH7y7/XIOTYGKix5dBhnrSLLFLtwXu7
23KXMu9mvq7TRdoWiZi4JSNbCNHKgBf16b7BYtsV/qiByBrL6I3O4lAtkRO7LtQ/mmTLZPsfiDjb
FZiBUuZNqPuWiRAeKgmh7iqaxc4Krg+kbyLOvQEVY+BxU78H2yNFPgywCMVBZMGXjqXGvUwdhdbZ
I3BPBUtvvtHtrEI3P0SwH5sf3GeYhVc8q1MzUcL2mdnIBDz+ZTaX0QDTjOiMmwgTyGCCfUpkJKoN
SmWE80HQheXTNuKP2bc0cZVnu3RzBClabQV0P7cCd7TXr79x76r7pnsOkum3CHzOSn8w5waWQuWy
6xXhQW8X7B6ZkE4WNZ5p6SqKqH/brPSv47IlDdSMoNBh2duS36ndGf7kqiWn/JnDwZaoW16+P9wf
b8urE4ijSNQRzyPlCVjIfaWsCBixfoPtLIUzvrqhvuCh4EehY82K3p+4P1rcGXKO/g3qvrjo2r0X
ps5mNlljHShVd1EfNcqLpVvzN7oTpd2Jem/9iplFZVSTEwYlechqlgInPcRwmXBPm1/FZEw6fBZ4
1s4uiLD3zPqR3C1pEZwtQdT5qHudB6lA8eaeCYQrZH6lLU47ivSIIVkd8vVmhPVzsnbmdE2sF+pY
Wiwz721XCwH/czVYUzwBDCp89OsPamRy4KPFPd8Q1fhZm2UUssSa6CDhFvhnLkXBuExhU6dzc/0o
oXUSFZsn8l7hgiqJtRmE2MyOJ595GEYpv6Z8Z67/WdUeTMlZx+fEHxewTBSs33UsZzOlVdn0TWhH
+fCKkeCFc/xNqnvtpNi49Wo6CAL59ozPKWnNJl/Hbn4VcjI1l/OqsElsvzPfPVBi3wAPJZgQpOvb
S1vOZ+0Y2F7ziboZc2mkSAAGdKR0aSc7pFarHkayMvRhWha2WwffAPLDZM959AHYbPqxiqNbl5Pw
ZZBHQc55ZYgaOKXXlbHw+txW+H2sLHt0Hyv6c1Zu7Cb4SLUQMLVfgDE9ifOshkSgYCZgfg0ZjhSY
dBthRGJHDWHJEuhMyufKNgyvueU2PzQZWLMQYPBjGtRf/wgpXY80QYp2o5HY701u9XL1/+hJ31Q0
IHv6HxGTcBIOSm9QvN2sR/RhJAy6fj9ae4EyvU36SU/wWMOB3ZBfN+onjH8PdgiBK+UKhWBYjJNU
cUHrdO/FzDA/zsDpyb/Pi/lcziK/Ef4btT6jPfcmgA9ygiLdWStNXa/jByyS4lD7cP4G4NOVbVH1
+iDJKlEOSkq7DqGYg+1hUPOpgHO96Gl/ymEN+Dc9NPAFGIxL2QvCTDi16afr1nKBjVpB6yj/vgoc
anNonhRDbhaEh8WBXkLCdwwTkD3jOWcDfOjLyvvixX/dOnO1FfNgabLGHKZFqOKisMWv6Mk1N7K/
YgQvr3uINQ9dKZFX3jWEFWHoc5QUlRe/ufEh3ypvGr8W7yU4rMAPsyyk0Qv5vq6GXuZqHTEIMSej
9oXzXBDT+iTvA0/Zc4fwsdeE4xov49Ba52dPXR4pyqfyzi7Dad4V0kjGfvvec2SEuigPVI1ydGOv
pYj+sEm2NXEXPeAp1KxKvHHGlcfQYxSNGjvTE2O7Esej6Yuhu2fMeSyxgsi+xoV01g+X95BpD7/J
QJmnCKEL/yv2Wt4yBCuNyYsuv58rhlgRb95V63TOlfcqTFCLRHKYZL47MNfDIR6YLgtIsiUyJDbG
8+i/ulTL/wD4EF4fCFTGUKB+G4PCFAOiYGFgfzpkfHoSazsZKTwGWeu4zM5FJS4QKc2dyjs7Rv4f
OyY134HvFtlLv60xy5Pu7GPPRJ2eAlrQrkE8JXR8EfHFV7jmdVzRgT1SksRGOHtOsCLnmeH1wcrZ
QVzQid84/EaD8bDhncPusLZgRCfGIzjUGxxlZXH6j3UZbBSmnVPdqgh4Ezjw5mVExeiuK4jqLsSb
+nQaT6GTKeOISJuEiVvbTV/1aUiBRfpq15RJkT5Y/Pes12PBiRqIoCLXAnAaqSMq9IapslolLRzy
KHJQ/QcnlDdBbGhv0UFYdEB3DH+bmTmL7hFAC+E9MjRrKawR2Mm0Y/0RKTxxaquKBfmw9j8rhHP/
6VWZKMw/8hzLv2NDUrmHmvNLPIoU0N0mFrj0wbu3NDScSZFt8+t5UIaJcb5aoRwlPw/B8lNMhW3l
vBr9BhMwocoaei++FwqcMsheyCYH7ui1EZTtUxXQQ5Wls1ymiiprKlRNKCTZBcsrf5JWScTcbfah
LjmdVwwcuidPmsoGM6W4RBaCtbsfi+MHR6STt04yolHde103qewJGH4CiXQEWwVXJO49mp5l4Z+R
hweSJHkk18bF6NJ4Al4x8NrynnIKk+kxSq3FNM7JkPljTYek3VTgF2g0G8M1C0xd9wPBQY7Ug+rE
XIx4eAfPM3NvYGn4pY3w0TXFQ3//KRo/O4TFDKVBpYDwGlT6r2MvE3L9Iv82lf85Fd8MzxnKvMhH
JNA+LY3v0g9wcq2gxGwxLA7oK8OfKCO7UxZjfyUyVARlRhzNjBTBvcWW0QjvE66OtHw4q8JvZz99
4XT6YlmL6ZovYnxEiI6ZNApCrxfMuS0Zux1lkqFJRL/yhK+rMNvHpZM7yyJIw0K5YzXz5LFfUbBK
XkVdtM+HAQTlNcvViekOw8oshTp/JF8psGYRFMKL6hI1Vx6zmrb7xdhGn1hB5QYIwxDDSqsyJpqW
z2vwMSJo1gWmib6LO6k7RktR9kpSyebx9RVZHB3q+hRPOBVHDhJ7PQS1xUSlXR2L35Iq/KPcOtle
wWPSKvL/OnOwp1MugbaFYF+QvFP4Q6hLmBpKjrMMmCU5AqsHsfYmzH5RTt7Ogt5kckUqcIjniyUV
6OjvG71qJVFlyXftNw0xXCIjHF4/li5lQNPC4km4NbNyuxISFpfkfbaxxa5NwXK0slf9TXa/j5cv
BA/HbK5XL9E+fTLzJeTSWT83qvhDvwgHebSi+Zb3xRQoS9xnzD8glt4qJyS/HC8XW6n/PNLx6aGs
4doys8hIi6mlzZu7UWkjXM/0szQVZRQeDTQ0TWN3TQhbm+BUa0lch7oMa+AT2tKeyQGKTyX6VHiG
/TFDLmu63hhXjmWHqe7b22TkJt+xiSN0X9QcOexAmQDNke+LYtd+9XFwxuazXVdA56p64ic5R0YP
jRzR57hcRgGJY1WGu4S6rJFnbW5/sq3wgY9Nxc+P0vg+2fvYvw4eyBejVCMzECyyg/qhfkszumeS
8IcZIeujH8pCZay89Ms2QeBimvZHJST+Bd5OxUBQhU3u5w2H+B/jwgk9BKxar+7+7wfKgq3l/OwE
YFA1LQmoTEbZlnmpx3H8l3w6PFFoIgSL/CUB8i54v9p5UIEV3vI5JkHVGvqWCxCxC9NNSy25Ukas
CL/1dodOsnpnPkPsbu9D8mt1MpW1pM1PXlknEgPrGHOP2uHCktbXvgMyvEEgmgng7AZzMRcs4YVh
GApGMDieJ7inAObCOCXRV6Fwwk8WZUyk375EdyZA8CQ/uQnLtBnEkqn4DpWiTHZWCFEgX2naSK7+
NJ2QZobGVGHauMwgjphYFmz/QIn2gHXo1OiGGBOKxbQ7ZxCzU1f00vEVOc3uwELfchdXQ7D09kX+
QSUVedl/zTxvOPiokqQpQDRUOuWZ21t8ekQVUUJ49osX8OIAIxN3hytapFNhcGJnMV5JcPxwKrDh
KEqxrxgEKsO1W8Xf5qUmkfH0Td4xMPnVyHQdNRRzEV3xoMCe4F3x/YH4xPInjmQKR4kbGt4Sc4U8
eOSoVpiAGnJTtde0vPhqHP/q7NRGW3DTGqQfMyJNwhzL6FmCXgP9umHmQBCMML2xXkkC8R+arXZa
bBNnocMn7mZV40nDWT79pDnyF0MO0lIvn6fjj/3f4g0Wd2OY0CJd2dQxb1vshbdNifxLdmi7JsIr
RejeITkyz0i5rPWtS0YJKuf2Q+fphCw2zF1qPL7pJOWjVl7X/T4aLOC9wSfZ7PxnW8ATGpaKUDMi
Y+6eBJ4yJHaswcix82N+zswkfOPWi2xGyUPx06HLNzmHm4JX7+MguW5oOPcRGTDEAWZYrCapwIAb
A6l1zwltsIXnBNf3rVOkFH9aGUz7UiLhIKBzti5BGm9HmwU0nD4Lni/eIGGPJiaFJgbdV4YoHKSi
N8/QW0ub7DDV4J+Iy1Sc7EgK0LiA1yE22MCG1pXQFIEWX1r9fZCmMW4FoVqZ44bTvjebDgUI092j
vXKQ1ZTTAnIZcPiWszI1NROOZmTtASvobJJ7+pwIJZ4nCFRNyO2xOOFDk9Tfx+il2Yhbn+AJolVk
1p9uCcfdM0rompsyVm7t+JhB2ZBypcSlqyvXw+0gX2A7z+H9kN5GQsfdPLY9V/FX27mBC/SUzWit
N6r573lgB2DmPRItVcY2fNcsV/E7f4grKNMBaDE2hhFVw/90VXeRxzCY9VszXCR6sSdA0zjV4nYv
6JnK54jQcqLZ8+a38htgenAFGtjzlCRZVxUPJR5eletvMt7Olft52UT/64UqYRSaCbSpjc81JP0i
FedhTZ1TFQI9Wutg38Pw92X8VAHYnpstKPU/EcGVlhOiL8Dx+j8kHXVEIDuoZX+2MiFS3h+A+Q+0
aHJJOAMxSHwZGQQbWoGf6hKMhYb6GB7+iy1DSEKkERy8PIfxWJf2x/VXAZb7uVRku4qfXdzg4y0f
dhJbewe0k/yu57+FnHGDCguDz2hNgxY83i8+7uxzyMPVKYFUC3BEtxftVOJHQEx6JVkcCeCtj3/G
c0tW9VB7ub7hBrcbtIVZ99l6JUHApP18DrikE7AYA6h6/7FQMP+d0cY6YgWxZQtK6nF2gBpHxA5B
TW0/Mlm9RvR3USYB3BI+BG+mxQab3EyaxwFLjmy2gfe2vdtw9PKBbPH+qKORCUYe9zc7P2HSdxse
uEldC35Uc8U0y9Ul2L5XdQOIpGd8uNN96dXS49AVVxo85JPIcMJHg3N+bSdWYa/yY6xaYytBhx0H
RLiCJonZ0NiwzZa90TDqCGwQUPbxEMQNcr/ivG2hqQZSia40ANPpwtsFBTW2Y5yzS9c/nXz+Gh6t
jyQ2RRjahnn95ZSdPB5We3G6mjddDyZD/G3Iif7WqanqIlwI7LNlqaW5Z+PQ8tXezc+JmKBL0n+U
84qlIULuerPYWXlvRVzx7ClfnbvsH4/Zsa9AgHX9s3+mjeoOUmfHWnZ8VVFCNuIhXCl+/dCwx95+
YIMgy6cNyC3UWKL8OopjnI6rts1LRZiuhLjqGCAJ4Tj+/zEXgVCBT4Wp30xbfTdhmQfBhNn+ENwW
I1HtE4nAbBGGtxwWsZqL9CiYOl6SXdeSHXRX14nuqnbWw9ryuaVAEF5p43H1JYVfIto/KgL5BdbP
ENChew1/0Y0b1g154gCbhbqTjOYj51iisEIsvWnu5MmW8kvOGT8xfATvy8QJBIH84zN0XUXGbEVS
B7jRjtZ1TXnQlzJKt4f83Lq7RDELGo5Xs2GuQxSB9S0pm/vpBX2BmfvQoa4vWUwOZDPNwia1c+eE
3Rxzy3xX9+bOeB1YTfzSrjpP89f7g24EBbom7QRJ4AldtDzVjqZMiGHXYFt5iqMQ/qr3dnFKH6MI
VuJhwJsrOFqdxaG9mCgkejErPjy1Aaxs1YF/pfTHGhDZBI5tSPihgEISqxnz5IbNSzzdwAxHQvme
t3pppr++pL32sBHPisHeQL51iFeJqAhyPHeHQuTF6B9VAY6KQBKmSkJE+Ukln7VH04BMj+c23NTR
SIionldlpUoFrf92OtV8nikynib5LR5XfnWDzSAdyXrvZYjZa5ioTL+7eudaUCMmVBqj/T1L0LZh
kX23A5bgBPg9YYf34O8bGnBi0eHfkgxvrumOwwhzqutEf7lWK5xkYcFljQT7TLqBlHf2qKWtRb6N
romGAAhicvgc9VVCNkuNor6zDRiUVFFvszWmTsjXG5JHX3DYfaRqlGs6EumwldouN7YeSAzW/ro5
y+R0uynJS0dfUPCOi7vNlJDDBqSZ+gLbZRpLl0psyWWTAgvT3e4KMCkblhEVrPDKrqjujYDrg5/2
CuTCsXId7l0KpPS1pvuPpHwPNjm5PnykBcsAuE7una+U3GOeFeW5eBHcJTDFCaDoUy+3ACUYzRT3
8IRCruWUPbg1jm+aM0xZ/lQw1wZFyMyYwd8U+UWJKXGo0huEdafWkPN31O/4xF5T6rm0+vdCB4gF
tERgaFJf71b6OkxD/Ac1pt9YkB/hE8NFAnp2pOCQn2gO59GgCbE7kc6OIooQ6jSIP4IdCBzSgRH/
cwohmHBF//KUKARaxwV7QmCLffUFoyfLAUJo27ZZmP7p/NAQcsa187Mbaz9g9FudwbvVVkTnHOmp
jVtSjRZh50YhZdFxHWOZZXHv2CPqWF7kLjXZIkfT+3UEKrHrEDWFBU0all/pjFo436QU3UIVZMdu
38jxphXl/92YzKRTVTGPHn86C+StNJfp575OTd5PM67aBkXChwTujFWjz+kG3wmnqqosaJPS5vjR
3VZ68Q9SzM5JOdMOBfI18oIV4jkRUg/SSpKLWohd7cem9B5QoCRraifBSYMCVCmwowvGHTSIjYDL
hcWGWRqNZxJyX1iiRHHHxFfKtQk4x2PNpkbB2E6VM8Jry2X47F4YnClcLgCNt5UNEU+1L8LGVEKd
CWPUpeuE5vYqvq/9IpN8j1FvqYvsOJvgwskUoPJxCyo1MULxlmjklDgZvO9Ev8+P9XHZ7Gx8sdzc
g/aCHBCla00rceNS1Y9mMYVAund5pU+5IzHZFBvqUWHpXFNFsvco8dngGapQrRyH4QXe6SYnHqzL
+w6y0Ve4oew2QaF2x+oSqGZ/vCjZfabhBTI5N63yH4EUlpvB99gFrX6OV1rtNQ//WFKqFtKYfrov
nyTkAw79ym0K8EeORNywXQ/vh+EJYSAJq9qSegSg0FAvQCuCMl2+ZFeYX70VreK4LdYVyZzAQIqG
v5bp+8zg1BtTJWNW/U5aW6aYhsRaO/wAJWlZyIaXM5qLGscenPlApcBjhtIreaQQuoVjtgHd2XOV
zisvvy/OHpVnzTNmqQByYTMLtuJUpFhTN2oyI32kjHLMdn8ws/qqHHNJNqd5DplWgVDGQW+pMj4C
gEENcbr2E1EwPLHG9IKnD1gqK/T5f/jgyXhYopeQ4uRwGPG86oddWmzG2m2IBb2DnsVM4RF3fIbd
25pZDoamWmRyMOogG+xHjYhfAiGoTJJOAAYw53GKXetUxTi5xhLYAVVJulLQ/900YrclEgfBPhjt
kvNlwqnOUlznBFrMMyEd9OsZ13x30NJiCyXntbuG1HlG3D/5Bl/FC7cYUZ92G3WCypJewhS0M3Un
J6SCYI2kGRZzm2oucGPKpJUu4SBC4PBNgQAmwtimYmzJUqm4UORfyojthaCIF6AtOWUSxrdpxip0
sJ9aCiT59nMju7m7WoyOpAz49/EAyaBIievE1KOM8DiIdFD3tJfb0ZoByAw82F3HnV85WpwPDCZz
tuMuS691HYZbJhtF+rqfW0atQOkEnJNWZm18BMWkHSfirOmCw4Ohmy4qkkvBy1bdraCUV0DJse5b
Fvak8iHHpr7P5j9UK8rOjk9HFc6UbivtbDhOkzQfLP5TKOqA6MQVNLhM96NoHI8mO4DyAJt7AS2e
UFRG0rWEvybqvEwG0LkQvVYfHUCrLZW9clMl9j+JQtwWq5pkU8BAj65VIi/EnSojzHnXs1FNpm0E
M/7nU6g4J9bTpx09OUHG1m6t/hZFcKRMgNSnMT1ICCPXEJsf9sU=
`pragma protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO��� ��:I���^�o#�s�G���Q���p|����}��w�!LJl�J�+�t�}ac��6�"wj����+/^�6�T �:ɺܑ�SR�[$�EY���e�1go���P� �`[z���sI`>AT5�WF��\{��R� �~�xLƂ�\b��Y�oK)��ץ$��Ё��2#��Vp���[B~���T!KՓ��D��� ��b�>�A�{{Q�5�2���W���^����y׻���8��3�Cx�e��٬�I���,! �y!�Wm��^�8�9�z�.Nu^�b:�ͺ^���FqmV���PX�G^��٧�&MD`Ry�-�qK\YQ�6_t�L|��9��������ֳ����"w���e)ag���p'E���Z�jL���>����w8�O��:r����=��Ia�5 ��4ơn�0I�����/P�6l���B/*��� b�`M����3]"�B�*�\���b~ʸB4�gکw=�n/�J���1�@X!�l4d�)�L;�D�%��p����έB ���
]�z��u$�fCĞ���������]<���zM��4����� �^,�ADd��<�T$f������'�M}Lu��� ��~=`��?�[��W�y!K����k݉2��	_������WpmԂ�@��1Ka�X$x�m���M��Llg$�i�ZĜ,�t��$�J(h��	h��`z�i��?��MV_����"�S��4�U�3�$���Q�T$����k�����So�"�ա�W$�x�R<E���q	�K�';~�g���W�����rN ��^bÈ��y���/����'�C{f���>Ѵ+Ǐ�R�l#k��V��ػT�"��yd��i��
�g�fr���б N��������o���M������p��q�*���ϰ=DW���Nl�$-����TN���r&�?����ひ�X����x�*�v���H��zQs��	�����,���I���k�K�W���^m�7I�;Z��9ң)ʹ4c!:F��+Dwt��Qs"�B�D�>"T��,ߊ�@��y�m��$����1m�bt�gUpM�:GO|o��Ǘ������p3�J�U��r�]i�R��.ض�z��tU��*�?��k���U��3�i�^Q틘�AN��}�
����K���F2��|�9�"?�P�e�-/V�P �ƣ5�W'I#�a�a�-^��r��ǣ�v�A�	\��}=̓�3���@�l���HY��X�l��7J�20�����F^n�Xp:�cH^�Ƚ+p�Y>�r�y�k��o=�u�QY.dTj�1jw�hx�7�@�B�l�iQhhY����d�q��_ dY����L�ם�m`��Á��.���i������Vk2/��Ko�m_�"m�M���S�.���ME�
s��4�.b�#��o�ඨ�����: ��D���'���7�&:mN^Q��_`��2��M�_���d*G�ʴrHk0ՍtIKxN
5�%� �FH�(̤I�c�[�o/��΢S5xxd��ģ����p8pA\��~L	��]�q#N��_�m�'��ѦY��P M�J# *�[�o���z�"�!�Z��Y�#���I����"��"{�|�(x�~6E��1-3�������Z���V4.�2���*@,�F����|�,!nҔ��F�3tG#���-&X�Z�y=���ܖ�_��$�$�.�M��5�#ͭ�U�T�{ZVgb�?[
o'�eH��Y�9�����g�&�Xn��{4H/ ��%rr�`q��5ދ��4H�4|��̜MJ�}��Q��Y�S���[� �s��/�Wץ���o�Q����_�����B�������
����5�?���K����CA�W�����=x������
{Q2f���5�ɱ��gI��ُ"�eŦ�,�辳�?�~c>�E��6T�}�V\aK27Lg"��0��@x:ey}�鉦�#��Q��c��
;��ۙ�ؘk��6�t;�h9�M)�P����:+;?���/7�Ϣ��R!�g��sRT�&���P)M!j׿`�9����ؠ���w&8#�.P_!v	} r����E�����2�g;����A~��CT�;]��)�4*$�����_��]��rV�רZ����v|������x�a��[sw�ۧn�8��A�D��#�����aI�Hn�b��6�u)˺��IOúp|�a�w,)-�IԢEd�m3 ��V���8K��� o�T�l�Z'B�̮��O9��7y|e��0�K����M�苮 ��"��6�4��w�AP��y�������016�]_A (.�2b��.X��Tc��ڴ���xC��LI�L��$>�,zd���9؅����
��'���Y�:1��p�
��ʘs�����gm����G>��_�V�W��A�c�T��<�YG(A��
�T�]���Y����3]��J��tn$�5?����
vݧ>KkI��N���כa:������&�,PUS�L۽ȘW%�m�g�v�����/�#��;4	?ә����F��]�� f�^L�[EGl:�?}Ml���w��e�Sj@u:�RzHQ<@g%KT�YKpX\8.�"����lp<	_�u^��9ʨ%�=���$�@iIJ��c �����,:���#�Va�sП�-�4��~���7�p��`�~�������TҪ�z$�jɪIH%�������o�~C�� ،vph��i$�{J8�������ʻ�
;��!j�O� ϧ���U	O�F��_(S��n *_��_`iJ�3b|E�ؙN������M����xh-�m���sH�_F�c�>�Dd_%���'�	k՟��\ �Tf�	*��}��"��|�̸�+KF\-�d�.��γ�.������ 7"�u��j�bD}͊�5@q��� ��ّ#�:	�6J*8\N}
>~�-�dCOmA7��I<M���uEُ��њ��W�'���"�FK����&�d&����}�^��'�=b�Ӈ,����&���%�-����+/�:�|�	���<Zڷ����GH�ȯ����u��R.�#~���t�HȥDe�G�<�VRr ���c�ѵu�$�1����M��E�.b)Q���Ș�5X"O�aT�4��,��tu����$f�X�lo��jңF�{iC#���T$��&�<��6�
�t���Z�ڞa��|�*<h��ʸ��X�P��DN9��� ��3uҫ��^s�"��P���w"����h�d�����Fn�,GgHTR�a�Q��&@����"#Um*D��P*!�<Y�㤬yH!\��	��mO	E��\����k��Ϸ(�	�s��X3�YB��\�6�F����U� (Ȯl���T2­�}(�H�j���$(�TA0ۛ��>�t7�,���d������)��	=� ׬��H^���r4P^;��y���&0�bjp]�k0�B�����d�G�����D�1@,�5N�k�C$8t���mH)p�Ah�n�5vs������/�O6iKR���Y�R���V���҈/�@�"��	\�e(�̤�5Ӥ9s�^�T<�o�4��������"r�.�N+���^�t߱��iwF��q�%p�5g�
��$��s�P��?�j�0NR`�oɮ�HQ�p9�o��u���bnk��:�a�4Y��O�*�iݚ��m�s�Z9���u�/����G �!5�漢�m=Kyy�7����M�y�����Bڄ��j��xr�ԙ���gZ�G(a	#���������e"7�$�sC�j�O�n=�FT&�F!x���%�����gi����}%+T�h��&f_�Y\3sï� FL{F�W�D�<܌Hye�����c�1�u��iZF2	�Q|o���_)s f 4���%�(ϫ��� ���T9b��N�iV�����r'@}5��Cp�s�i������z��8ͯ}"B^��E�;�з�OL��r�M����c�'�}���%���"��[5ıN���߉��=�l�x�䚡�fz�����O6et�h�ߪu$�u�1S�4��E�Z�����,���"�v�5e���ʺ���;���=��P9�"9d1)��l�AU�o5��}4Hk��aG�g-�`�c���/>���0���;Zl����a�)���sL��� �g��p�I�f�%�$�(��E����~�<ֻ���0u��*N�(�ɼ;���٦��ō��FR��}��%���Z9��S�t�s?vi�Y
AG���RnB��5e���1[��~m~�����-=Sɵ�K�"�uU]��+���L�E�9���`������w��y���kd�m����.}OΆ ����6Si���K�����~[A+�!MI�*�q1l,��[x�7�����s�zB��*���Y�{�\ i�y�a�F��V%�H{�ٴ���`��w;զ�чA�����øM��Z�H�m/f_T��`ˀ�H��)��YQt�s�-H��;.LxO�tS���D+ס�16U-f�>Wx>��,�J�3L"��ўC�Y�!3^���=�7�i�9�X�����%<A��d�%b) �@�$�.M�{'��wn%��8j؝����`�F��#P̥&���-�L4����&�v��_&�ݘ��'���ڙ��M��(��N>��+[
=�a�F�<�[�Ky}N��b��α,���G�a`Ic"Q|� �n7��[������jj=a�Z��Z�xZ��~��%�x�*������I������ p
ED�K�	1=���jh�&Y\���!�~+�a ����{���� є�HN1"lg)��"��"!F�%�YG�&�����7&�p7��`�K5S>_�k8������D��L���*���7J3B�vf(b}q��%&)E~{̬�#XA�m\�1C*�V��7?q)�__��BS0�7�(Vd�{kUp6_�ٯ��0�Ĥ25�n�����Ԥ(���<��8�c�he�qԲ3� �7����[T]� �����o}oGk�i�7��B逼�/�	R��5�[QdU%�X�����q�z�0�dL�������6�w��ዿ���ճ��fZ�T�ՈX���p^� ���Q�����Kۏ/9�PAzi�ob5E�`��Z�r�
�e���[���x���t����������x��u��m~1f ������Q�Bc�R.c�4LLn�5Ο�ī��VWR�+�,5��b��>�����4�6{�z��tU��O�l��ޙ+�e���W	�V�%�Γ	�7���pD���x��O0S�z7�K��*:��������}�}r��_x�5d�p r���n��A)��/7}��77���sq$�	g�-�ItFw�tp$x�|5�\�ꞽ܉�����Vx�Ig�[�ک�����"f;a�e��y�!TA���hǑ���4Q�����b����U�����n��@�em��t?}YqJ���i����m+ϯ��e��n��\{<�yQ���"�\�v'����<��9:p�0��� �ͅ�����W�����p���_:�M����t���Ý���6C]x��(�l5�J�`��e I�@PX!��Vù����$���8H`�B�p΄Wu#�$��zJ.|��W��{Y�R�2#���߭�T���va8̏�a@�p�:���bR�1!&� �reN��=_~�Ǩ��e-�ɕ��y�wF_,ִ.�	��U+�_u���r�	�R�rU��h��W���E��ξb>�6���$�&�>?�(�����c�&B�%5��{z�ڶ	�:]�3�z[�a����?l����<cDG[-��t���[�	D	F��÷=K~��Z�#��}?���=/s�P.���5=b6yb�:i{����TmHi'툋�R�$L9\w0E+����.��|�)[$�����i�+,}����,�,x�Nc$�U� / ��0�Ln��= �1�Jk/e%G09m=ě8MS�7d�;��^wm�6��s�	w��Dn�
�qS����tTl�a���癱����r������EVR����(m"��T�����o�h�(3h�������@��/���Ƥ}j�#�Q��%Lȹ�$�\�'o���0X�������5�H�}���V�7>c�]�y>*f1�ѫ�;�^�{���w�@>H�U��٦���6#,e���LDȶmF�fˬ���af��B!	�PD�z8����U�J�T�ʴ�l�+NO���n�-�
?O6<���Z�qF4[yFb ���S*;���
E��C�6�bͫ�=�˵߸,��$���Kjyި�N下�T�{2�� n U�-�����H<�]:qt� N�ַ�
-�h�:���e�ںє�=��>�\�;\%	#bA��&��#bB��\�,c�mU�=a�r���ʌ$dQ�V!M߀֤1��}���ʙ��#s��3@R�!�jQmi�R��S���Y��,X 02U �"��#?ȯZ'������}&�"BEqx["C�0����RY�^�NP?�U�9�*�܁���a�X3#�D	(>��pc�<3TG���J�K���[؛��#�|��]��T��R�Ϭ�K��~4�/��2����{��aB@i:6?CQ�4�׷����3`��7;�c���я��2�V�燦\Z{ޑU��Ʊ�_�c7M�&W��4�0��X<��R@�%.H��]/�u}z�7b���I|���?wlw,��.
�	X0��r>�1���(	�7N%̯�^10�q�S��m��hJ��&O7J�T�����}�~{�#�8� ���x��k�q����a����v��9�sp��O�Vb��7��D$sV��{낪��`�^�C���=|�خ�/�%p�g��|��%]�'�#Nc�����^�~��A��'7_@M��ֵ6��yF�y���2�z�|�)ǒ��cC[e�_�R�"�{�u�ݥ��S��)ٕN���:A>����[��Љ����Gy�⌰�݆�֛�j�ᐌ��[ɼ��q-Y�$��r�2�����X��%�ugP�,�x����)�x�"�ܐzb�!�HE���νG�c��}P>A)��H�,��R~��y��M�i��CG֚9F_s݆���;�*����y+S,��e�d&(3L��l"��^�h�͒(v�b'��
�0��C�Q��9�t5��S���3���(�IP_.y3�]����d�b����x��o<a�Q�N�2��F~$2E����hGM�����9��+r qF/�A�����+4�f=�x��œ���t��;S0{nB�Om�JY��آۡ43C-ۚ��^�Ԡ�]�x�Xh��/�%d_�����A�N�y������xĜ�2i�oQv�'��Ȃ$��}�[�R<:l��.��~(M��J�8r��r�7N�ᖄ�+�� R2Ț�e��8T�iVF��Ο<l���݀�eFIBw 8�Vn�چG�ٟ��-7��;s����	o��>:��,���N�]�\�����[ON���2�2��'3�j�0�"����3A���'�$�\�}�IM�Ihiq�1s���Kߕ�1+N��H�P�c�x��tH}c���L1�7�Op|�y�1�U�0����M�5aaf������Ƀ�㗶��@�o-9�C����ܽ������X�:����7L��3M�;�md����&�ш2��z�'��sn}'�,�\[����>��}�I��}]<��ã����ϗ��Aċ���/s�O��45�E
�i���R<`�L\�����p�,�r�
K��1�M�sFl�W����&-�u��_=���f�R57������O� #5=�����D�����@1�S�|.|�:��xL�d�an�r�Hyc��,v!�Z	����B0��/r1�-ܶ��P�b"�G���!q(qqs��V��c	_�Cի�l����� �s��>ө>�I�ɗŖۀ"���J�Gg�Hf��M��*����oLO܆�|���ʐ��V��l �F�ˋb�"�*Ta4�I;���#.�tcN����;�H�1�,NR�5A`e���q�M������dRX�	1��\ׄ'�c�j-?1��(WK�� ��hbGom�ey߬�*�vp�t�r���P\���S���K�v���m]	�~�\������cM
O���-7���p�5�{�)*Ý�����x!�K;M����aCN2�^�a\tv?�z�Se��Ʀ��c>��1�^�+��tԴ~����>C^�����?l^Ȟߦg>l��\$��:�q�Ԓ��,β{w/7#2�]�k�"�c��Y[������9�5�0G�_��'-��f��"�QŰ&ڶ����@�M�J�Of�?'0��dpf1�n�
�y�D$� -���5��Hz^�Ȧ�.��{��{��m�����VN�߉U~�b&$�*u"�'㫈>؀��2���k�� 眜Z�D:Z���	��u4@�`a�ܼ�WS���	�@�����g���$��`Q�v&l����h ���� r����0�DH�iA���<�d�/y}��	��� �q�6Q�YC�?�����K=�_��'�gc[�wVB�
Gr@�z�{l��U&�ܐZ21Q��3����c%�ѥ�{)���v�/��%j��4��R��mv����2�h�,�om��e�g��NB���#I3�)��p���?��F�]u�<F����/�_'�Ԋ7,�F����
pu����N=�Dd���׾�H�I�Vb�/�Of^��DHÈ��v(m���q���0%<������=VHs�o�_}Sl�����P�������V���ڝ�e���`�[�)=��,�o����ڞ+w'b�϶��$�2ȑ����%n�b�di�A�t���r��dé��7Ƭw�2�J��`�Y;�5���u����� �A//��k�����1�]�<��_}	�tLy�؂F;���)����3��13��@_>���$8*����A
�/2{�}�w0�9#��L�pmj��݌�8��\��ۿB�zU-Jl�=�x��Z��~S�(��@�^Z���>����	��f�ǋne�d| �:�-�z6��w���+��嗸'��^j�����;f�۲.��3l�qV�_Sz�`���h����߉&��_0ݯ>q�~�"��χ��"�����٠<��K'�ŋl�%��t M�����HSs43X��&�,���L�G���F<��J�H1����t���9��w!T+�*�W��E2������7��Vj��>���%��K��)e��T3߸jy;J�K>��yz��V�	g����g�AL�)W��^�d�i@1���6�9@&H�F�(T�`�_��8����B��8�k|x���>��FE�;�,�������j	a=��[�7�md��gߢ�Wǣlԙ~彘��e��������(2E���6��8ԇJS@��>���
DaJ�w�H�����kS�Ӯk���~�]NBh0�?:���$�Y��!��w\�%W�DEN����s������w���Z��on"u�_�����!�-L�h^�kw(0��	<���'`L��X�V��I�����<��0��!�8�ܸY\Ȅ	;�+b𫚋�
�ޚI(���tա��	�3_������2+�s�{��1�9��q� �{>klW�ګ�jKh>��e	� �E�G`����o�+zK�*+�!�?!��j�E� C�������Z�^^s]CQ��i���T35�<P��E��Sc�"n�i�!/�x�/F��m�N:Ƨ�;���<SR�G��N�(�)Ů����1.맕d�D
�]����
�����|�T�_L}�(�,+����1��w0�}q�4��cwV�;�Eގ�m�Ȧ�:�7��O�νO󶑵)�xx[��>�|v�i��XD�G�A�w`Y��B�s#i̱f����H�n�ZY�s�vke�W�(�
��֑����n��ڍ7�E1�d�&�&e4>��H憎OG4��>v���>�$W�IM|$M��!Jr���\x�_B��*��>���c;$3�l �7g�a�q�:'�׹��.[�5CX�b0�9����	(��V��������D�����yQ�瞶�~��ci�'�BA���D���7jD�ch��Q�1�Pޢ^Q��t*��OQzg�f�r Kk#��DDM\J�c�]����c#��Oہ�c6�t���\�Q"#|�,�ug��}2«{�ρ/����u�e~
�A�w��y�dҫ�f7�D![%Hy�6P��86�<�"���� ���d�(cm��(Mo�F�m�0�}�.'UjLe��i�ɏ����
7r��mfBVEׁU8/$ax��V��K������L{���Z�3R�ώ���l�Er:목��� �SǙ�4Yӯu^���Z��+�m���5�Z�K��*��G�0���e~��i��. a��<|��!7(��%���W�(�M�9M���a�����R�P?gC�]��X�ڠJ��6���	2cҘ��^����:%�#MR��(WgEBָ� ���3ۭ�jp�� ƥE5f� ��SxM$���7�^���gR5N����_�8�-pۉh��i�N��7!܈�?&em���M�����k/y�E&�T5�;R�GC*U�Arl	�}�V*@�����Z�+A*Ů@q�(l�<$�
������[��vFV9�}d˓�,���	!$SD'��I^[Û��*r!��V�ky��;�5�"��U�d�S4�W�����[ɜ��`&�c^�H���P^�H8�o�8���T{���������>���ft��9���s��qH�s3w�L*5�#��m{����;��j��V��zM�]'�I��8ks�rdy/�P��E�=��T+���Y/������%���c�j6�%îv�~���#n�ר�J߸�"�;n,m�>����;z��#�G�˄��|��c�*�P!q�ǲtU����ab��H�:=A���lf5�SЀ7��n�%��/`F&U8 ;a����`��R�10�4z�NI��0��t�䒘��8"x�>gn�=������OE�]7"�h��tu(��Kx`��b�O��,A�RH�x^�����7?R|�M��R���t B{̯��l�Q��Ȼ ܿk�9���s����������Ѩ\NK#r{�!S�����9X�1ܘ=�kyuC�d�NA.��^�w��Gܳr;����|�a�er��B<�ymy�nD�B:��p{��q���	��J�y:	0X8���!��As�~�ѫ�����1H����i{�F�<Ǩr�9uK��^y�y�v��kkn!F*�i-����fz�s��������G} ?�����?f�<�[|C���KS����s����y��C��{n�un��	��� \�KG��1۬�xǴ2R�v�B�(�M ����=̟-蟉��L�cJ~lɔ��9E�Kek����KK+��C�G�J1Vt�2,��Mh|\n/���<����2�P�1b[�W\��</+[/fϡM[�Z�h�6i�!��:��	�F/E��r���gl��W.��sU�:9��H,�,6�g��Š_G7�PD���Z��]2�g�Q�a)�j�tO���9L�H7c�����<񪴯�MR��Ij��cj0[����oA��.�_�r�NU�g�X���ZZ��q{+u�?����]��Dx�uB{���~��C�#4y�Alyl�?����ѳ����_S���������
~%�'��O�e�@t��<"��#ĚM�����������;���O�� \>��L�}��=4�?�^�Cs�Zj��hc^��vU��Y����&�{�'�o�_��`�!��Bs �z&�}�w��@|Er?��aeg���厉�h�d�M��G�Ջ�(�7�X,%EK�͖�V��1���x����RیG��0�z�GO�'@�S�
�dk�jSZ�k��۝[���ݗ��^i	�f��Sc9��Z�Y�Ai�ܣ�X]�����иS�o����:Ȋ���j�eĵ���Z�;��5��4��{ϛ�c�u%��~ ��Jxz�\�b�+�yc��L.%�k6V �R_͐&��=]4^�EC�]����qʄ��#���	L��������y��>�� ���u��;C��$
����϶�7�P�k��O!S:�������p�|���÷�����"ͷ�1�|��O6R�F6�b ō���/��]6��\o�/)�����M��N�T��|�eZ��[�;2�ݶX_�E�9�@�X�C!��Yt��%�]%Y�6g�seab=�^�C"��F�B�KE$gfMO?-�1�j>����)�l�Ӄ�4%T�njhXz�H 9w�6�dCG)8V��wH���8��#L�P��x�a��z[��d,=�w-*�k�mk����Lx��X����y�qx�ʏ8�~�w��XȨ�Q���m�}��K�ٔ�&4NP�$òcf�Sk�4��OxY-����(Qr�@]a�0��q�
��@A�n܇�䈑B��f����hB?�� Y#e�}W�4i$�	E�=���Z6+O��6�d��7��^�^0�I��з�����b��-�5�d�������QU��L�ԾY�TJ2:��P�4�b�����	��6���,[[M_����8�ğ���6;@��Q�_L��.�3	c��m/��(V��0:�ri�7t>��d��<���u.۴-O�S�9C���!�FlY�W�"D?���*���ά-�{C���Қԯ���;�U��[1�4�-̞�(O�D�L��3���I>5���DIPܘ����������.�n��� �
�i��+��{�o��c#���n�vUv��Ֆ�N~1 h,��ſE��?�vUy6*��8���S=���2L��f������X���8����-�z�5�9����Bܛ�:c����Jb��W��.��:�^1V����0{<i��P![����������5^h��uW?s����؟TIPx���URݻZ���e.Ei]z�-/o��8�
��,���=`���[�+HmƧ�c_ۂB��~��>x!�C�z6P�t�b�R��rd,jϡ�	K�5*n�'���".�?Ѭa��l��8�[�O����q��G��/fa��5I鹃5�����A���<�'0��j�,��� 3x@���9�O�$Nia�E]o^ �D���<���m�@�?�=s_��ʈ��u�|rx���$��+�ң�푗�T���Hk�R��%�m�HS "��^����S�L|���p��A\�$�ɐ?���|��T`�� [1>ܭ�)���F��Rت��ށ)��	�����Ac�veJ2c0gJE�"D�ź&����A'��H���b�PWg�[�ǧ���0m0�H"�3��	o|ro����Җ��gR�𲒙���� \W/벮�>z�ywg�����u��aGu��*�~GBuf�u�a9e�݂����Ȥ7D��#�vw��v�BY����nC��:E�ʮ�D�Ϸ��L�w %Q�%{ޏ1eD�8�#N��c܄�!d�*N%�&7V�����r[xD��$���S�����l��8xǌ7L
A��Kc H�A�|�,qw)�L~�Tr��~ErY�-Yˊ�&x�; }.�TlG�CQ����J� 8��}x_�|�MK*8)��[�:Uxڋ�9�O�����M�^�L��-����Mn<�=4�u�haP<mû)@�P��Ѥg�{�V폙)�?�m{MU��$.�Y�7�dy%;^?��3�#q<����P\�74S˶�������g'�f�xP��8=���!�Nx_�fF�	G@C4��܇��o��R�����Q��O�<;��f _SR� �Y�Qd��`�,��T�O$�@�Ɋ���Xf,j�$�p���"1�:�dbݮ]��,Jσ�nD�ka�6q�s�8�!CQ�;�Z
拡OJ�f����ls3;<Y����o�v~|ܹA�����eb���	P�H?6R�h�'�m&mP��Bຨٻ��:Y��v�(�����L*���/���
QY��bs������Z��� �5��!�iv��c�t+�7�8W_��Y�#�l����EHc� ��1Xp�M�s�h�����ڑ�Nx6ܸH�x�8��6��b��U�q�&�G�D��2Γ<��+"*�o���2�����=c�#�v[��٪w�U�@��n�E'�UpA���멸�q���#��˝��В�s:E*��OA�ȴ��u���\�(G��:��0���-�����@��s�Z?����7Ix�*���1��j/!�
�{��T��;싑�u��Q���P���1S���x��E�
��A���([1!�b���{:�?�\�ϸC���/z4-;N�Ƨ�NE�i�%��S�qX��x�]��6|�C�[���)4E�����)��8�i K���H����z��4����A�l�0o*t��t�3F�z҉�p�z�jʤ�/>�Tݵ�K3�!Azv�!��]6�b��?����w�W��#MK>Mi�7���7dՅd���F �1A��|G����/���7��ư��]�R���T�nR��Y��m6r�[����ES�e�������#�d�W̬�to�EYكdo!�t�aw��m�c�i�M�7X�,�:.���3ZA����u�v����0A�w���3�6�����\���g�����w Bjx�X��HLTZ|�����k�[�BP�V.~%�q��S��V�=���E]M1`�x����(����y��z9|���Ҳ)�|���eZBc ��RW�HD���}itXN���<(��R��� �1����tb��3���S;X@KQ���Lm���}
A,��8}L-!z�
;���[�!��@i.k�"|�M�~�0�?%�W�9�,t��C'� �������CV�|��4%�+w�� ��J�C��%Ը��w�LM��y�lҫF�oQ��_���\���(p$4s�FQ ̮D?B�v�����u���Q���|%Y�]� �[��RyÆ[4U������1ШW�%�1Y0b�J�(�"./g�de�ݖpNOj��.�pI$��g����s��nD@���LQ���J��SP),Ì�vv�����n�u��U9��&� �0�P�P�CH ��NG ���Ii?MUKp~�os�2���'�7)BH�S��w���
�.Hs�:�`�`���(tX��8��|��=g�ޝ��T�7����� s���� < �y'����.�ր>�����8Z���b��+������n�E��#����>hlP��o��g�����A�yV�]�h0�x�L �!�� 3L|,F \��Ti�b9ߐw
�CF�&�^�GN����e�bǈzlַ�!�;�����n>���$��1�d,�� =�R��E[ 4�5���&���S�|#Fj��&�h���;}6����M�| H<*�;L�:�kɽA~�L�`Q4���2P\�j.˒���88M#_b�P�k"%���q�g��:�*���0��ѿ?�e���*�<X�*��B��(����ZU�oj9)x&�:ySw5aT: ��jP��M�#9��6��R�g��kw�nq�"e�q�~����Nk�����²�	���M0+�0 ��#	�N� ��2r% � P�g�?JR�f&XL�`Θ ��m��4�V䋐-�G�W�L��ԧ����/��S�lw$���gE�q5��wz���j%��h\�̅�_*57dfl8��,��:×6����;U�|G~�3��~���|&[B�o�$7�P	1���=�EcoR��/y���@�c��I=g�U�c��1�/W:�~Q�cMe�����c����!�nu2�u�-[���'�C��D�Cf��{�8������bJ���w?'�q@�'�����z&/C� ơ(7÷�Dz�+�+BJ�<c�c���* V�.	<nfokJb'F���(G^��Y3��:�3&#�s�`�z����G���R�}"����JF<�F<c���2�<j=$�=s�+���]�ȹ��@_�J���n��f�������UC�_�R��y�"Tx�����k׬UI���JL�VDɢr,ן��b�{�m�.^���j�:I�?�"ԁ]	����ܲ�1�s���<r~�f	��M��U1�"M���s�xh8nZ�tS9�"�u�x&5�م�ıJ&�_&�4\͗�����&d�Y�=�Gpʒ.eݥs$�1Rj0&+B�us,�#D��L���o������cL�2�j��-�lmԿ�gj�Bp=������[���y��a���3R9,�t�4 �o����\���)e�6�(Ǜ����߉a��G�A\F���㠂�\?��g%1����wa���&a�5�s����g���������,ˆ�ۅ/t��|�3l$� �݇�>Y'dnv�CBt���=�uԬ>Jf"v��Y!jV�ځH{���?��L�|�g�ʈ�/Y���]�'�嬢�j� n�y'`5|�y*#z9<�S�:c����'3"�O��9E@�,3�������@o�(m��e�1!Vh<������vBnY�3����nu5���5&t��m��)�I|c8��3�5�DL���4SbQ�l��e��z�QX� �`!F�/�~���O�(��y�W�,?ݩyN��NsW�����R����[o�b�9��H�BCz��c�m���^K7���]�t9��o�$� i�*�`lC�Rd�d�u�|u(��l�1��H�!��Vjc/|'h���jH�����*>
�t�O}(�ʃb�]�+e&|!1�隹���=�i�V0{��V�Cw��}jj 1�������,��(ƴ��&f
7Մ���������+�%Ɛ�\�޸ҧy+ �Y��m�1ά�դ�;�@<���&Z;S�U����3�9+�=y���/���o���
^��r����+q�Xd-�xӤ�iѼ���5��*X�;��I�m5�$����ҵ�Rk�sy:�3��^� U\��ټ(�m��c��:
ŌP,���q!Z3��wA-a�Ё>��c��`9O�G��]�ԩ���|>� w�s�����X�GPu�s/�k�I$��'Ϋ̠���N^���\ ݦ�x�d���O�*ݏ ���X'�PH�	?Η[��%��2��W�Q�o�9 �W ഭ����+Ҋ�[�&��rn����V1��7��l�`n2�$Ј0��/%��$���L�{bq�­+��$�`�}��Q��A-�DIN�gm��:�8�@Z,�Iс��u
e)1/��qA:��	���#�^*(@�x\�$�O*n�C��;�´��'�w�W��Ӊ�9�3�������5�P"��O8�3��ڈi51���q���_<A3�&��$\I�Ё|��ԚQ6�բ�˫�[���ʋu�L �`�&	�'�f�ŃKZyuۗ�83�pcm�@�畏՝��F'����n�0l��(H>ӡ���TKIb�B�8X��+>��׍3�h�� C�{B��d������v_�h�҄i�Ң��`�!�큫�)J��S���x�����p��7j���g-��X4 G��aA�ɀ3J�:=�l�R(�h(�ydF�}w��LK�tRt.�ϥ��xF�3lP�2 �u�@���1RF$�<����Zk_�J�}#�f��m̃A�N����#HS���7����
�f��z_�/U������s;\�}T�ܗ�������1TG5b���)����Sތ�T����{�D�Zv
���͹�>ȑ�Z��P?	3$���x�5JCi��"��q/A�����ؓGR3i�2�H����)�mP���F0L�6���?~jN��߁����ud�`�4��껗��Z����ZwR�Ĩ�W���l�z��_;.�Mqi��R���%��TN	4���}kDi��p�X�VVvn�>\�k�۾������$%v��� �iǦ�U�f �n2��#ٳx�+���6�.f��KUi��Ӈ����q�F�up8hM��Jd;./�A\<a�^��aQ����=��L���Q�~fL���>8�_�v��5�m��(@! ���2�9O6����	�W^4������Iz��X�����������O3%�V�CxIZeTB���1�EM�7E�-����6�Z�}�6�k��CO�Q'�Ń�0='�^E���[0U5�uI���75��Ɉ��Hy�]�߸e�֟�
�����_�6�Z��Ŭ}ٓ�.�;˥��mv��ˍD2��qL�S�����<�'�T��I����s���$�O��4���s=GE�':]�@W��Zfx!�}�����=U�:(�l�=��|�_��L� �!�
2Z��� �{�v=�γ����z_��~>�V�l�@0>o�bZX�|߀c0V�� G���Y<hzN���\82���l�g�����?W7��Q�㒞	�|�}-��Dn���K�)��H�sb�>�h!R;E�mJ�Pk.��1�+�������˒�)*�rܦD����DS�Z�Π�����C[B�A4f��P
��H�[:� '
✰����jh��x��D��֨��� 2�7���3.˿{�Y��zE�,��9{e8l}��>68�D-&�������j�����c��u=�`�j��1RY��z'#�1�Y� ��\l��"8T�zE�X|���U�H�II��sJ0��}�.�u/O�2Fr�R]�$���(��j�\ǜ5����;����,�/mM�ݻ���po�$B�m7�\lgy����Ap�e!Mť�W�����(�ݫ�Ǵ���3}3|��}8�Q���5�!�v@�g���j����ҿ���/���ч_��(+QQ-tL�<g��3>j#�X�Qknpw?���	��=�����.y2�1�Q"A~�����f2N��rRz��h��صć��m��ۃ36N6i|�;�� ���L��J����JaΡ}�Q��6q�y|��	�*ǌ����Ә-�&D�,ݩ��خg���֡;��E�r�#��8���&�i\%@{�1x:J�;�݈�p��o�}O���y�V$2���l��
�n�[�)Y��)�>U6���ح�ο$�l �졽����h����}	ulm}��R ��,���B����?2���b+FP �����0P����~�[�c4A8~��ڻ<hq:Z�N�A�!�*����n��x�j�?Y׽����X�0r�8W�d���<�3:��T;Yո�R^nF��E5�����u���j+[����C�.�߷ �+C�.���� H��k�� ;b�#�I��F���t�Ɔ���z�F�H\�3U%08	m���]���������K�ȅ;r.��T��Y�����@K�}^����@��]��v\�遚Ϳ��ծ�;t(̳����i���X-7��~�����omCZm��s)F�#m�D/��,[Z�(W�|1U��5�&��_�<����^�W��.��QZ��!M\�=���6������
�-�o}�T�>>��qB�?��q�l?��)��w��N͚eߓt���c����P���2���������Q�X>�|���M�Xb`5Z��z�������I��C�q%ң����S%o��t�����GT�}�I�d:#�<�$�e?~��������k���41��^U�b:���z��犾[�����ɴ!cF����R
��<c�Y�\��7�(�ҙX��0Xp��ÿ�~��TW�nq7р�S�=��T橫"�(x��R]=���wpB��f�ҿ�5��S�މS��L+�H�1Sҵ
�Z�>�-��lk��r8t~sL�pU:Xѱ��9���&��0�(E�^z[M4Q8hl�^P�=�.���!���� ��|����Z\���u�&����L��]Q�|�TY��}�5R��IU{�:$�1]
�kl�V� UJ%Ü�vq����cW#�#�X��Β�;p����`�U�Gz�7mP�'2^i4>SX$Q���e�t~o���?�o�`��
�Wc���_�D>��v��)���d�S)K�t����c��,�m��0�%���͂�"�-�S� 4|��6J����ud���9��ࡃ�+��&�8`BmL��!��7�d��{�g��R�uP�ԣKf������/E�n6L��{t����И^@J
HVy`}#�q��غ�fd������~TksӺ��j'����9Y
��*�*�w���ߏ^����z����j��Oe�]�A<��y�Oy�b�/�V)����\ֈ�9���@��N��=��$��<U�TN�gq������"#���Ԍ�<�HdnU�S����-�آ�Q��K��eu:��p�8_��-��r��O	̌&�<[�5td���h8�A�#|U&:ؐ���
�\��W<��MђXVu����X�bl��@���ivo�3���.�b��.D��-�Ԙ�˛�ט��C鉬 O�*�M .nqu�E��❑b����:��r=���#�/Ƅ��$�$1,�S�S��`���X�tx%�m/ͼ޶�,'C9�۳�'�a�B0}�,^�?x���(�R�l����0`Y�=1B
X8�c n{�|F1�ID�$._���[tݨ���?�ݬ������_��*Z�u�hmR��c!<���ȓ��r���<:�g�Ih��SA�)�MC-I����p_b�p�X87"����"�>��ˢ�Jh��j�;/�~<p���3�0c�`ND%�	'(Μ���"`�ªM��>ë�&BGfO׋�H2���u]����F��H�[j��1'������3�<zI�Ӡ��0�F�{|��|Q�R�3~]��oԷ�<Hy BԬ���4���d��;�X�{-M�u�@��D���@Y��KVR0��3�'��^�.�7V����,IҶ˥M(���f�ͧgeZ�,	̷�X�zj��l���0"Tj�#�T����+5�妃���M�P:B�i[����G�G1��l^��������k[3 �fZ���L��y�L˺���ߚ�u��,��J�w�I�/R��)ՠ��L\ym��<�)Y�K�(���OM�I7��"���e# ���\���xk��r��!u�e�eB)P�FMZ�l��>�\��	��"�]p����=��i�>8�	���>H76��< t{!� �+���de��1^����pCd�Y�LI�'�1�� !����&$MM��
�B֍� �2�Z\v3��L:�h{��]�^|���h�d���ژX$P�I{)[t�� ���;�? GJ+�C�C���⃰�!+Ø$���е����2H�FZ�a>6�dۯ����g���(͓���r�������$m)V&Z���>��7�B�\[��h}U�ڢ��m>ї��yxEImD�ahS~ �2�)6���C�JŁ��Cjdg��!b�n=��Ρ���'xe��üތ檾6��0:�$UJ&�����`�?�d*�#8�\�a�z���f3O�kB��	�}'~A����yIґ�]i�A�U��3+�H��&�����c�@	�#ץ9CC���~zZ�3���V�<%��,�#U�jU�z��iF��#��̽�2+��WY7��F��V������Kኞ����f���"OR�aיR'(5���!�B�)�����ǩ���1�{�g�?N/uE�3!�'�$Nd����OFR��3��J@��Q���\�LNF���Kػ'{���0%=C�����75�i����^�<�
�o}���QS���'��m3i�'jߎ���ESB��|�ڇj<��ΉO=T�'<�+�"k��������W~�C,�EG�,E�s�1C�NG���Wu�
A��埒����0���x��>:�k�r�E�?�%��؀cpF��֣[R�ɔ+�w�F|�%����?��qf�|&�^�>֘��^�����R j��zOddž��Q;@����/8� ��>� �3uN�T�2�|g h�a_�qS7u�/��>�4J��l�6����0�-�K.�z8@��Zd6��d������/5|�|o�i���m1�F�Uy���)�FI�k\��)�q�l�W�}5����Wz�0|�l�/.l�SW0��8~$�2d�S��%w�K�im��Ha�	ޣ��(�.Z�D4�l���$
�7,�6>]8����S��ح��)��<K���N�ӕ�ђ��:��~-�4h�bN���,гں��!��ۖ����	�+��7���V�^��E;5\�x�������~l�fE��Ms*@��������'n$K�N���X��m�Al? ��'�*ϛR��.����	ס�o(�B`Ó[ݶ�g�j�'�
�B�v�hw��`d���ޟa�ӆh7�N� ��m��d�M��k|��$J3�\���i��:д��)9�hߊQx|7'���&�w^W�c��B4��H�cV��?y��ƈo�R��&�@t�`�F��3e�m����z��,�yP�Q
X܊z�I ���>�_烃��W/e��
=Í�ݍ��A�I�`q� ���S��j�#|"����t�M���wB�ۣ?B]p�!0r���خW�!$-�޼PF���&E�J e�o�KZ30}�p԰	҆����>hO�A��7]��Xd5��8 ��V)}�8���K���i:����Y�_c}T���Ƒ�i]�&�ϕՎ�D�	.e���D��
�6雓��:������ڽ��I�N�K���@��M�:><K�a�&ٲ��v%ȷ,c�X1A��sJO��R�6 |nmTԱ^�j��q�|�O*�᥿'/,��+��E�cb�{��٠�LB�"&И�����B��s��Bz�^���z	UǭYRI=�\�����.Up��D�k�$�A6i�� i,6FS�k_kq����ӦA)l��@w�q�ݙS�򌾕.,�&-37:嬲2T��;�m͓�1�wG�D?5���@��X&�?j��<zo��.vD/x{3�ⳏIJ酋�g�Z\��B�ܩ}AF3�`m��Dj�9�t"QH�P>�w;��,
��縓��k�/$.^a�Rt,�z�9�����(��a9pw���j�sW�yG����n�����	��-Z�&Áʌ#�7����h%
��.��R�q�7���z��
����/�d-�)��N�G��{�#���c�<K<���'op7���1������|x�m���;���P$��[z�gd���Ҟ�`����2
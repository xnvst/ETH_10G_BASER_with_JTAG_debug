// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:23 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dByIrKqWANy/OHnqkZoYZ9OstpIChbt2eyAQU0D/g5jqYvTej7IzBIf1XXX2kcf5
b72/uTOVA9tdHgICqfvS0LhQJJW+WwSFirQ8tl8RsDmFYOI90tauNnCWiqMdoGMm
J7SjFpa3QnfMpfvFwW2LoYT+9Z60DUkSddwrkEAgneU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24432)
/+zuSyOJNpBIWDVH0W8KAcmPbuV6NQz61nccYU7/eoPAm7kYuiszI1m3D5jx0+G9
yXa4fWVuaPzhEPJNa7dN5t5t6uVx2vjph8UJb2lA5Y5yAjGtl0IfzSXooBgUUozG
eIYpf4AePoBmcMET68PFTWHzBd1ja9I9uPGU0AOT3r75PDBUj8OZJoXBUnAkEqgi
jzlEnsXTCCDRHnziRBPOEIX7THw9CSWsQR6uii1zIwFtKxLNKF6CPpjP99hpaUJo
WIQi5wRQI6GJiGvFnOyu4FcLGw9mEncMF3NnhbBdaosSAGqsiqjt+JR3+8AfQ0dj
qg0nUWrUYdRcasFiYi3NYxF1zDYqMHw9+VI1rh5RvcfAGWkiwtP7vF+WiQFkZKT/
F1Vf5cybyECxu0n5fDDZFQ+lHmXZAeT/eorWvfrH7aJ1w+ss8v7cLM8cM72qRX7Q
WwnG1AFEtZLwaQoucrU42C9tLwXM/OatQjOmnwd1CAN4eFw+/36AsQ1ZFDxj6pFg
hN+kU6RIdTtvmvZT9LU0IdutPq3d0tog9r7AyZpjc5ENGCpDDQ/VFEKxlp7BWYeN
uzOtIkUBduo9FWCJKQShdx0RCDPiA8U3hztu5BAQg7frozBNDyr0qfOLAjmRqMy9
fgDImYRikaY4rG4X7x+OpWuATFM8kePEomg5FxUsJ4IOCewJcoaqSpP65J1r6XU1
kOA3eP0kBIoOCGUdfxM0VmUEUUCCBT6dXiyv4BuAR95ViE8+OaEgraWISfeVC1+Y
VwG1n73WpmmchnjU8KAHKqY8aZ0JRgSiVIPKa7HwSU7f+CxKbDZ0QOcT6iay+MEx
hyv+6zEIWvTSsMSuZfG/xNA5IB2YgM1n3nmDhr2uka26oztqm4OokF8AA5ObflmO
J6kUfGYf1m1xVRgpQLbPiJdSciGupu5HapaewT0ialjvK96nAoompIlCrLxu9Pqd
f3TTWEWymKtcqwpktV5aN5o3XPFiqhTOOBCC+2jAPei5qsKSGYtQJWAHsR/gxhmq
/yScQQhuaALog/YTc8vHpp8H8OgFrjgJP2Vk7OyqNVx8PLhx5RW/59iafKIhMoLv
eLxaqAdp/bhdragfpGQyVFlJ2+7M8jYMYGWhIZ1SLLhNhZHaG3CbRo75w9aPajvt
Ls3sYUyLhv7BMGa3ZR2SSNjWb2UhMD3Gk/8spcjPfvGgX6O4A6j3G9LB7ftCoQO4
P29liBp7LGPtB1ltOm5ft621xyi6Ro6f/rOsF0T/n5cPuCEPlXtK1cHkfdK1TpkP
Rkbqh0w/LdPTvw+8wFoGUlM8hDwUN3NzKVj6kfoKywtdEmSjfTUwdez9UAojaxY7
Bo3Abm8nEzrTqhOA2UC6nlAupKQ+oS/CrlspDCvKCHDzHVO68uoq9O996kNE/1zU
8gn+/6vdsmU31qTAVY7gShyLDQBmvACwmEcqanzijMQ/0Lv+fj9SrCENgtWm+6aD
e4MliPkIpkXm4E9K7I1OgQfi43XRRIX65R42HvfewD+UstevaoL0Pr/c0wSLtj0U
dNTqeeCtTIX2hXFxzd6vFS8hgEPyCxw0uzTadhYJtSxkH17y26yb93bqJKheQqAY
VADRnfov5LK0Nx0YaHUDcy4vWjM1i1w/itZRHl0iR9jIjvBgXABSvUngjNGhyM5z
z9CGKH8bgp1I0lhob7mjxT8qypiatayTQmez64K8It7l24RyXGtAOX7lMUhd12SP
jYxfbThGtbnbOautWMTq94462i7SpIJ+oaZR3LEDEg0LFIZNkqFzbuv2aZjz2eUo
3v5gVymTb5swQ+RSt2tjiwK65uFMmOzqSoUFaFnABwDtpgSUCr6jqPBct/wH240Q
Ejeur+PBJNUKhF+3XkWMUv1sH35zy1fIdeD4jBFPS5CJvmah1wOrHahhE7+qJWqf
prnEnaD/c7m4RmVIdW4tkmJNAS69vzaUDMN0GG3NsJ73j/4wsera0LyXugpHlI4t
KnKt7nNweZgm092KQPgePqGbSZ207htmhu11ym6peBzDaQxrr1YwbD05QdfsevWK
4mUsboNDr78kGtWOYe7EP03q+JZP+JQECZSgqVk5nyDOgO7aM4OuXV2pP9+wqk49
AKhBnbk6UiMGG/XqmBGkM8ucaIBB03LOVS6kp8GqRoyjTHP8Mn7vbToKdbHo3nNB
ddWd1gwIcVW77QEw2vPI8aYYbyMCO5M/iVYEWE7lTT8aTAWIbwfMZ8WszjJZQ/Ay
5olZkH+fvI2FWAWD7g3MpbRF3eDvC2KhAl4kHUi76XER1TlCOi/HnEeDNGigtQpz
Ie8LvhIKR58BJdbH1jdaov2a59WKDNaDtzxZ64fTieRJOcXk+t3zkgF5D3zxETEC
sbAHjsjti7PdtpBrBtmmQj8IaSWvmPcwFl3nXlrYSoZsShVczv72q0UnkVeMFYoI
wexdE4LggWysLt7POTMvNx8lB/XctBW7aLEo0A3z8Plf1GhM/ODQgvuR9LCaDEVE
cufvCsE+VmwHNilwuYhWCo0y3R+vLd+qsZJJO7TBsbeG5s0a0ft/60qzxWRLnGNt
tdMjxxiytSzZWgkqDmA95LIKt3wqhaNt87WeQVoI73C4VYACAZcPnw1PEKA+68nL
9zRvlLvTEJwduhihTNI9+AHPpEuaz/kZoFxUX2z+NW1VpgG4o19roVE0itNNBe/f
OFVw1a2Dl4SWO2D/rvOKzleYAniSP9Z90HZvdp1sUyeQXLttAFuxfh9qV4kQTgJS
7Cyy5MrwulgqsfSYJU6d4xY394W75KTDC08GcMj0MAVeX7Ia5UFIs7xfc0uPyzI9
MZzH8zKWQayrrdsiHHukSY2qmPi1AgUfDH9Rsrm0i8hC1n50sbQgDKJG4zZc+uV9
KX4gwDjrdZJl4v13MC1bDamKKwsKxkIPoOB5LAC/L7TTzUbxnXULvxnms9+PfCdZ
ICeK/hNxDj9L7Vp8B6l/vlDNae3sTDJ1vtpnaHxHov9MnfeiSBd8eXAOE4JjuE4N
eP1OkeuOolr2hA4ivg9jrEcbZUqPwK4GbWsOdZq99ueaaQrguaMnrKsHSEH/KUO9
Wkc1hjN72vTKgZr8k0NFN4o511zEEFxJpFrRs/1XPX73RShbaK+B0IDmeZ/Fk1a/
Mcsh9S4mvQJfy0jVvo/RkgNSsZBGEE4tMTK3GnwitXTVAsry7AHVXeXm1I3mGtCo
CW+Frt5T4izGoOARpsG+3+n3sfVIAcEhtGbwHH1nxUlqB8BmyVR9tW9yaeG874AZ
MwMhi0GB4qoXl5pIQMkY6PxvNFMC4hk+HRAn7h6OQTqyrrHfjiAb1VkO3Pz5ykPy
PrYARPF4s0BZ0qJSjFvY1Frq9C+c8ukcpHFcF77KEvjod2k+oAjmv3aoK4GFUtBx
3RSvxSqf6xcBDvRApDWfOTrGyUYV+vJL/shLlJnlTxL3lvNwSfGi1Y6s6UUjEX9C
tRTTvP9cwV5koprtB4pAEmU5El1fBehbHURzIy4tCj42lVHhAt1XSx/cTz9iwvxQ
QNUYuwclJgYNRkXp+oP9Kv/rqycEimflR1It0jZhhuSlVs62MaQhnzUmAT4rjilC
3HMWuLyuFOqDZpdyUdspNlBwJvbpBA69zM5t1UJkfTHpgFfakiRTTGUjo+e2Y0eH
3QLELcyDU0UOO4mkA52Bf5a24sMm3bgNr9sD6ICb/XBlR+6iK5uh34ohg655yWWQ
JcFesf2BCOzq/eenLSALIyQcNw0AaBScp1v0qXKVWSE2Q+JzDNiKMlnd1UzfDpVa
X3l0F2BFVQogiU3Q3nNldNkTMzMyIf6gl36KFTOFnkcQKr9ToIBpuQHnYbharvWZ
eEhWBGsju4KSFg1TS2/I2/uQzk+OHANp7MsC8kECcAu1QEeoS88NnSBxDn0efTiu
vYLrxYW1fTrhmRbPq/C2TZU74LcNb1YaXn3jJNkL58TnuNRtuQsTiFYXi/iwmd+S
6gFD/BiicpL1gZB61VsG11w4zRUw6wqPkJ45T82tBKJ7z9OEsvtt3G1rloz5r+M6
1YWacdyKsfK6FVZtuZ1u5r1caIoe0KOasHeAxE3cJjhOiGqRqOpx+VsRe9QWSUbP
Y3XlGHBu0l0OuLwLg+xnS5Trljesid808KCa92+8tHpVbt5qiKt6f9o1aoOLdvWK
x08IXybzuRnpgGGbSDuTYaRNhXaxPe7bVmK7PzjZ+d3CEUnO9IRuX40Hdf/Zved6
7m3KcMyp+Qbl3Mq1+vZwLCX8d5+hwAofGI9YtgqrIbbAwpxIQAp+icop1CFXzXmt
CxFBd6PQkPcxQxjRTOeE/UrIK3JjG0+uMXrh5Yqg8aoKgQgmDW4Xh0oUZHAvgnpW
JRhxLp354EAlyM7UCvVqzkafGLJGiN7gcxMjGensYMay6HgwwdhFlMYiDzqxBHiC
BL5QNBUN2k6YvFwmmfKS9Y4zdBiFT7BdZJCwBXvtHBhfjAS8twTcH/mZGaK+lLOg
arHWcxR91ulFTj97+wzQ4cLMwuJJE4hMOMRy5LNedK1xfBjZv3xliCDVxmQy8Jb2
5wlVNPFvkQAGy44KDYySRBfr6ZUdhuxscnaDgj41CMWhFwN7oVkbd9e9NcPLv4B7
qsywRpgBOz94ybai5hL8kBuB9csYbh5hG667V4Z3rNb/r5y1LGI2Xjgp5sas5HNR
hN1Gur3DM/JOVRL3FTvnzlPQdXhoZzyvRsSOqVsrqufC/VZeQD1GSESpO2noe5P5
LJXuP8JI+59lNpP8Fp1LPu3CkbjGKfn77IjXg1+QnRj24iuTUyXcCQW4Nqpitxdm
p7cV5wWw5to9+l7Ceh6XdT5hGzyR/x5iRmZndVHTWBiaEbsAgE1OLbcrXWk65Hxk
9Qezzjq0DwVYgN0WEXPQpyVMibyEV3mzV8WcQhE+tIY0Ar6zwCTrVf4jbOr7C5/8
uvTXGMBI8lvIeYMc5XcU5AH2DMhvxrDuvVdsfuDjrMoeSGTbVwxx3/7EK0/jJOVi
kUW8w3VpgYpDoJPZ5D2Fk3Ibhks79bAQG2GuiADiifwU63/iZb2H/xaOeyBM38q8
Qreyba4suPwMCxOhrA5/uv2zsXDZH79B8BI/oSzY0ilXCHiTaJ+lo0x8DiMJhsD+
4cBHYpSaIfWP3pgyhp+hOkG5OOfOAKgbUOjnsDbDOTfOKMFqWH8vtCLUxZm9n/KE
OQkEAggZotplwjhksfHR/UOj/uyK+vQ3k/4QA1WYabQMGVDAEAS3ntJG7vojdcWQ
O/8LgjdHi05D6GdLFaItuH/rf1288uUcz8uXnJ0FMap6E8fhhXk/6vXqswEkqnJX
c1wqi/CuWMXZeOa0xBnZo7XzXbre9DI/7GzMS00+MDsHY37XoKxTvPPgy7KhN8v7
YydGEp+HyityKBAOVxjnu63bShEQL2wOdzx+rLfSYk+Mq25JDDrwDEz/+f0Qc87i
LvL3130xmAZUR9b8jISPuiYsT/fUgy/ErIvzuPHZOxsvayA7KIoXhtqaAx0HH9Vx
Wp2+wnrdTX7diZ/vcdIOnRLEZKc9DRreKB9J830aNrbhr/PAWZlZ+7K14bL9ps+t
31NTtU8C57nnEmZFv3kU5N6NHCJI4h3SC/xVkB1kMAl1RS2kUAltaiCB5EWJVNy/
ux7VlH2LeaO2jJ9ZVEHNEzLjt8VLbPJEmwZeY5a9gX44zxAmyQEjiLBNQtXZSwwU
IYWQKaWTz0trl9mBuKFqJPPW9YUKHJuNNj99m6tVg39iYhgK0wHDw6IuoYrn3xNq
j4vAIVruO5XMdmLFiC8GB8NRn3oYsweJBQBX8VKssFooGNoel3dw3OLFYjEqjlb4
IRLedQi8fOXeshh7xRGQ7RI9DRnTwurSYkQ/k2BT9ORfLR1A5BXyKajLAfTueAfm
tQ0MFa88H7FWIfUYrRvu6g2/r5qUxtyk3mW2F2IOlNZO5qlYXOU1S9krKhEgOR2y
pQJEqlokgekl/Mw9lq2FOmdPefoLA2q2Bj6W8C/NrkKThDMXhTTfCAD86fy+6W3J
2OUNNVBjwnQ8JW0IzmhL3XO3idsKHooy0DYZW66NeSu4UVxiBrKKMfZu7I69pS46
tnO9M0HM4jK45/7gouHSGa5D3P7EPGndTUgbFI21OP+XrBxgM+5/0nMI6u0ovx4U
IW0yyUbiPsq/qx2DDfWoceI3UH4MTex1fYHo3vMj9gwCGLixpr3fcVKs+8xxsLUe
LAxmA6T/0UAR4kFpl57cSVvAYJ6j8J5IMJkh49apWsQ20h0ZsnTue9XF3MI64PxD
sJS+b8osoErk1VOg7pTf59h+C+VqSFm+RXe+eUYhODI9aYehHtPU1XgBE5DX6eB5
kom0Ee4CSsix+AhjdLPb4xZfHnkQ33nlJB4ywBRnDGGmzXzI80reR4OpYDBnP+2m
3/VXWz7lEaBGAbKYceMbwOVAWZN0wqYhyh0WzcQMeYb4+w+dC0eaH4VpeDCCrZst
zPPBfHfjLGnTl5AEJYgL6S8OSHU1KQ1ATz6xTNn3ZrogGg9A4SaQvzO4busMIdqR
1l0F9UrcvEMKHr6kIMFiQTSOLjKoUoK3HCFTribGmuhpQ/QCTZv+EZEIwbed+ea5
irshQP1A2ioum0e15PIpzdmhSJVq+LfaNmqu6zmSLno4a9lSZ2DXQFnV/0/EfhwS
3w1EfZ8oZ6QxrJ6j45qpgs4ANugj6kyPk6GQfcufWrb96WPSgplnmnfYdiQxmcHw
fNMXUOXSxl8eXDIdgSpRhJ+djVMlEoJ8VLOMeXvCq85kuVH+MxCN8OFCndXcmHao
orTSGxGuDVBJ73PjmLIdy8DemlRif/sZsLLPHUK26csILdTkoHzx+pwVfECw82pt
T7EjcHYRZWEnC8PFzGQ6m6d4V9/+dPSv4u3sfRGrfcMojm5wQ7Q3FDBJqRjeerMH
r8xsDCdfpYtdr43BAkb95eC7QW39wCeR53YEXrlez1N72S09UrCVrQ7sTOK4Txyq
h6oTtCgmKeVJ+yXTfi+IuFmFIZ1GPRYKv8FwzRkWVEl7QrdXs7TN20MM/XhDUQzg
gpUledX8AY4TIt1yZE27EMpUO2NZVcUfwrqlsaPexrMohxE+ajh0vD8jIWqJw4Ic
YEG5lbOCSN7BbDbOG9KzUDqCTbw7PPSEigog4yKOiamM1oGMiF94jBZX80+hC0dX
zXPY9Uk9nu08Nbsu4Cp3ApN0DS3o4VD7MQJ+X9Aayhz4UVuhld9A2yU5m2guHgfb
Nq8uoWIuMk7dVq8yF32OZ84QL0cZZ8ipDMCiG1Sxg+naZ0Bn03bwG0upXVW3rNrq
rSuSXrKUWDeClQTRCZzwoDqhb7TtAT1T2HoY+gWScyKHtZ1JHr8rtXCd+6TzzwXE
RKqP58DGOHxYsiHV/zYIxqaW3mhUe+6+rFD+gegYIqFs+G3aqt8vhhDuGDh9jMpb
Wgf+HGTrFKL/sD9nw8SDOkDZ1ceMtzQxySheOv3rNj0zvWF4TQKyxRawa7n+BbyS
mXR8j4kHIqmGb3JdjzkbQAThD0JT5rklznkhWOru8av93yPSa1ajQW90SihygFu2
8UmmYdvb6XYcSXuoGCrxZ/kNjty5feUgr4TJ6avUAg/mzqO3Ve4ssOmALU3t0Apb
FFIGSdZlI2xwppAbhHBtd+1lXti0Z9Ggaq/CNDLmLTft57RwASkATZSqY8a4tNvs
MTLYaG7X8qLes5SEyxDK+cX0F84ldrXPdhCfWeEsSiSHHOa6xgs1AtaKFyZiss/X
O6go/DiSOe30P6VMct3tHN5ZIEYUNBpqZxB0VNqJqzrnnraosgFRIdWHwxqkBL9V
ONSTMz9l1moxloHwEi2A4F7KU2WiLqdW1rs9rdwtgDNPr1N0Lfli/sI/nBYanK94
rgd9AFhDA4H0pYxRnoH05gGJYdipeoqjNVsqWSMKJSw0GZWlin8yTxufx9pgIkSy
et6QqmHuAuwBxudfnt8KY72v9Om0YQBTNYKr1yhBecP+RDNcURnZdgr/0ailmATG
HGx4ddaOj38B42vNREI5f3s8zMdqpULuR0c3gZ5aXwERV3sRyPoCm+YrQAwHQCOf
U02qP5wJDDmZV2821vQ7XDCarJJGSpneAOwZsP4au6fefXS7xZV1bbtheGWFvir7
ONLwWq7NJLD1zK6qmWmWLGbyHZjRVxgC/p29aa6yzwWXAe/8DGrc/ivV4neN6mxJ
3iQ6g/a/zZfbf+9BytnkIADmaPxkNTnL7CHz9x8gRYf4NnQyUKTzhYEj3UmlQlyM
t5vQjsgl8OvM297Q3qgt9F5edWxANx09x0OESVWm62i07HXNL3I3uDnc28efpYW6
o0tLD6EksvK3Eb2IHVyVAtQ5EOolGO1IMu4SspN+0HhIBJjiZ79w0Eg262v2iZKq
zkyyBf0OsM1y5emloLBlKRvheajksnKkprM7ayIFf64r9jP0xbfD877qLK/0UBqS
FRaO25gBTxP1Tzztpafkx/ec8X5CgWfR46o6c5F3BKU7RC5fsrQ+DFpXy5G/HZr/
pNesicAnzemwOfEKKB4+pI6gmlKgO64K4un5QxHooR78cKauYXtx86cdJIAopCSs
JBiUVhKuMAmIfwt0UMIUJSc/DLzcSQ3lLj1bMFHwobkVZBSZrZdH5os++ZmUbjiT
hPhcvr0V3mmkqe2YMNj9ar6LmCIlzkv05MBrsFf75M9jb6IVEBIb0hOq3Pxizcet
2+1MH/J1C2LD0qvXSK0d2OpWngaHjAmrrA5JXrZVUouwATAWym1ImeCpgObOmLvL
Vs0IDovtt2kpQVyo1/X8qBuSKrHELT0zbnkomyFKYx3N9qJdzv1K94cbCLOSDrF0
ISkDFg9UIggI+dVxV2w9bUBRTjC/w1BrWuSgjdIYU2CRLqHW2Q4Lw6EkFy0qPodZ
q3Uw3MBVwfTuzWs9fX3px2Js7voc4fWpprpMq9aUAaMz8sMXRRc9juYOyo3E1AlI
1Bn9g5Buk2Ren5ZM2L08Gos+ogR7Uyc5CbUuW0+GrVxSnN1YOv/9IJQYVELKstX1
hBujj34Hh5BxywIA+clGd4vwUJFHhHT0A+TDUQMNec5nZfbFfaal/sIoqO4RVirj
R/OVSnXjOaXWdSD2lWB+RJHaE7JBMtKq9X9e5knb4EONP16ghwOFMWhq1rNk74cB
vaBf/iWSPxbTf/+AKvRDbJWKsLEW5c71jJG7axHiB2bWtvBPHvw3E3zs/+BIdwpY
oru/we0ukgCD99kr4bFDh+TOAEZD1Le68QVl4J4jkqu46LyyB2jGbASsiYHvE15k
QVSRmcyWabrRs3/85Ka728F8A2jXYoGcpZDOeP5V9alHsVRtRIIGv/KaO0xaq6+R
8/+4b2ztftlMAbl7E+ThrBmfmDGAxvg3V2pu37Ry7uRmHYQ8uTFmOAk/HHctPMnr
He9kmdwwLie9oR3ArQaE59uuOl8d8CuSZ9/4q44F/C+4zpWJwDmLrUC5hkILsa/U
v94cifeLp4OJ7SiZ5d/ioNUvQUAl+Z9M+YDBAfe8Z+51DwhytqSy06tdCqXJpPOJ
uHZfTD+HnKszmI8vpWzbsmeVcoyHVqanxtsWGsw9JXH7U5VbdrwnlKG802RgEDgA
RUfWLM9026L9hX/wA3OlfnVxRViRG35WTHv9W9D/W+8ujZ79k53ieyLWlo0L8JHY
sTPCEniqGXpBfYan4n7A0361fE8HifBd0BFw/CQuTPGbp5xaP+J0hMvu7JbjhYhE
f4iOrSl3oXcPG1z01CLNwEn57daDjIKWEHykoJeT0IzYYDKEvkvJBmg0zz4L8OvT
IqTxs6gFcKG2zk1tLwK+DBFkexUy/pyYFtqVpTxt5N6UW7hTqdYffsJNUbK0qyD4
HnrOR7AXgFIEfdAdYIEforh3uwiTrSqOCLXYuKVl8CCqQU9hVMw1Binau8sssVYG
XUYI53VuwQfmPVzFiUFOX6oVRXycA959TsQLYqknBSZ9zBKqBbHL955K3EFPMHe/
H7AfapqWczIKqelTfxBaedEvEYL9HpgRbkpU0YSre9A8UgEvHVrxZLADeKJ45kHZ
sjF4PdxJb0mpVd9T5rJ5mQ/9GeNc4EZwJ3pMeefR/1Uj/YaKwUK2tCPU+M2dIhxm
IYUSwLWCsF6u0Dj4eWEnz2DFWo1gfrpfhkd2rPp4fQkKnb2nSKcdtIwO2czXVysI
otbqeVoEWruyhnn5o25KDRKu1x9tNCUBPTIJGuhHu8P6TE45a5q96k3bbQw4z/WG
jMCdvFh6J9X4zjTwwVQLD2UmtJj8LRl9LSie8s8eNqLix1F+Kvt5f4Rd9oXV482J
WxcYHdzgKyq9pDOsjJCUn6fwSvol36Yrz4RcfiRHM4qWh2mGPrMjoANeP9Sgny5l
2WQe6aOnipKnmxr9DFGYuz0RIagt5gvJVE8MUFWAdwEHLDkgo+kQihnjQrs6KjF+
iug2lDCT1+/H3OXwYQH7r80/pxWy+3SzUSQkSt+t/BlTxmYuWlHu5bmD9Ae8T94e
47BgB4jB+0Ep7vORtzMDMk/QoUGxIt+HgZBBPY5NBL0YM/UwddCfhdStBYT+hKgc
zj1G8eN2Z8wbuEDhzd+z3ODNThLNg/tx7+A/2O0xOtjQPV76kR9zH/pIcfzph25A
D0iNkNVCTzxghO5Je9Q20E156S4Ic47LltA0tc8oHVzYT8KNVNtSP24+aU2FZDi0
DDeSbqRpYJ9e0thLXiAiuXf4B7OlJ/ke1gJTS5yCZpqzujX0EMA/+1kjp54QpoPP
jvtgpsDXZeAVQ/vgvLAvRsHut2YGTsfk3jjMQ2B/KFOJjcyK41fODLgGPAImL04v
x7m6Kclz87quYqwsAV11cRGkslTuzg9fUW+3eZl6Imqq7fPUtRbZ0Avq5E13omyk
qtyV2dAmUz1fgGT8MxcQLdEPM6FUgyUNu1zCjwu76A5OxC21/R/k0Vx1lmPrmxVB
BQdCvpKMRGyytE/bvILqp+So+G1bu1GDPm5pQ2s2ohrPy24Rq/9R79sOeOvnkeMW
qlsmqgXrT+xXjgb8KNBzfYhNYd5/urC3K2wPluGQLWy+AjBXPmxzr4I+neyvrID0
4UjR2813eSmn+Odcfwdh8/LWFub7cl1DdiA2bYntPMW+lplfo3hVVplJl0Vup7fp
KI4gdebGZCurFFDsRHCvVKLmWAoqSwom/4Al8jUwZTmuhjUOWI1S9/Q9wwzeJMTi
OJQUU5DgKoqI2BIr7dnhT4GQaKcg4DZa8rC9or5EmJt8577/pCb+VGPhgPdlFPoK
55Xz63IO4aqvCFrM3WwH249Fvt2pkeiVGAiVRsysvSp3t94yr82HGrGsjTq7ziSu
6fa6+qOZdQDVAiDSiehylAGD7jzZdCy+rfA/iHcUPbWtiXnKmG4uiZt1yhR4Mn1x
wWHtARCvJn+1LJxgs6hINDyo8PjHyM/9BhPdcUFb4po3oDM6mYZJEYRrKtIlZBat
/AUXskJeNojbMCP+c6/Oh0lVVW56A/YoHRHiSEfYFn1KIzt5kGNjeof/liOAadiq
dW+GrK9cYTiR1kKIeUbWfYU4GZw6rpYRfjJWctx8YgdJQ/n64vjZCAhdNF55iGPi
j7ZxeElAlh/h3HMKw1QwGCSQBCtz3V1+B4TmBPnsFPeJycKWPZZ/bWoMI4Rk1gS5
oIpQpJGLlvjODFyUTtXVhpm3P/BfRRTf3rxL5pKVc/l4hR0iz038ajyY9ccKpnsA
FHbjledlxbMwFhnaTr6rtssotUrKHRoxD33F1URG1Eg27aoOA/ddk5rWq5hO5YLx
C//4qN6+zGsAng+sVJ00s6UIBc0hqT6X8CxxjFV6ukiz/hFCW0gAEfU7b+ctMAX/
anEzyIjTOYc50d4fdXhwVM+ogfQvNxEdH+YzWQ7leIXlv9rc8yKRcWQxzLi8TrH2
7bAZx6GpFDAUQXjM6K/Xhtm4qExmWdxzqAlBYZU3FF5Z8fLbhWY/cVqWiue0827R
taBi+tgOxa0EeW4fMwDDs5gotc9jz9nq9pA0HetwDtj87b6xDj0GTY/na9Or/zCM
dEp1FMqn2cUKioXW05cT3uY/oaV14akkcoMv7uQUaYu68CDSrqjvOqQ5V/7dmH6p
lcDEwBu7kPioRessZq0FdfcpcjDHZ/eo3upXkSw9pJIALdnPdY4DZw/sfqLZcxqJ
dOHRgOY3WdpN62s1YPULXPDuIepIj5zmPHtxFmwG5vhXttiOlQyliVFZBlb/2zR0
96xCRCds5m1C6iOas7w7CCDm6uoXb3FoJoMfo8fy7WVenb/i9oyQ110+f4o2OCLY
fAJ8fU1YnZ+7ZH64yCRtfpECTCv8SwWlJdEpw/65nZtN7dXSo888GnmT1kJJrYp5
s+EYFYodgfc3SyWIprrYOTao5TLupynh6vnMcNPCX2uORndcvHSvFOKtJnR8QPeT
OWGXDUz+FPFvmwLaxJgY35Mmhe72VATpIkg5x6YI5B4MfS8E6xMyAT9P9mcWiiIF
lFZqexWgfc+LGWgIMaMuPq+qy/VUVoDRPZoMCdDKmMOcgwecEOci6VsOrjV/UwyP
kPffh2e2W4X07g/G37dxYRlFKPy7KiKxKcfoL1npZU8/rED6Gub4rTu2n+J0tlPJ
mVbxqlUN+lfcCHoukZTZPURxa3Ui2yENiA50nQefLASHofCbtoJKTHejQ2AfgBH9
di5P8dhNWV9gp+PlSaA+tOUSk9wxh871TaiO5hyIR3e33hrFsaq1tn+lhCGEeIKv
YjEC1xIeaKbwGQSV7WMffgi5wsdJnx4i5wNQ2Om9p4IS63m214+c/qA/v/+7tK60
LZe/EYMivS4d8b4znDVykWc9n6SEk+i2nZfqoLwD6E7llHTYiY4Dvy432x96mS05
hKgKNU1lqCP8JPMG3uSypw+LE30FCIildZ5TIRDpKAyKGZUFvNsDvhovbbUdgMoP
Ch6lMg5/HCUYODQ2ogo8hR8Z1NAVVl/pYq4CQzmd9Yhc+OcVo7FP0V9VgORBc5Rf
DB14eV4Oy4yFvfnP38xcNg01+1vZqjhpVTjY1qyEP8KpeSim8a+fQ7UVsqnXKYTT
PCFsT+2YepiaORw/oetv/U+mK9ZSbEMIBF59PtZBfQMY9xlv2BvldZ91f3ayGaUX
wmIUYQe7ZhPEc87QUUz0PYnhy42czn5xahtagfeF7cS9cArRIPc+geRjua3Q9C8P
zwIDmZ295WXgusgUJo198IDyjpqtxZVwcgEk6VXlgPjVL3+3xzSlRl5H2QnLpGdB
eUgPcJNLwPp5Pc1zMATnlcIcUXbsB756ftONjlkpiLRAAX0M5FYyMTmPsrMMtGXb
VsvaJkgJ5IFCziWFc8UdfJeyTJVMXQ6VaNN5I8wqamq0yOzXthFuuk5eYZXr/HLa
Tyj5stu4kQb2Fj5mCkpZgB1teBi33gITX7htSlPprsh6J/Bbsf/78Biizw2yxYu2
ARukoHN5MyDbsWDdwrQ6H/7+sDHyYKiJA1VGycy7RiCZI7kp72s8cF+38dJ+hemQ
jovrnZ7EZoM8SOWv/XpFfFRSE3xMgYp53sfyDKqQ+9Xk+uwvLy7u/6/S6pf2EVdg
ILnp6oX7V+ahEJle7jAd4AGsRI2gSRbdS/yly0W5R9RL4VGYo4Ux2tnqfA/NpHO8
ewiATQRssPNXZlj29YW6D/prW4EQML3oK5AuO3URzgnSoURSab1lZYKyBtrioCQF
bdkOS6Q4l+j28zjgMA9tvhJdeOnD1DT6njg3iS2ogTp5dMtL+GeTPubTR6qqrPs3
h+eA86u0swu80GGv7bLuCf1mIlfy3ZlmVeV85Vz2AcLzXlT9Y+aexDN6kGBtPvu+
k01N73L19z3KCToVhTnnq64Svoz2C0UIlESzWfsb24A/FZkmWp8JU2kxpTI83jVJ
R+xobw4E70adZJB/+4c5JfBmoU8Fa2/Iyn+o30ybz28uXCo+6HqIPL1ngsSmJS2x
tePjbuljeYN8t6KXxeLa6E7Rxf8cMadPbweHTT3MzPqOOQ+eazB3q6HvyCuzHjib
tYI2SfbgULwOhXxvaAl/yF4LWRlRvAypzC/X4h45f/CAwQX2I4orfpCbercuDotX
S+c9tkDXlZpVAK605q6HqS7q3AOr1gFyJS4rqaYYaX7Kb2iKyWuuqruOIKjxXywX
qwUPgJN4tsk19RqymDoZM8upZeTuFFaj4t8tuNxlvjvjuRfnIGAZLYANYiGnSQjC
Pe/Gs4acnFko++Rkr5hqHYi0ZQ7ln8gN2n280DQnQX5yLwwen9kP3BMpPsFauWxD
lOIiGssrhFwUDVyUVSDurLwxYKz0GFNeMO18+WoGgN1L7SRuZCT6bcL+plMTLhHI
hgSQWEh9kcvuYgPzxIScRGxmOCq6Z2y3CRniEb8je8BUZfx2LKGMCEQ7oIFy+9i4
7eUH6Z3qcfScAddtFDy6P9yNtCkxW4lAq94G1eLMnmc/sPPaRy4rFTvXT52w9H17
+0w06c9x8nqyCTawFYPLahibnvYRTsp9UalIk4ir5t8qmodf4eRa5Zjp0om0805Q
b/7bTX0MJc9598/1booqh7xeGGbc8tWjy/3B4VbKhWz874IqQGdCRcPP0a3+8AYa
uNbL8BGtcZ3C1tzlud7/YyeO5KWFi9UULUrORqiHK9bG+bzbTREUQdSicWhPIeW4
5ndDzQ8ICFj3j2EiyNqVlC/ULSfEcckdLxdrzSa8DYklxt5278W/Vqze6VhKUuD/
mI1NCVA2PC44NbOYq/ElsOsiHcQCsVhtsltEDpcQhFYE0X8sYDxHWj19Fbb0JakF
SFiGd8A+ipC9UKDXXPatuXrKLgtYGow2dwBcwXbdJHBi8XpT73Q1Phz0uw3IuKOf
EC9VHuk9Hqr1UtzuhUJWVxqIX2QN3gjS6bwGc4nBJDYctGzEoILfsa6U9qiQs0sw
QnRkkQrGzi6IBJtmgUPtO6IXQeXaQQQuSKUe9ajGPME4Ov1vRxMuuUFcbqjNwcHw
o9KH+Hht9j8u2mGQfR/666ssBMEoQ98JoESV2iPG9ERjBuaz98TtlJFqNHI/DHI+
VYI+vLqIf/8WJDsLOyY7CX92Ks+6I68qq58R4BBsQ/o7kz9ngaTseeuwEWN9Zwbf
YPkg1r8l52bHUvDL3SIxptNUkcoSMRDS9y90WbBUyyZvlPp71LEt7sOnaOz+cphv
gJ0zT70NC+iX4Fs3I3GNSI0qXcaZWciEslk/pDeBDXXsBEB6TDQrhiAkdtittaTt
uvJeJgVUlgkksp7y1VuDfSR5lqNmUpNJXWFkSIE+UN3aTeFFwQLUu0fq8/4HbFep
emNWuH/u5l1L75sT9VIbBWWzxzAU8BhZs0MetyPLXY+6q2hwpWzRa9OefhkC4tUt
R1W8/jsQgkmclPxN5OAJnEfoV2H3SrnzoeiQxIgGTCcgdiYPHO5AKjcmPVsjq0vp
H3hAWHmkPdIQgLSdh8KAzrK1eFCHZQc5EbeMBziPnLfSgAZtJoBqoDvOBtmPK8yn
K7SELa29vzUheH+dAGmieIHjXLv5WaznpMqALGmD++M2sRinQLZibLeqq4x3WENY
phYVAmF4xb+YJi723ebuzhY0zim9QrwF2R/XE2RoFqZE0K/D+L/bth6wmzxbXR1L
7phgNyA1mI5oALWD4+wXFlf4lPssX6utoFY5ztM3N4BeDCL+eYgjDQCRcKppnuAk
D1OmAQy1mlSL7mX/Lcvp5M5NszVva8hY6zgWje4SQMhkEDCKqu/x+nHH34aODUbm
Mxs5105CoJ4NjbdsIURmp0H0T0g5Zkw5nC4XhKXmzG46cwQan3tzNJc9wOmClMUD
eKrYLShv+GC8YAY9RGPr9aNP3S+uaiBLukqG2LBi0wc7A1SZWwClrHsyQd5diQif
N/6tN6y+bPvi535aHZTsk/3Dy1Nbi3XEHBzxtytKc5XAxearhoocoVFoniJU7gZP
JVQAzmSSdyqA+tV7Wh8xrF2OiL7KiNs9HNk4el2qkG7yjQM1WXpVEFjF2PpQEj4R
puzWAIlsTOUT1tvadQXXKQNBop1RJokiSpio8oyUShhgF7szwMKvnen1NeenLcCC
XAGeHLzaVC+phRzO3lLTnxr5yVOma8INhN8ymUnaWccmoe0zgolr3tbIPokMTldt
CBK+V32CJjSEAK6IFNoqtMMJGxBi89bs0B6BH0XtXqG3Gg7rITvSfQ2AAlpFRrQP
eA6fh4tKVzy44n8CHjAsZYsm1IpdZngtXZWYEl+yLv9u67Giu01/v2CdAsCiI/Jy
aFC+ZrzkRJ98IrXzOiiJnmk3MImsg6QztLp262BCkv3iXuoCUlnxr1VwhhHvVi7W
0td8HJI85mAfmX53AThxHvE9Dm7COcfha2ISXssm5v8ixP3eaJz2kj+/a7BdpVtK
2AsbxvWzDBNf4ksH+PwH5TRvFEo5F2WCA79cBsH20VnoY1sEi/Wf19Ni31KE850r
r1M9xptNhK4S6VzzS0bdP5xNDYoXa8A0B2S6+p+7KjCdYzpsL58sz11cCfRmkViw
Qzfgfo24A6cK79PgZM7axeVXeNaxKnIwXMKcYXPU9bcqRTbb7sWg7Byx2J4GPEk1
rBlkA98JAUWkpi/kAzDIuP7iLPjOhdOgZbwPEvQ0hthfkG8xoMiQSs/fX/7cgqmp
Fg+A++u7RgUjc56PIN/183N0pW4+Lt3UpSi2i/3jmFQbw+0/mXCkOY1OQYUHuo21
Q6neaVCtzbNgb+pDI64DGlN6UxPdPv5Mxa58WWvYDE4wZLgtvxvyy2DeY3qFV4QK
MKY67ej6suEvNTI/DU+D7/TRQ+o3ZhehxSFkf0JJ9Kb4Y6E2v9bJYsNLRnqv6CyC
X8rLQiKp+4s44Y4j0YLj3omRcuAqmur8+AUWgUaoF0lxI3nKQQLXng1vTsf1I9Es
LD+N/M3LWLO9hlSQGE+KRaKRQRDT2ylEn5x1B+rNGqZBIlypReERm4Xa+4JL6pRs
DeuXh4BBmW1rVsL6FiBDkStVkrvozAZTD6MDGT0pAFZL0nSlV4nv/+vN/JBPMU2f
i7CBgVm6B9WON2Hw/Xljrx7oUO8PqU7NlakIIHKE599Atrp8oqSQ4a/aodCSvtKO
lsCPAqDe74F14U+wsvRqSdhK8QKQvxEL+1osKFIoen37F0FHCaslgw4OK0Qo0NSQ
NuMVvQxgMPeT2oOg7f042icyCWfZgjAFp9DHumF8m/xs2FNld5HU1PIwm5wr1qZO
HcfSyQB6vua1Wal/feRa6uys51q9aDQGMiRrZl7w2oUa/0CzHv5ERlRNnkQyDdt4
6SLXzkdlnbjTMQS4/HoBiCtrwCo2/Pzc6OPc6pEcha64ZnX+CHsfZ24qTCI2HLLu
0HlE8GckkDv+A00k2CPXOhH50O7PKwei39puo7wObLkAdM5p8MhuftHdiHtT1qEA
T6UZQNNPmcIKn+qya53HHGFl0srtDXBOZMtivDXSqBAFTBHVeBQH5QE7H/7yaKeD
n6VL083kZ78XsxSWl06GreYay8hsmXDgU8Aatks95TMa7wjrwVcv4IK8G9AhV0mM
jqMo9QU0bMX0YTA7yY84Fo2M04H8m5QiaGMxwr9NW9+30Qzupy3joBcbsUxWebYJ
ZyG82+FlCR8PL9dWkY7rtdmAuAIr0y9f3NVXFf7LSJx2Z1tDSpmdkWxG7w0fIohL
s0uo7A9GOzjXDYcpNb9+O0YiCGDQnq2ETO2ei6R4WpzYu4VaFWPlgJ/0HB0z4g/u
qD5a115NdqzE6R7rjGl4O0MZ9KYTopxUn3ItPUSz1KBgpwqNPMLQLZaM2PkdpZP6
qLeNCJLQQIfQmCvisZig3fA1o1ebgCqrq5qbvTcCwk3/5TqOjcjoaCnbpo6EEwK9
KVEGilg0m4FqsydB1s8fRn8wO7vbpGWXvYilB4ToF/HZutB7DRQA7HG0o5nvQGTF
la8x29mVwCpcM/nB6V20mofuIjYkpKPaCDckdN1A4lmd+iIYzsSN8jLChF1uZAKf
LzD5ZL9/ufXxC44je0f+gvAktpncr3aAmE06kMUQrXDWgFk1Ve6I6NlGk9jTMdvq
tXN2VzpeX4lcYNcFKPrktLlTNi7zZXa364v+2DBgC28wgfKMWDdOiQe0uI5c2DZh
mJRfBHn86Iu8AstP82xGBddfT3jb3ta8F14uOFa3u/gjXhHAXCRohPYSrkx6w6Nu
gsc1PK6NcrZLrbC/yDhLKgl8ovtDIg4WeFBpuA0ewMUBNYGCgGYTp8Ak4M+hE5MY
TNJMlsJ4LsQ2NkGnhlCEO7/P9JPs8JkQwHCF3fB1T9PcfCFaC3nX9byaFB0bZrg8
MwUG2+3+7UZnHLdZviaTme7fHUgrLJTcw1kncU7dKeEqu7VXJPvUjYLr7d9BthuT
RNk0SfrsGikR8AhXmBaUG27FAQBjHZ1ajHeTZk4pS63wVb3yFDT6u2HvEqKs/We3
ntpWPFiSbGSthM16Rcc9jtrLg2dn77DJ06Og1ckELS7RX9KxQOWWZ51SrGJH5TNy
vl/cmuJg+A6Pw4WxXcMH+gMQfF6PSVO9YyV4ejecEy3UdI6JHg3L2wVMZpTOMc/r
H+3Je/0YflO7GXWYXMuoV9bR8lReVLahh0FIgQEGtbCNZD8atbTheL+EYvxxuwG/
wFmjBFAtj0hx8Bh0Cx34ONuHxdLu/lwBjdxo64/ebbvEIOIu7deXmLtgVRAl8/YN
SN1NorE+W+Axqh3ii0wQAOtW5U4EVpCRFEA87W3uUbnf1NOBFX1NkzxGv51NOMMT
lAbECkQsk2E4IeO09kDRAcxJ0otxi9dBUtdn76SSxlUNKuH5H/IZwoOP9JOWDFXU
qWoXxJPwZr+7wleGI6c3stltIV/SCVRX6mIisGRxCrAIdAEiF7hQ5ARinMpHoc5S
kuPdHQ8Yw1gmy+U1E/N9ePaYfmq3WNOavWMlpCD1HC757d+dYgfPT9MxsKit75YM
Ce+SGbbCHymy5wlA1fcCr35ZdVGrkMklQxFkbabi66/G98rerXUqzjvncLjlLKRe
Hu6l08sNVkLuJ5lWSdUwc9/ZIo7G9/m4AwzYd3ooADV1Bz2HNpYhfmlUIh0aiXuo
kABU0H3nN8EUyWHehgJfL88GwYKBds99PFvcWuXVWb3nIfs46qv4GbdrGyEIpYCb
kS2vqGqN9mitjdUrLbThfzubMT+3/CrAr+JVRgx0jZzxXRlSUWd87nlGtxhagcbh
4LCiMp+bsTp4xVgNzQ0Q3HBrl9sakzpKP+PIJ3DzQ2k8SXoHj7v30lShmXgf1UWm
xv4BpgVU4WocG98IVlJpoyVgqQ5MGcPXO6ukc/5fYrXuWSEJF9sMvG+0MBgSKGU3
xdBZBVrO6lTsf/Eq5QKDFTtxidNBzHzFrrFl1PMGHZGEhKKMXFpBZ0qyfxoEalbL
UYFDDHjRgLE63UV5Q3juw1cqu9cPmLQTXBGL5D76bxbWqon4h7kI7nE/7FQuuCFX
TLRdUArXwW9pT/WbmydhF4PdQ/1fYwHIY5flpkvfu8IT1ipDbPqs9kOuDTIbGBkM
b0Zj8mN7irSJ7fycdLopITU0d6TlTSCv1gNwYbdg/5zSBHlF4lme2dkdDzqrQmOl
3L5s9DQAud0RjZqNiMYAiunP68mv0gxOVpxAGddDA19PwMJaacE1w6GxTGvUVXU0
qhTC2EBtQsHjsqfNSZpS5bjli1YS+kBho/vaaars7cnjJ8u4iug/e2zB1BXicfs2
RYkzctroqE4k2zfP6vINiTTmMtZhIEueZb1XfhmhPqCJr4nA/A7RNLXKBH1ouvYY
xN1P3k7P7dmytVnFzA/BJ724xUnZMQLx+/opwiyA5b9RGfISdgv+Be70t/J8+r9y
+1IGJg3Hh3Mi0z8E1j2ko702OWzWG23/ronoWv/b0WiotnXHHLFWOaEuMA8Q2Guj
rcT1hXWKXbCBPj84xkzgSt6gzyaP+2qqYYzT3jX3DLZJJ1ogkfYqImfFPcULSkXA
hU3//GVgzDvTRONXCTjbnsIyPyDx5hP8omO8KrseGAGsLQznIksn2g4R3FrV86cI
BtCoG/GtVOmTJPvCmpA6Tm1FeWyPFf6lph8ocid2GeTk1ro/TkFok1nwEy5kemJQ
ceigSUCiTJdBAnnyB4KCRjO/znpy6lQ0gQYZxvKVyJYtJ3+msvKJOBaH8cBFSBrI
0kqegZfggkGBRHX5hf8Ujc8aM1MRm3OZqhXTbqovX68pC/LW5G/LtsfO0vGu74Rl
YQ4T7G11KIXW+O2fDB8wb0f3dEKkg8eVJlPX1+ezPMUmF3FSJ1ZTqPDVfnaB2JC/
7Ik2HS1DLR6iYt2Tjf5n3nJubZAiQcyYw2oV3E/udQ+kFCLJYF+6IQtsyl8ftFCU
aO8uyWhI111T1x/g3NA7uONdT66ncp8t47/Q5+4KnpaTzGB3+rYyjUu7BPxQBOaE
7veg2FmzXUxEkrdjcKWboGYUFbcVpEcgCiV9xrC6lTFug6+IZSScXhcGMI9ooYU+
m+E504AdqY9+WGFbYvsSa6/QWac5pJIyI1Xoh+6Yw+89GRoZ0eAaefsfEflIhIBK
9P4GFuUBryCmj2hE57yOkImWC+0SMUUrUzqH3sjxXuetu3tu/t/dvBtVAm76K3Wa
h5Yd/0z2ethYqhq6M9JFjUGcxCXZzKKycN4HE4XyIwiCqiljrY/ZjU1pwoN1lu4z
92UMjmaYMdMWPXPJgzz+tsiv7HV8MfT/KtQQS0c7ywbT1sXkaRnqqAagoW3I/fOG
NrtOeMirTarwa3fp0pzltb92WZ4g4PSa/tZdmzItJ5kRcx4I67UuEiObcoAZ5rCy
FUkSZPBgzt+/1jsguoEf+YdESaZdgIR/swxTFDKFAWqnpvMLaaZeXKyYqwQdpnGj
ZMPbiPaX6JwyRmnl44+AbJpbeZ2Qu3rAYWbVlKE5c9f5VDh1TJld6/vH1nx3zOYa
F6fu+/ixqkJ7++ZuL0Iq28UJ6bYgShFjK6tlf+VYwpXzgJrRhWpjJjsgqVx1pdp1
AJakf+HJDFOk8mWMW+vpHZgcGEO0ahZl1iWYLd8vFw8LdfppqXIKUwMxzW76Ju+L
1lwzjt6xE63CG0vTTpnDtlJ3DLATWIS+PREgUW2NsxfYisvVQWrbjZFUoFVzX8WE
JhVpPQOWIIRKQq15+m4ZZuqbLU23IXLfYcdNwm0YpYQja7pUJ4e5zxhwRIJZG8cl
1tQhJhn++DE2Yb+nL7CfIXHMUMHALFgIlnaePfg0l1l2Q2BotHl4gTQ/FXTtUDLw
d+gHyiXEj0zawmpyl0idsSwZo2k6+WvMppVtqxHs4n87RXbOPOXruFPNs/N1v++1
CM/xosDLBZ1S5S25A5mpEbsea78AmnfD2RuaJ3oSPsCjX4K7wR3GMcEJU+0ipKjO
HUDCMZ45wRuHaUO3SCeipp9I7FSxHl3CRtPJyAMLtDu7JZPJ4z9iwA1NnoifzAiw
KQinsIKod7dRJZC4glr3Xek5Y231a/PD/enNkSKODBb6X6mPEET3pYx030pks8L6
oWKa8prtn/HJ62n3YIOFg8ktr53s0dr50YQncX3WILsvnzc9JHBZvDhO+K0wKlfb
mXLdT6cnvEpZpoXa9up2wCLVcCcWa0tuBDNfM/8Jv5jDC3Gq8jlnGkeGE1Ol115B
DOqGvSwd/E74CHkjqtHtFDX9DrCmgNq3rfSvIN4xpYZMEs6nlhwVEI8nRHf4qYhh
trt7owU2NX3SiJValnO8iD/iz1op4EAB1U3X7sS2dPO2fFnOLnJilXpCywKG5HLl
F3ZI6cLG9eeSR5/cvvzGdsJPudlBF1JLbKTaaib464Tp+H0KTyPI/c2QYcCjTX4b
ayxjwVuqFk4nLeUkL/Gf4TGfZAuqmk2qIFRzuWrPMo+2jy3FdNl+UkR6f8U0zM9A
ilte4hMy/ngexAUEm5ExA938S3HXIrF3kR3H9glDaEQL+bQ7hJ2r8FkZz7gUBLmz
wNd0NBfaUIfxE+DetzJf+UtQZe6hsGJtTV1of9KFmbE+OnyR6vmWZLg8xOvgYYer
IcpbDqGpx7mciv6rMPVYLx6EV4LqPxsMSXlBGD0WObDmA5v6BfdB3S/eAuC+jfy6
FpcRqylcH1hRM2iLkb/q/fmDwUuiKyT68Bwmu5MsBKuwk9QnkRWhLw/Z6o3pTgOf
GN1SwTa4IUSqeUnc/bfxrdJBdR1DxkCRyPR2txTU6Pim3MGXbGPrInoLWVZb+ykd
W10jyeXl7TjYsYbIEC1sbcrPUpZBHfSKqVeYxKTrLSg7XS2Fsow6Y3R56SADHD13
Ua6J7jlIPVb7SAvlM0bEQmS6hAFAW4zI15MmEVkcvKcKdnTbE+Tcr0PMrzszcOov
G9Gr7ybN5VuYImZR3N7Hh54TIRXVeeV/7+eZLBns68YVHjMys9AR83BOH6xGSJiy
eEmfeOJtjmGwSVas0CckWmbwt2UqyUF6kpduMFgIVcjNP6HoqcZzdUCSjPIeQUL4
yayltrSiTLD6C2Bf08p9R7vhtNY8gDJHfdjsIn6M4VdnKOknWyzwT7hW+sdtqioI
UCOAWauxg0jWukGJj5GEM6LcB2eYPVzRmZ2cmK5CAcl7TyPV6bFpiWBAfHySyslG
bPVgNx+lsSMzERFWJoxv3u8hqOZzg4oZ3681ajofVmR9wFpaZYW6qoluR6br0Mp3
bSX2WXFpeAq98oh5nu16OrA/3Vh02mMy+68xs7QhcQnEzhmio5oOSSsaTLIUlGuI
+FbKemPDL2+z/na2c+oee3J+0gv7OGiiwAN0fRMBwyxaiGg0wiZnzeNAwEgiBcPa
OfsNrFznytTeDQXQCBqYUuOYqAGfMr2nzD6IXB2bE3CGitVVmdk6mnucl/a4ypAq
Jkh7UKb7aqF9QPB3SSWauYo8Aj+BXhHi7J9N7rk1syHugpFi0m5pitZ4/6F7EWpE
hjA55NGX7W76M1t0A+xas+CI2vm8p4a3WDFMHPfLUqOCz4OGl8AxAswskpbh3Q/A
+cMZWbzEeKbW86tU6zFo4W4IHm4+3N+cTulxWT13F6FRlO9qlJdoLCZH6myXWonl
iv8aLdVLplEbOVqVsFoHRn433IdbwrS8M57V6H2r8W9B+vLZWeW21Lk05rxx47XA
oywYdihp5fCLvV7gR0Z0GCVIpUTlEdC3b2mkItY8VZsI9cA6Pl6+En2qwc6XB2cT
jxQyQGpGMj9YojY3zMpwuAWjqgnxbZUF0F7sH3CbC/tYXMylFKEdL3SifjFgK3Uu
+dEyilULvXVAwHCvPy14LznxLaY9qUavWasvJWYFzturdBxxYqRc1e5RNUNNUQx8
7TYgOqhclqw+qI8KpNG4gfWkL0xUpusDDUXjr2ertV6OB2LUBN9znURMtGrK69Up
HJMjN7MaQx1+IkEfnwVx5I+sAH4148A+dmkir8Jcs3pHrgCyrzzWvI0O+tpPcJ1x
caJbPYp4mxKrFPuzp1XAVUqwHuMey0001JzkzKWs1u37jti3ipqqXaWPQlY1/7FC
wWx7fyD09z+ppLe8AJUD0aur1JFql+PXlwK3Q8B7cPWwmI2mSe7LmSf0RMvi7i79
ulToE5c6KJCiINiMOHRKA672lM4+Oz0DDETmeIRDlpDTDjzCfN7TRFqh0zaaQZ6n
8dnVhB4IAFDKFsCVCVN1ZIM7cXi3To6+cIrw7OmNFyQSZV3VJxnthtEAVufQ4xHd
CD/B99LdWSK8ubVcQIs29g4ed1C1p3x7XxXJrRIZCMW/HhkaN3X+/rjbbzUMl7BG
poANkFj6MCdkxLQ72Dh/tiAS+OvDf7salKpc6J4xTy1NeNbe+WLppvsp22JynCZQ
Uvkb+gJYnrZdYV9exA4ldC2BAt1TUlhS3pwoYWEas55EgrZ7cZa3OUDyL3sS8So9
GXQm40Iyxlyhyg6xOr8QcKPK9CuPEk6qM2FHYbMPWiLDd2CA4C7IuDW02zndlexn
/jcHMWtBp9gRhM0ra6Q80G6b6ZV2gQCpL4WOm87PdaCtX5lKp0U2/MbfiVc8AKTF
Wh3D25sJbiOddqPckgnHr3fnGOi7QpKE4gfizIjGOjGiGyn8/zydNTPD5RncnXqZ
ixkaTXkHFE2dbComkmv0p+XKJa+6cSsrFLK4nDO1Xv7YmWLqRvcdsrWpRBkj2hlI
l9a+3tb8tNnTNiCajHCuF3xhLH0T5FmY8nYhMFKz8T3gjVyEq7tbOdIeRGYV69kL
SVbYzmH0RAEUZievgICWZJZgjVS1cKAHyW/n5crk+5UX6k7LwPo8LtDBKWLKGmz8
pbWdfk0PW4laVCqXkA4sANLCSHiBykz7iqWrAtJ2BS4cIlY/PV9DAGxJfTJ5V0Uo
/CVce4E2vaj8mqwxfcr5QLFXZ9R5Mn45loXEGfJj6wzUxRAUBayexOMhQzZEX9YI
PE25PkLbxL0crlBC9uw3wFW3kjGAS6bS/E/6jbJ9z3h8+EmqLjSvZ/vX4AFyASF3
InbLzxvKCIvOitTuyD2fQKiQLJi99zcAwCR/aJ3Ti0VikacZgI96CAaQadhotf11
1OwAaA0hajA/0Ksr6m7S2/IbUCGV9sShbMdMLGsTgYfbUKK515r2mqaZf6nsOqtP
WxqlxeuiEuh5AiA1NKn7w2Wmr08on8Vm2qLBTdmhelJ5MaDN3efgAZ5L7tVIEPF2
3M7n8VR2wgb+QFKJJL5la8SAXdaDo5Ml65qmjXtQtOIaBLf5a1cmfHw6g1zQfPXm
/Cv7tSjY2tylT68mKsipUEo7gtfi0yrNm6vzJj7hnscgBBgTDVfnjHUSgrrxTPo1
r7IIZyS/7IvIz1QUID7eL9egVYL70KmafEw3X/iGWPUxcZzQc32iZjzjyRoKXx8S
V4b9Kk2Hkqymk5qKCLc9PGbleBMGWdJXqohLWoxdtLUcfPIorVZ5zVanso2E5m0/
b+6qLtC2fEZPSz4pw0GL4BaLpstrdl6ADscsXvYve973ZtUE2rPabfb7l87TO7nw
3+Hn7179IC9ejtCbxwSqouPQga7UVcbRo6Nn9RIBQ9gc6GhgPUKXDVBM90qkY5bw
trv2a9iMJLrQCtI4vODg3GX/QeTQTgN3IUQtHiu08H28LagxGbNHBmKaemopSrtO
rmSRPln6FDooAwTx044BDShIewILQpeIXmilomHo040UGv4Cw0EL3xc3TettS1/M
hM6UjrBSs10apSOEoyEs2YJI+rROEVjTJH+kHPIM/mj+GBwfPsmzc6qJc5Wu2U6g
pvbFvIaL7wywsLIpUApiNorgMTaOVDeo33Oj4LMO0tjb7ewxEjZQMlOrf+NS6dxP
HWfwCcqH3sKZvX+p5VAdAY4iwtotyYSo+kivFojscrEuS7i7s3eao/14u9NqVZAr
eIazF1FQyo7uo9Pk9y5CcrvbOuB7vkUohuKAvZFxeQA6Xw6hbS+VDtfEtdF1xLuh
HBCjAApKgW3EJtgC+lEuElMlTzsI8sTpzWb0VsNWfrgXGRmFFs0Z2LmQH6DEIBt4
TR7MvV0CkO290YFd/kP63FTdNn5WvVjKervw5/l/50wHqy4DkGKUa1hcKvA38rji
vs9JnDXV8p34GsVUw0Ab8bNcz0rpZgGxDUa3+cuugw3TCyrCgiTQV+rV4GRCmoTc
IDHtWWGYgMC67DFAkTcichNctPv8dUPME3EvkQiJy/ERnusopcIE992UfVzPrjh7
6FLg8clHzb/HmpnZiwxQFqh7UcReCA0Odgua9/mKdftovym6b2orSyhBkldOtW2y
nxQIqGg6JMD6vjGkgA7/LoGQTnh5m7VM+lK9i5YUs53nM0Iq3teBsCl79jvJg+oR
pRPwYVzKxCAdyThQLWRfpXFU4GYNsFfoU3noslHQpWSV9SJz9b6B/NzYfgL5kBfT
gegq65ZMlRRzhzXNolSNzm2gepidIrXY1pQR2uJNWSvBFsJHmKhWK8sIrSRuy0Vy
lUfvK/JX8YguZ49q4G7nuSrcRm/7/NVgvi+Y/ixjYg/h23lGAf7FakIZlhG9tvfQ
vVeC7PesoPY4OhWlLgZGQuMlaYcjSrd8FO4E54pbS0jzzxH7NiwPY2f85IrgmIGe
fAaKK18U8A/wTef69iBejdyGVQzK7ENEP9rzrdu0vEG8ZwJKsYiFNm1DFlAvUKqn
1+zyunbbu5bAxRwC6WXCWopulAQH0PdldE2so6/4aqvARdUTaIiEZ7feam0S3188
AaXLneTJo3uxWrkLGDZdeVNxREwOXp/MDHrIreDg2vdL8GozVotEcT7JMuWthnrq
qSURo7B7W7tqzeESbhrRFg1q0m8FGtSub5G8dplKe3DQof5eMUjLTEo1xsGS2Ksn
4aSPn2srfCVSAHzijtcUCwLB1cc7qfCS8f5wW3/Mib2eLiXmBT9TqUiGaJb+8hT3
K5FcZ26A+bTecOavOdRvEDOwILANIn95ZaCun6XGSeRbYNDyvBnClx4m21iOtE3t
7tiO+KfWfWY6dDDoIk8+4ZhHzLbT0KXLxtYYn1hNHOAvsR9jHiSCP3HYXwj+dXFl
7QpHek3RKES84ER7wxBMyZsodfC5TIt3aLq/eU3kXzvGw5rWvleEuP9XJlbiPGYU
W6FZCOrgFqnrqoYwZ/8Ug00lpYdo19nWBU2IWxzzTkyTIHQIuoret9qz4nvb8Cye
4ZE7zpxBkX8nJmcXh3380CHkzHz4izQRnNXBLQ3pkpgvexfN5NYTErNNTsAcOQHw
aO5xS0DgteHWYRGiVh0aGiOYrm4wrSVpAsBO6nlpi3/g6WDvyQLHhKqHV0VWPvEC
fhFOR6CQEeeDLVafLBaAfAoAeX5T2BE3bCtLWn23i1IGDDErVlejJxcNGhKjTVni
8wQ/UszKDSSvyHoXth6c7raquNVE64XE74nlc2eHLsu1AZQ8tt2wXZDsGC4Zb+Vy
iWOTTaaFK9GsPtYxZ4xBFX6YrBeBkLqysUIAKSM7fbE4eFXWMqO9fkvTNWjm0Ikp
dD045s6zctGmWnHCcfKVt6WRgYgEEMHtQUBjH1XOgiUecdyTiOUognRd55l/GN62
CDBeh1ocC0Hk3Kvdl1jRJ9nl447HTo0Gb7UzShWTk6NcEdf7Q8nkZBlCftBPHcm7
d7+B4/U4UU9/KfUhFHuesgnjy9fwWOFk8toyTz2P4XR2/O6dkF995s/BXqBSDvXg
LliKY3bpIiWWDah7UDanm65HvH/YJQmf4bkDLsOtJ6K5Rea8al0JZWZK0rmYAlm9
qVDjJ3EBDWPAnS8+sdLPbQg93QO3ygYhBsj57uUyiabTTxvkBj+YeIpUuBfooi5I
YDtS3ZHqTFvJZWsuCLG2q29nvM2wRiXZZFkESz/2jWHXjyDJ3HBNqOP6Emz/tYun
9RYnO0SaVupbKxCe5rOCg7lMQyn0F01/mEJoRoeK69bT1McGbYGKd/bHBCPeSzk5
Kh9dSsWBaIbY8iCrjqEwXEm+Y4FJ8Bcdm8vYt6rnTMYLlqT1aX11NQXuS3l5XIID
fu4+/W6lR4lbDy67zQkMiCbowgDvvkptaplD7Bz1eOSLMn6iwE7ooM/tro2c3Iqu
S4Ws8yeBw9/muRfgtM4ZWrk+LIxgwsvA1Q6k14vFCiHUaSlH1+kqfCmxC82FBllI
lT0JSHFQOx3VIHSbH1OILN9X4HmVLEvaqoUbkDZeLMFpysXlmzya36IwHAT7WXZq
BLxG0XRjR355Qim8QVS+ss1lQqFvTWzT51lE7CMqQMc4hSHyyCUr0bsLL4/XttiW
3MnTfBWAE34NiyMt+YeiiJQqy8bThqzzz6QITyMrPGSkYsNQpnnFUqUktC7LCFYD
WZUksbEZOaL/ZCB0v85QP6kXka+YcyQlfI0gREg8mvzHCk3hWWrhZPKkjdRkENsV
335wcHN+D+8RhFuKe7liweBNmr2Hw8JtZrnquE0uxl/LmKZmgNzSZ1l6ci2Hoa3l
jZz/BfzmJLlcoVbO+1cB9mlrjRIkVECs3cFDI1KojBf9ZqFXdy3CvInWyXvK/M1n
WD70netOf6i3G5grpV6iAwyOYTnv0BCRsQWFOkBSzRZXFhVDMw0q+AYOfTu35Cm6
NDR4yhwQ0ITqyB8muD88bVfMluWUETqC96iMKpK+S6MxjP8yopmRZeen68g/L1vV
he2tBQjLk8jcND70ZBvlvyjvnXx6xyKec7CY+exePvZFmeAdAHQq+gskEeSG7Djd
6+mOWYTRHKXt5GgaF2E348FQPKwptqfL8PevaxVYsfU2mAR/rnxZeYAJjvGJVTQT
8mGswpqwxqXYTQqIvSIMocqQ4UiVCBIzhW27fchp9JgNsWPPTRQDoYRVaorrmsGR
IcfkYkbtc9aMFGGT81bAcpY9j/0uVcoA1e7moGFgaUYcH+Rid0EM0vC5W+uw/5J1
EzzJ+4AX1gXdQzp4oGroBXVtJNVnvG6l/cluQtVnyBb1//aCtZlG55vZZDPEJFM5
MeqnkZ8bfRpzFxJmrKaii/3X4mexYSbz9UVi2okLO4dL4E6IRqD6YpILA5Z2dzLk
2VyEmB9AclLZvZYUvSUjj89wfeytEbqSn26aiDfRt+yDkesZNW0EQo0ycd5wDH6z
ImEkrYUTc8R+Uy/MP0Wyp4Osy8UvaDisj8+3KsN8NHTima9mXCHt1W45rf0Wj90G
h0yLZCIdKFGdYzmPg/cFF9adJZmRpVigkCliOVQbehuHnqsVastw8ByfSWeRnx7n
d2RxTWXJaSv+UO8fGo6uAMy8sDlGkRw8AIYSRZ9c+bT31L9S3s2sWdTapFjMysgk
i4PNIWwK5VUsj++JahcGe3SPY3O29Wtd6Cs6sr/ByoD/EFC2ptWyXbOeNBm3r9AL
QazvzXi/ccPji3ZQLTGKEzKHZkomWFmJTOXPTrFZcESmtt2ikqZr6SZNH/X5qqym
pW/RnM/2szIhOiCYqZKK2Rrk9xHitgsc3kBEpeah3t1cmIt2b+WqRPJ9DFQ96za+
OcQCsHElpUNlik50l+Iehm7CSzDtHaLKnsDiC1WTUPOsAKSxNfc+lX1dA4JuSfzQ
C+GkRhcmSmqYMdIFNoaCDorvpUacItYC4LUptziAUIV4iPBSGqOw5u+zFoUXHlut
uzg5mPfTbrkRYb/wmNGkBzKzjElpajnSiEA+9EC8J8mDlS2EdijmgjZEJbF6hKvV
5BU2tRzRVElEPN2TQFu2AzmSiwZpP2QHsMU97kZnZRBzTkra9si3oUM/xC5lxLN4
Z4eHDb90sG/uWkPwJI7TwAbsNYht9/aEQSd+H6UfCJJxcxFHUQDJhTy3f1kzv9aL
yl8khvHN/h8SIMgJHMUEzGnuv0NHekcBZelSoHbIXhZ845hIR8MfX/apNDNIYMfx
/ZCK+MGOoifSfs+BjYXBN7CIYy7U+pFt8qDJOOnyuBBegI0kn5DVAEoMel4h1Wfr
Su2cU7DyJgvOBsfJwgl9hlLueifgyx+e+biY9I7Cm0Br6++FrFJJSKd1VuYS+kPF
mHPYH9LtQT7Ec4vq+oM5tHQeZ2tdn1eL4pICqAEFghm1fsQyF8429i7TTbXeXLkW
ux0eDUmfLoDB+U061oDULVi2tpjvHH2halJRsyOEcCi0i9+M6dZwog15UGWsTsIe
ZMclWSiU2yoQ9Q04DN1bV2KmWDbsNq7Wv9ts/JjOtXA+IFTkJT+bbeBZe/usx5S2
uA6dxDcCqJs1f5crXz49bDEzJwt3Yc4Q0f0CMYhmWGX0NElJMsQjzIiwT3BgBvzS
bixCBpmcufviSZArT198fB71dZhW7ECiEQRI9ZaMOP+JlYFdkSBGNLZ5q0Fv8UVC
wvFgIHiGR0+dSTVr/sMSHx6pyX6gE0uKfR10NVvOfuDK+dHkJsEYbX8UgeThpFDd
wLFL/RyyJ8udkncrwHe8FgfAXQMeBAaMla5LTrUdhZqWELeFOh7SW++0CqLMofoJ
xG4sbdF9klOQgPNVcyoFPXBVR5BBsbjcBU5pV35kYuvCPi52fS/MI6VPnWcCVxxO
nhfzQe/23VoSUEdz+Zh2z9R6FIEhJGKfEui8ppgSu7tNrlCwytZWVlomyB+nOG/m
nRMRgHQkInFjW2tY1ygCAcMB9jKMeLMHN0e0FbQVicixLCi8GoJCOpMlS6F8Nlqq
wOYQj13FatfcysEZzC+YQVXreqjANAA9lz4+Oa/pVYN8JqsLReixz+CKt7mgUdN1
/Rp4Ab+ZcKGyQbJDeIWs9vnyHRCKCSTRlUng9EZj4jNq1Fsp1hxRQiqzdSeNaW7v
rmqFQnzU3uIqDNt60jI8ObmBXq2/4fx9Ds3apjdGZQjidrWMNfYyYysj6yyxXVRH
eD8NPjk8sIDz+3aoriOfIMDKPIyz7NhcRDzjpDn9yDlrtENDoNdjxQy2dy5U0AXB
BX9xz8BjSSfCESPkbvHwuO9eRnKp/8Ohyz2GNrC4yh5ruRnOTQoThbLNxRXW2z4t
34v06jvS5OAfRGbHskbCaHS1giY7FaTox4RxdQYpUGFIY3iQQ+0hBIho/cZFzYB4
xsduLAlNEVqskbPEl4HrXkNkF2KqaWnMM1iQjaNMzU4J0l2ugdRwSGA/7v5XjfRL
bKQ6gfESvUgPc7bGMNOTehZ5L8y9OKhWCMGAbQtgsv7dY4WOyspmvT0YQEDadNnb
tizE1oGdaKSvMXEra0ReY0vuXbZ7um4+YmSjBrAe0DygI2iaPxHzujLyG5khCSM7
5433iGcnSyX0pFHFPOBqoT/xMv0Tk+Ud9H9d9jkL7qPGjnSn4RjbOGvR2ziGlMr2
A6vfi/2OlGrhkP1xZZQJ3htTwf6rXuNjQmzC8jjNs8MNeghPlEFjFlmtdCnS8JUm
quOrwcJIfAB+3bjVphSPZrynUPE2dht4GLX76LNEfjiws39ioreVq8IioP+wVQ/X
6SllsreM+gGEOoLeTIJnCB0eVaHGJ+F4yl8F0fBDUH7iCSGSCbVly9pToA7Tarx+
5hTLjQMeddsHlJdD4F9UTSzNp1nApeag+XfU7B0/XQZvT657xVaUYjRNyvwShIVt
8PLAoctNj41gUPOIMQlV7n7j0YJhHdqKQVob49ikwVhARiqSt08zfRdjGE/DRzvj
nxG7A0HuJRtiUNCeV1r5pImTN40ILEk7jBYhoXuMDS5ZLtfXCLJUXFyW8UqP/QdX
jGwDIS0ylIleBEWpStXsAfuvjwlO/fvCU2X7OYIMISv1LS1vFs5r6ONvCikYIa1/
91XY2QTe476C5ksfvQiPgOxwNOgNWVJsgTudlFGZ2f7JrzJsiq2U1KecE61VdaLu
0HXFpvO9mS53vwR4APfnWK6HPNIkawP7OiR7epdJQVU3tmtQ2VKHLFQ/AyIyehSv
bnECsfkdkzqYfIsUfY3MKtpLYwvGU1sF71jp+CC4tHuBDzxwlAyGYshvvpHPGlFL
zP8JZxxxpPixcwmkT4cQiB+RGNJjYctMHMksafxarzY1eguf62ePkeL4yeqJRAzq
FlvHN0wyQ2svCY6K1v9IeqfRmY169vdBA87my4copF/9PsNGP6eRu9fnalhtRQKn
QsxomzMeoPqe8EaaL7we0wofrWaC2z9Ja2JlNZWiH+NRKJN1UhldGhIr6gDzpb+U
dR8syf4TsL1aka7d3tEq/kV4cO65eaQYZIt/rZY0vwzZGgb4QHI6T/O81KyzQbLO
H2XqRZ6Jp5dXmPi8bAbLF774wly7v0XFYCAxEHGbkEnWnGTiN74FvfAZXACMDJu+
7Gxn6w63nq+hPwpEj3eJYLNdsAJKT92lGzUCuGG5AUd8GUqinhZViKqr8PQHYnGi
bFzYLjYBui+zgurlCiz6v3V8li5nmSTT2pLU+Nl08/rzj/ReHHASIIfUcRSnP80M
QtLcm77n6IHOgOBgnN1wp3usoEmMldaajFcKqeQzJIcI4toWGBmoeJ0HLXxVihfC
a7p3nGEvPRHypjvB/+egKRQ7ZTxLTKCBuaPATmiwfmsDP0BpOS/ooJUJtheG50XO
h03F6B7w9uS5IFoixig1xlH8d4AbKFdIWJ0pTajh1T2jyUGyM84ZRsn3xobh1BcW
xwt5EogZ5nfV/vL7SxccwkAS/7nS8xbo71j+wxDrIWy4wTc5Ul7kuDEsBUclUben
rMTgDCqQOx8cnwXAHZsl3LsqxOFSd8a6OdfW17dxMBjoeu4FdvbNPaIKOLJ3wfA2
YEHzqyPvFCEnFmJC41FvYtNAoT9bURWnYVc76SWw1A1J+kv/3CGk5QY22pteQQjX
KiDaSXCBLp/SAuFCXXb6aZ6OQJJpuN0qzL+/Z1iKwIRxpc7zysOhdv6rhy6KupgI
nZZL5SI/oLEQrkooM2Zjfn/jv+50YOaB8sqUXRd2/K/azYbtCf6ceyyhmdF+fqvd
CKViDg4MOK9M1gxmtYJhutJYRCpVPLwXFUWpHmOLy2EhptlvgbKZFFNDmSHQJwyd
+fb3eDjViJl5HOxR8fY2Ux00ZFEa1mz8VsnqaUP9LzGPys84fhk4TTJRxJ9HbFem
86Tln+qTS+GJBIPtvwd76ToatAI+xYM9uK8XquRYhCUNwiujqs+JbBUXZu3XlZx3
edjqZ/W8ib0zfJH48QOJAM8/mNL1iGMdWA+qOdwBRL007bBDQk4fKRYG4IpGDVqf
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:31 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H2RGNRaiDKZ82du42bakRYvjS4uEGd3YI5yxA8F0IjS+4Ww3MPlWevwmfr+5iUy8
ISId3AxgtsVUg9b5Ne+2pgPoUKyyK7mbvSlmVfbGFtWCTZeVrWalDfN05tARZITe
pC6o/Y28xArHRDT5zYW8pF4AY9opOOFZoXh6cIi9TbI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25104)
RT0yb7tVXO+YWlRUv82ADfeISUHRjUAMWmOV9JjroS5Sy8jNFEGIRkoi9weBmgTo
7OvRRzn1zTV0MMyrkS/uyZjgPfBvp3luvWUc+tQ7uCWMUk47mVfvlhfQSFZbYy6V
+I0YuBIWLtyXTQO7sz54QYLlU1l/xX6/SlbmIQ9cT3taQ82n4A41Kdsz7INi5w9D
ZGh1ohjNoCGOhFAIsx5pgjkwUofQEsZwN8YQLrMue5tkAkj4S3P+CVJ0xVvGagRj
lTXO1FAzsVLqOEpB0ykMLNbnmaFVE0p8FEfaeV0xaj5qmW2MlMJrKf4a9EHbPBMQ
zoNuvSHLBVNICE9trd918NVoQ+Kl4cCBdXsWUbdccquAjx6LsiqVGRWdnuKmhYxM
AJwS63TVU7Cr4MEgvnKLsuuQsRxHT8rMe3PdDU5ne9XDRiye0rgBm6ZINb/IY3LV
1w60On1fTDA53zy4ecsAiJizF//ZiVYEktmB4bGHJP9YXJ1axhIDsyJSHkTlhwyU
8Ix4+BV8kZEiZWvF50uDalXiFm8xDwzaFg/+j3armlYCMnT643I2+kMCWZURvMx7
UbxJ7vIEp82Bh3sdzrItREKujXnoHHftWjG0mb7ZxVLiuLbOI1F/BGkCk5uIzq7J
IloYsL2+xcaBQZOlt4UZ0JZw6BXl11hIPxZ86SJPpM2sU1Lm2OEk84y9N+dmpHha
Q0cKGtR2lpkF6EUToz51uVPg3rRdolF5cRjsjCDwTBE2ntdHWeZx+euqATK4a8ty
UdGs8ORuB3ptrs1koTMni7Kw/9HyKHnSCC4lcfkp/JM5UNSiaaPNATFNuZl6iW5B
thcjB3NP6Q5eXYRHFuMZbRQKQRUqtPOPnpuCuMgsANR3s9B2CJCjhVrufm7+q8Aj
9aN629cBdU+e/Wb6HItueETQ3Ak+Nm4Ygzq7jnNCh4tV5aa3y6sfGuaNAVhWr2qP
q87RfPNiu6vXNxfek1EewoqV/S3YedqP/bO2BxNjSCV46mOJpe+a2H9UyPcZwp3l
sOo1FWinfhO4QCZy6MPPWwJBNsyTGZRkh/huWq8s8ha4EKYdlUs+UkOn2wizqkK4
3fttfeajVkCmWjsj37Kve34xyXc4uszALV2jm/Pi/EYTCELwMOzTXV7Hm6lYE7vH
aj6ph1G93AhLTqu9JWT6DMZIbpbKwjolvlpdmyiGi/htcSJfyS9RP7bbTfbAOgof
1/XEFvZDIA5o9ESCGD58MJnKULPEu7YvdEXhARozY9n3R+pSJDkHccXk5/FV1tUK
2/caUCCOTn6HqJi0nhSaHvVXQhsdpVbt4DhqDvIzy8AjrOB+kTrjwYhQTmxtWvi0
uQPIWjKEHavSab6K/eEu3+v6UtwiKw5hnY62IxMzRIrd1qkRMBRrt/oFSqusw3Qp
DXYleYajoM4kGmIXhULvb+g0YzOsQDDpLanm+crnHXYx8wMlYRHYaDYHaA+119Ht
y67Zcx6kCkaJpUUd38E63eLIMaGoaMXPvadCiCxbvtruQ4PTY94AoFCvUxeFAd9D
DAIpc+fzdExkQoQepwdKmNRWBgFcLf97J2wxLgUzNUpkSNHOUMn0Kuwi4YXh5ftg
FEshafhskfW47WO+Tz60RxdyAh7+jJAxy6B6PeShrwPmSy7+RsELP2qcRlynFbCy
GBHG9/BmMhVr1TGAoI6xkuA3XYFtCAIj2l94umBmYMuiLNWt0jikDEPGw2b+me2D
T9m4LjD333cs6i++aSz2XoZCEU6Yd4DSIYrt2WFXW1qSHsMR+4YowcQWe+v1K2Ky
nKajeqqLEFeUvipfLMrrvt8DAe7cI7z7SQ4APjTFjzmxREUbTSGLKQjPaA/WisI8
AxVOGqs5wWxf4t3ygtIxKhVMy08c7dlLO4TcaKZBJD8Om+BWwEN40AGbi0FoQnlh
f64PsnUsTzYEgOsm0s9pozVARmOFtfEXkl45hkLZ6yq2J6e5bkOrN8GZ6xQK1MtO
cvZEbb+5vMwCKZPI37T23iLLpR3xpGyRkm/j8O7APORk2MkZornEbq8Xb4bctMgH
iGqeBuUR9nfMpGmNNUug5KhuPZIAfbqQhVgiaVsfL2rWgaLPw/iQmrRVs1qjeXVH
5Wh55XR+rCjkL6aL6MVZ4ZT2giM/7G9Qwb7n4GkUTarAh/O6RxSMh0XcVmv0cPZs
KoPbpjTUXncGU8a4H/UbynmhcqwGheoS7zKLc9zSFDPyz7rD3RU4jib8pH7HnrEr
CbbbBIdHxHrYfuJ1G8X5QiD+0ThBAbhAOpBpJKqBrbEi/R+Ap4NyyQZEIPIVmerR
tlN1ZxeaVr/Vtf0YD1DcdoCPthTlzjNruSdnPxycUbYUWKqrt3d/0zD9NzjBxpKZ
TYiPGPs/mBYM99DYRMW2s8j26DnX3OKZHtluZc6BIvtw+kW2iXZAkC7RtDXK4nH6
0mJ2MThRWPFXy8mLNXqaWA/DgydkyXEx8rjNmZR7ee3uQRvCkEY/BO9hOFp9XmT+
deeMvKnwqI7sQKeAl5qOvPIMBEt1NGX1iXDzTF+NVUrgjeY1t7IEUkbEPGtX759g
On8lcsySETVPvrptIIEO02IThujGgeotBQQdXd0HuzVWQWPdHDUZ+kay2c2E+20J
ApFQmXgAhRxGMH7lY7Oj05O6kw7BIigseR0kGQoMQuEHHOyamL34iaj0Z4gAUvmA
7qIaTjeuxF37DaIA0BZJtR17hayGtDWtUKWhqk4BWh8jkgRSRj/Xsg1M8qZGm1Ia
EwriKQ5Xx0YFoBdlXjW+aQRix8for/TOTxYpOIFE7DZymkEFDjk4tt9MlwBiBw7q
vfquBpU99K7nnKNLNG3oMOcNyrL4zr7WQtSQwbQmMN6OWYiPVlBoU6lNrREyQ7va
1ToftEhJxCOs0Xd2DekmkitNMQqj7Awzqir0m2HphzLbFlcne4Ug+bm9t90wG4wO
lQrpkO1OlbdU3fFKxVjVgGQmN2bXxsQPx1/vqbQAepyM836ep5JWJ6I5zEw6vyGl
Mj99gGGjvSU5t57N8R2jMa4W69WI7dbujPnPxDbTJcjPe6svthkSuFpC1ph7e2fN
FgEgFSjMjPwHHqg+sXQ0CAzCiEmoSHdsqXo6nMie82iM/XU6IW6UIGfz6RNqXxMm
JPsarzE+Kje8NWTKeYaR66G7vy9obtG25/0J8TEUV4z3JJL/incttXAwv4PV424b
2uPPUVOwu5pi8T7Uar/73zmflPhxvMASmvoedXOrgN2r8cvYBxym/YRwnXU99Jnm
JiKO1NXBEY0+7S/Uz67tHPXmOy0ACnP8Uel49i47Cu/evNOSbto0bX+PuZoJ21k+
5cC4M4zpPOuTLWfWqCJVd4F9FJxSec/ROOYpW24bUB+OAd1VcKgmn142o8ouYYcK
+95bfk/jZvc6w/AW2TwOKZnG/nhj33f8TMFHfu7UF35DpguzGQlON07dryLB+ad+
OCJadfPTBTY8YqgkV5v/gEFIN53OKy7Dbs64EGJ0gY68xiKr605+oeGm0/fG4LBm
XwebY0qApMK5Cq+iONhM9u1dirRGZMv553JlO4ClK1Ji5rKILhw9X7+qiulB+rFc
dUSh7kDuXGqiX0PKXHWMVs/HmTeBcYrR59J/NME0D9PdsCV7J5dv5919TvVvzGex
8e5b0GDmv6FwssIft0L9gn95oQJyGQKkIUy+TVOjmGixKSQACcH8nVJhXvD/HP1y
PauzQE7FFmY7YXNabNynFq0pW0amEbTsEgbsU4aTw4K5wpGVIuUBllYhFzp8Xv58
hfUU813I6DxmQZ2GDYq+L+jCrz/VeJGyyUW7gv4mF7euv6eaZcXq4Jk0NrCiGrGn
kgEA9IwyGt0BapmMqyBb0Iij7oebcKSv46j6Byn+/uUttpeA8gXfiY+d8LcFJ5ZP
5YQFCATSJLhqWkpiZYJUjKBAkyyCiVXXgp2gNHLXaqkQ5KLTA5EQMD5sAmDy3h/q
A3+z1pb7LxdtUkYGVrZ3nVSrOOzQWSSFhztF3i/eTPGruh0r4VqAoZSxQ8lT1Pxr
JDkKIIbtyMv47fiM4PRE8R9WRjlqVFx2iz93huhpwVTx2jTd4aBoPyu+xHJl5KlT
GlVPCiTSWuSEBqpECIH8zbV6TE0gkUo1yjRO5vU8/gwk/kRqjcCWzxxgVqFxB/Ng
Wxr+KlR1BX3WIV7I93ym6XIPrmdbufoN7QnGic6ce3zzgZ99Wclt5rZ8sE8yLYLX
1PwGjxWP5+Abbeh/c6P3vR/LxtiDux0Xr3Klww7Mr3oortrZXlu6RYsbsLla/x5s
cygcKcKAklt7qnC7e4vukt9Z7WIkQEWABSz8sc/BauG8DJSzijN9ROwkEN0lMsI+
D8TflrxKw0ljFd5Oex15jadWpDMHdQQlwnh5os/3a4SEyXRu0ol+upNGXpiGT80Q
5y+VZxwgcI70tucvtHxtOLtNqkLGdHlgMnHI86cp3rouSvO0sKtTRCbmcaY9XEFR
I4CJxZADBu5p49zvlvGXJMhz/7Y0Z3NEzdcyrXliLSECzyUH1oO+R23xkrxDil/A
21AwEip319m4Mf+EVofIO0zyZMZIci0cTZc8yuDXGV/coPQHedHkciYp6BL0ytSm
qLz/oXBFlgZVoKUIbiQxDIVGrvoXHzd9jhdQ2Ef79SLgjzKf5QneJtO1qZDoawQH
uBVkuw6xjyxfrFKCI68gd4645mqFwX869tRAsoGLc9n6diwFYqXkiiPLVWqQgCHC
HGI3tA/8PlwgGq+jtn83PBAxT9GVnFLOtavfLz+d9jVGUgBZHgBtTfjupV02vN42
DFDXptb7PJM3iCnq7TuFlI1NPV/9vpwXtE968HM5zGQxyu+N5AbN9xuhzp0XdEqC
6zqGl70NVHZGIjY1rpJqu3ZGz4lHeDIPlXe7umLekJ/dv0wjr+3lMwSwyBefRqZH
h8nuTdmnexQiJRzTHmHM+/5R21vg74O0LP5s2Jfxm3kgVSKiq0zpqrvOFDRuVSK5
NcfxHDRrApIwJfv+Rc3T1qGkxP2Y1Xp92DVnBGTw5QekF2lTFiAFD3UU93AjXSlM
vZog0d7X1Dwoff570ONvWkMp++xT/40gmFaVyjvtXLfVx+sptrdkCb1FJPNIRDyv
aMj5o7MS41H6sxAlMHAXFgic8qP0w+GLeUfU98qC4HAmjV+Y3Z2ycuE+hr42/tBW
pAiDY1Cyg5sMNgwRk16XM4/PUo+bPop67PWb0hveyxpr0gHxDo8Chw+wdyHzKXzb
WNBiQvVTgh+9uRXhHZV8nIVVnfetmE+CW4MUmSdwBC53WPb8M349lavrYEaxaNdv
CoTmDTOFKzfccsvBFhSWiu9GmgGYe5vizbg5dXCouzpbP+h7ITBke1sByID+Ixv5
+LGLBCvlzGyjYMIE/PxJSz5pVEUWgMce9IffB1pbiBS3luMUTe9V/lyJOC7NQsT2
NW2m7c9EXep39LYqpsvGIVftEp5QBORY/a2wsxofdyKORDita5EiHO+XYVW6CnBx
NrOz3h3M3tLJ1fIu4EyjLxR7wosOlT4VHYLAtFsqHtO3Mn3P/ASUkcsOKb1foQuW
yMPIDUMJ4+eHow9TzRXYOwg4Rkwm+3TWAOYCVW3iq3qRITPZPfbCOHLkag7YUEfe
p1nrVM6jY78VE8cpc9pQECOAITe3RaQxM/xWqBvJVPDmRWSD9fqsOHFJpO4V1s8x
5ZV/nBPCfJgqRB2qG+BuIBRh8NPPFDQjhk7dcAdKKW9p4Chpn43ZUJDCJl3Sr6op
9ojGPYUFUsQ1+mSSWoXMWEKsCp/pAFCI478qDyRaOmzjfse2iRUd8lvxChQ2yraZ
fRQa1SwosgculSwnaIYK2g5gt8z5zarfafZSAGS68YQ1oWzPuxRaYcjBSo/NUhN1
TEN9tyn/q81yubDIIseNhsMiYOEkoQNNd5TonrIKB3PL6TALTK1hG/kkVcpuw4HL
N3XEkwrwQ7jVF3esLd0CqUT5JPeXnQ0LVLEI4e7osMSHnl/XgIcVW2VS09bQrFMy
T3GP5IOxVcMl5sHlzsTRX/6pxaeKA4In7Q4vJ3R2/A3zGd4tP31gVdNd23KVsSLq
FiUtBC6t1HPjwRGZkxD20mS57oPx66g3NIQ88PYtR9+6frKhBo5CV7dcvsJmGBAx
dQDxO4I4O2vLeoix5KG3J9Sfp78JUYAnod3s5h62Is7HWJCnPe1ZDLptqnGAlMVo
mRutYf4F9hx7Q93HKl5Fd/lIuUSSOqKT6ImOkCsEZH1cJAJRXiQwR480+tW8wrbg
HcCMQXh0XKXLwgpHDjc+ABDcXauxVXGcVRwIQklA10yLIsSw7vLTSoVQiMI2y42W
zEREoSxH9O3cVaT4ac69nx95r5ZSao+7SzLPH2koI4hYkHOdtCnKTtHa+ox6eJ3W
ohmSoUhu0GmD7XZmCheZ9MJFCiqwDIZBX3Glun5GwaTTxAwg0tLfX7phfR5GZ5wP
FYr4UNtriHljfVJN6aQ8Z+vYMG40XBPFQw5xnVLXuSSPNQSi9hlesKyVKOkbZ7qD
6/CzkQ4SfsNKr9FZAC858igPTWWc2Tn1KRvUFR32MTmEjoiGJKfoEVfjRfFEGL9H
mVlPhXq3AUT3TKxNCZnaHzvMJxkIA+oLyvlV+1HXdmpW7VcWSAe7mfP7DmnkwKKo
4g+YBtMKk6AcZTzUxBD7OgPxL8inBmhZYR4rqz4ukqBna9uvqlwMJe6HKXnedUGj
DhXPj99E8W322xyqp1B7JOjdAT3Drw02wmBGlBmvs58t/u+tdNQ6pRnFP+IEwBht
FGJmPxAFA4FAvwlGpF37gLYr8u3TpjwhSWt418lJlIVRO2j8apVA9nMTXelfSclX
8Bmy/v7b7A/RNOmr4WMHxfIPuwg5ZX6WZV5NVWrNdY/b2P+pt7wJ9cDw0/TydHui
neH6emWH6mhHp8uJKlafkruxiMhC7Dg92cmX40E7Ml4El6x4PKtASPPFFGOpab2p
PNCBtIyN7Dt7Qty4MlSpIvjqT7L8fj2Ztlwf9lKvy2tac77siEfquO/Ih9R5boBS
031UJMW+72fMY8J9ab86I+kOEuA7zB+eWk7kFyGTfxpJDbqUKTbMXbcGIyxmbW6y
NdvWdAd4A3bBMBhVQAhrY+BS/ubIlYuc2hi7mWJgIyRS0gaIeQKeQ7f30sKvr1rh
V5XTd4k72Hs5qa6VjTGjVJJDfiqFC8Usr+mWbkw+Z43CiKcJ1iCLFoQ673h1mwcl
zdkDHZ/EvKny0thJ/uITMXwGoEUF4QgggG5N2H9JeLqjX4xR0ylp61M/bH5kyJHz
ZKkz89VoM8mDJT0NpEFKwHLp0lGJBCNl+DEO/mLopmnFo5LF8QlqvhYbOI9pfv3P
GtzUV6dCk1ijtWiGDwWs9qnlFycK2q62Fv97w1Jd7UDiDn3pXCxMhej2EVj90SBG
Mv6yGQvKt8coP2OyfCJUJyJUnROAakDfgCCO0Dt+TziTWY+rnjm1g8YoLZf1vm2z
dl/R1XkYfIIHT66k/rozzvGrSDe3YZTqYbAstAJWKj+8N25YKqqlnGW7WTRoxYAy
5YJbe0+IGRcpfmyS3fxlChcqdANmY5fzcW4+CEQ1zv3n3hauZVCHHX+eMhANplJi
HOQbz9Im4NgxJ0k5/MSZy40T+gk3T8rsU4iWtpM+YffTmhkAHFsGuPaPfp/eFwYq
RcGRZfv5bafW8BcGtMfvcJWE8zliaFcwyEFrJr5Ruu3ggc8TbjO87xNkB+RCXp1X
OTdX5RhKtcmMjv1R3UuBvUPTPAOQldVXGHW2nKj3bxcBJ4cDCWBMeTNAciC8wn49
YHqQxTCkCoqQyk/9lXI3p5ijWEWG44+fHdxd1ve7th9K4GDMUSQR5FHK/BhU8wqu
DaAAS2pTNgSNH9X0J/AaC4m/YvUdWbhhqMykCjumbAO9ZWEn8mtuIehaZfGsboEE
4eSghXkelCj0PlA/knt4MH76D0CKqgJDSybrhPWX66gVrzY+fC3Ulmhex7RnNf/z
1SQU2oZVn8LbJgRYco2Ss5PU/o1K9kpWkVj7VANIy5WPoHPdVe1jVhJnSrBknpZK
gyX1nY6hzn/VFC8Q2OFyocKxnYArUop6Oj/MCeWeYH+rScfTX4zn4ydGFWB4g8EI
/BOWfVl8kKEZibMpilTe3xyUU54+4LWF5QqkmMw8SmCifHZvItUG+2uS7nrVsI8H
l4vYymKAmHGwSidHJJlYNj1AtkXhYQ8LQAtQOTTTonQ2/rsDmcBRsXFVEn+ZN2ui
pcva2iwhrP8/YEwfIS75uBSnt1a6xYT8E4icufTBA9g+ojX2Iwq16krhTtRkmlJy
ZUOvhj4Cu1tk+DiynFYGhM+gsHHavmJvyBTel8fdh3JKCzEf4u7zXhHJxnZbKR9o
mQffRroydCep/gk+RgVnNLiAeuaBM4jeZdYkeu0yDx9FlAXkjszRofLvoRVvYbdb
7SGvZYHSTM1of5TBXNtgscjzInSGnpyYBDxyaMj2yNsO6F41gKdwB5rAaanFhPDh
CJV8UBbV7AV107lYkacBMbckqeD9THbJmCxBffN9G5rNeRALNdEiORBOjMtyh90U
3OOkSDDP7QvU5Zcuam7GZRjg8kXKj5PU0wf3KQahlXkWpoL1rnGYFRNNBbhmcrpd
6K2bV2GovqatwInHCDKIaZJ+fvjb33H4BcVd5NsJKRmkPZNtGeLv1BfuSMKnbkED
7zXbBoF/noCPKYYsCUYkpK4tbv2Nz2OZJuHbbQIgSW+aYZ0nQ6EBkPpS05aQ5GHg
4Q/Cm7qZ10vQvnK14UwXVQtfh5jZnkow4EHmC82A/m5fgYFAeuM0rcFVqhAEO+vc
34DVLbxLH917ffapu2sH5ar3PywcT3wZaMF9JCCvFgKQJbaQafrRg0HCtERvfM4a
V5UtzawVKsue3QZEQp3uZEDeuMNYp0a0QozxHnh7ngrTEgs4RMuOeNJv3CBxx7TZ
eKGm9lmr4j+iMWWjtq4jJnG2qxBe0l0Ez0QBVF3ikkCWGXw1IJNmXIwMVYu15une
FcwrFTpWxvts8+sLN4TsmxuuMIQlXfYdJVbfwf8q6Cu8rVCuHkGq+w7hzcVdSxjY
p51lnzk9WmQywPYL2ZE1z7dNEq/d+3nZ8RwolvvYLEsbfEofD297Y2bKODDEO7mF
NQe9RLmu7w7wfQy5Z3nniRVv8k9qIy749Ipy/2oamuU4V7GbwMFOUvQdeij3HF5a
wXVeWlKpr0Z65PjhsrOqI2/1/HXlWNOVUPA2Ez7vkZPq+oaFW8Dv8UHJCLTrj7TR
MPsoQfAL5ueRygqnLtqvQPXpRMpXU+jTtscPyNP7J2EbGVR+n1orPHbDGochJCq5
K0tgfjS56o9QIa0ge3rqAL4RHjmBjF65TYb4m8p3sidHnbxllaZEULGiDrpCWQ8z
roL7DZ/GRFU2OJsLrg/1EUDLb4R1fZOrQbyXTl+cdLCsCfPEqEVZgrTKR5pOwzhx
qix2Ws5xJF1opPglH89j1Hw/XVIIuawEfj9gl86rmvSO5usjAUhEcdXgIL4+tUp6
/CKPakZU20CSAL5eAEROg86Ceklh7+Ie7eI40AhaXK7rwMWWC38kcPpGdSf4uq56
hpI4+snhseoOmmy7m89gcLQg1S57oyF4HcGVSUU21hV+LzVvFG843Fhh7ljSqhZ4
f/kTmLn2dgpomfUVk2tgmlLzlXnb6eIwVIqkc6dMbWB9exgF7kwsmiSp0Dz00UV7
QKR8E+gTWCCzPD0NQHtrcVOng2AD0hL9UxSCl0yaZAy2kE6BW3tGLp35zivZ9nJM
hPu2GCHnFY0K/r7C8kCq8fmIH+VJwhIdZFk9zierY51rRiy8QiP8MdmO75x2ad+B
4EY5zxM+xKqN86cBQMSoFuzmi6oabFRUg1ToGuEcmoa6sQ47p5Il1PtH1gCSjBfn
n3CzjesNVOwKrBUZNkZKUxGoNft7oCF6MsIG3ch9lSpa+SB+5ixaMOBBJbpedAeK
4aHebzRR9qj28YYTzFEeYqUYOT8yCBKPmim39WsFBF1VIzj2hd3SPGvX3MYa3PfW
xybZAAbNr/C6ukFnD3x3Ax9cUdKg/UC0PttN5vsZXdTEJagC90BX0Z9ax47g9gz7
XHj7b2KNLSoYsQBLHmkbfLLEeIN5HDc/+ey6W0WbUGujOvNDlVl2SZJNz8Mg4v6D
z8ZnBtYHIWmuVmpePZcSGSpw6eeiSSL0COJRZFEdwQKEB0lDp4GxOEa8Ao2MpW70
AkMepCnY+CXHkmX35i0rccH2B0mOWLRA0IchpZiiKW2FvWQyQehcwMbKYjZ8SyW0
ihsyZuo9V4vv4snOgMEwFmXD5FLOY64dBP3uM04/ef+Jh8reuY88frSl2Zy0tYjz
UihWQIcvXytwZ0/Dfb4HMNLvCB9hRg6fp5Fs5MnF89KMy8aVvMj9FLGib3X04Afs
xG9tJij0Zoee/mObuEfcYG5s1qdiyO+i8tbt6Kt44Gl58KWslc1xiBmrf26xFP11
1t0tuU1xCB8VY72rPrIbZQnbhT3r28iZ625fFlXqGFrX8RVWfxsqwKX9yR1M0nFU
T8PPN4TETjxsp4u3pBiIT8NrxVjp6IzAbISKMY8V3iL7mEa8ubBpzN0jzdlmXlN+
uhCiMgco7YJTRYLiax3GfOfbwD+lZ6R9YGINNbPBECQUWVV7Ys5gpCH/ahOJ9lhp
jOf2f5vsIkH7UHk78QWEH/kTWxLyz4k3roNGwwkRStEvUuRrTp2H/y0SgGeqjkxT
Yc0iwf1GRETE0EvZGuApicC+DyUcj41/LIrzHXqn0LjF9eyJweMxBvDeJujAXF1f
cTi4n+DK5XBCvwAOGkVgrFd/2whUSILQBBgZtyWmkAFx+BVTsgtIExIfRYKgLX5Y
xTG9yNwIarL7FXViHhuYexJlS4h+Hj4gdjLQWMs2ZapMftl9R3aLjSGEG8RgZauQ
ngOtVJfOK2qh+n67+bxYUR12P9n3BOb5NcmIwTqWoyywtOrxMetfgzNgNqC0QFEN
Pn5lvSr0pxZKtP2sb/62zGEw+GG0PxrB9YxNIFtWVrYj+vSL0OhoLv6k7RKdNjKP
H+b58KMTZ0QZ0KeE+MyAGOefYwFS6PpGg+EdZRri/P15HIVfcc4p3Q7EbYSephrP
HhBuVNw5AslrlGmjJa2EXAHnrLBscKFkFsRKP3QaKfDjmWbNV/tSDXhafHT858Mz
9xI6VczCPg8xp0/twFCNnumOtlVs+BA9K2Q8RB1KV0yGP/he4AQzKAnkwp9FTz9/
S6ION0b9cS4nZfu6H+j0eCGc2kcXT9gnY/IuhmHSSRpUH/V1Ow1XaudVv7SLDull
weBc5UXEHgOL9usrftiCgo88XRlKOb1ueUkBAaS/LeQW+IW65BWLMPn5rB2NrGUt
8WwLd/ZjyjgrO38uM0PicCEyfwNnzopW/e4mDS25RkVwRWDd3qLNCl0recNQp/mw
Hm4NctW6kKiwViJeJMlerE3dJ/XIYoiPfqqZC4RGsFWtZ4ZzvjOSxBwvQtmLSN4x
4nfD4ZcdvnqirQK419ca+OSrrrMAtoM5Z1iW4PppUYAUV0MBzavxqRzO4hEPKbOl
YC4jnYwb6aILRabYd897kviChSV++6RdYRVYq1m0dsGrr2MNhtHVWUU0gq29Mz8Q
wnhl3jKQmwVH/3pPLzziEv364+aDvOhQQOxq5zhzQ+cv26fNcuaWynADqK+KyWbr
xyFrCEH8VZs+9hWzGMNVwNKNY5MQ2nTw6rUAM0avvnl0HWlf98cHLlOGojIjGpnD
jhs+kGUpE41zo4PSGsry4c9qRZ+mJsczInkin12UfOWH2x7De4BT3O5bm8gprqzM
kOPRqT93eNPhGpZ0OsNcHpfAywnmhDDf2awkoth11Eg4z6Dw9QawFcoyhOIY/Q2r
md+4NPfdsFwItz7hb/oksPKxMKTrqNv1yKXzez9bQImeznjjJ4hVxL0Qj3MeubOM
UL6FKVsvT707uO57fERM3raN4ZFBJJ+/64bVE+q6AFA460xNbef7DKj2g2xQ1Q2R
nyRaqcye0BzBWbtERTDqgltTnls8RUHnRfJ/RJlXjGyR8bdBeYRPw4qCpDs2qUzi
5JkVVai9ecnszJM4VqOS1a/z5d8PW6Wkr8tWN2dCg8D3+Yf6BCSL25V+/M9l5SqP
nqqkwVXk4Lr1CYmhFaodSXgI4ZzR4VGW3uMtL8MpVu50AmJNKL6M4EITlQM08hxN
K5PxO48VRivwzxCGIHbtQwbt5oJuh/3QcFZFRSzABIps8AHghD7Wig4qSWwCFF/e
KJ5Qri9p0fHiH4LvH3eiW65vvS1uqYO//AbsjmYjis7YT8Q50Vu6VerTEudv0KNs
1/TsTZr+GHiW6vdUqTgh7vmhfoyJt2PIcYFZt4mNHYVk/8ydt82/d9ioc1D6SclG
2A2DMR5TWkWc1/P6bNFrc6ANbKQItdzLDIhtkh9Xhig3dg9PyEQq3tus6h/YFh86
SB9c9KLTjayIvOWEjj5/Y60pyjvP5Rq4kh4Mpy6vATeZoQ06UOyZ4P2BHSq6MzvC
pIhty+sEDdEop2JULDu7TA8LJ25GzQEZrHlNLSvMFuxjBPMrT+jxNj8ZdU0Zdbup
OESkIL78iySXgKKAPEuntOQ0RRUnLw6qtN2PNh9PrXn+GoM3Gd6eV0ufnf2wLc3Y
+kY2pEqcrHuB0ex8o/M+kFBdfbKNmIZiZAvRqmF04RDTfv+8IsD6162SMj3Ov1HX
yIfhjT7R1M5AJioHbidyyB0GuHoQoS+hiSJk/eRdCnutNJ2shKz+UNgsuE7s8rhs
xQtx50gvSij6WagVApT0c20h3n2QcjiVLmqkRmRoWX52hn+URMdLTQnb2nC4pIJg
llO3QgeRV22mYXzs0mzLh8nhXFZ/IWguZz/yHNy9oDKleLpNtU9IRGuNQSvCstSA
xgCM5TxN2zLEYx8a+X6yT9Zj4xdUFih6TkbJOx9pNpV9XNMQtvYXHGT8ZIyt8sAP
h6bmVxvP0nnGjZdieiplDSzhvZMeS2C8q5poYIGRlLvJ9azkEh9yGuWd0HBjZkHW
raV1cu6g3kQE1mxfBJdMmMfcTNyebNbOScpzl3F/q9js2996lRk1Gl5e6FSQvom4
MDCCB6kP2R9uzoPk2n2WoDo2Qk8hMwEGxlZzjCiTklMVP0U/x+nuZXym8Ft7jpSG
L1u2CcDeXgZI6kNnrOl8NbZiZbmnuQvQd8k6qL2PLxs+jN9JTSBZuCUxM+jsGb/f
5ZC/POihHQyoX1z4EUvPeRXVs2MYjv4c2/7ePNrkllESmlA86Zk6QYUoea91yBJ5
5Cdj7jDn0QvswdfobFMXcKazDp8Ys8QKcSrj2+S1ZPHPOJWVG6z9bHeG7shy/S2E
Ef0fo1rWzx2r2yQpoC9lx1Z2nwbxinKpqL/5rEd8v0CdOSKqJhKMyU9Ex8/o/kGO
9RlHpqyJskhFNvFuF7BYdinihxoyO30H6EGqpztsAHswaDlItf71L7aCyXrhBpNM
0sK9GpF8s9EooJ1Or8/a9kXXHAal2zHYbmyhLXv/ia4z6Vn2kMh6VJrnnLmJrPae
qeGCaDmklk25sRyAkPvfCeBvChuAUxsaznUpZBJs+Zi247UL5O3mW+xbynHDTHNG
ER5qbWy/3WLlfAp0nqqKfyVuLf77emxqqiWeCBBZTeIppfocC3UAdBKEg0IVb7f+
mcHRcnMZ/dVX850QleLKqzXiD2D+eDqoMtOqVE8JEzJm3/UrwgiX48eYrnHwdhSD
WWrAMcvs56IJ6RpP3HeGaGITSGqU/cWq89Z8dZH4rz95dDuoQ/2jnPEDQvInWOWR
KoM20bJTCgFQz1pQsMauNQpG22rX5GZV+Wlev+VUOfJW4R9htIwA/vRzWxV6W/9e
ITr3GOFQBLY36SkUZdVcIb4onalPaCz/bUn5IfRV/NXj9MLYklJbOYcJvV7jEG1i
i63uw6jtArVMErUz4PntCSNtKvPq5HiTgp009kwVHv5AIGbE1PgyHCR1ALiso7d/
h3k/14xszmyrWCBx4v7VbveoFsNeS9kwr6e9m+GuocaUzlYUBwA2fQD5ItVHnKIl
txEp2Iw8qkw4jByti+rszPKGN529fpFzsfV5heV0agTXqwd3ByYMfRSauhbGyOAp
fV3ONPuGiavVYLG+aZsmEalg2QqnEC9WojbGIri+FhUEDZHwa8tRL28WU/47zE+E
lmTTAVP2Eln1gqXXO80nZ0/q1jV2bxCKz2zxtEiDxuxH9vc3jVpx4u8zpEwM2fIw
J6M0ry3+m3UAMOZivFrGmfttaw2kYBMg32sy6kuHu5D1guTvIhD7QXJFVTD7EE4V
x+VGv39WUha9WW/exra5B+y8HxEC3rRNgQRWN07pY9Oeh0eYQL+lZ3ZpDYSSyCgh
Bsz4sLfihywoh4aWaW64ewk6vefznIKAbZHSCsjJM5HJqy/PvosF/ARPf6+GRUuU
YzU2MWakwQeRUb5Xt1QBEW0HGosB8FFDYkKnP1RpdeoZg1rndphB1c2ACRSvQyql
h3+noU5SiSjGURJbkwSObkcbIhzoM2Duj9bHkPThGr1swYT/Eorpq1yjEn8DIwJR
9OKVLxSdfX9OQ1Rd+G47MxEq2aj+ga8ik/l5BJYo6ifYEuusHw1afiTGgvjPF/4O
58jZpM8mP38rE5WNT/byZbD+sZrJd9N8Gp3+UFcn9IoGujIuWbM9nWc4TbNdIjF/
rLuN1r3VumbHQg9HWCM9yn3UguI8PQ3RWt5qxuSDGABFGvKQvfpXUFj0hEMPN8Q8
5zSjt4WCP5JevB8AXXEXRlN70+Bw+xz8NusV8/q1xJigdUmSuBNHYZ76dH7lKh3R
CW+/P79HNwROoIhUSL0jbXVNXhGP/WLY9jXGELzBXjv8OrxTWcrMMEy750jOPXUC
ltt/ALDJuIXQs7DzwjuwwXvp0Gk4B9RC/t0uJWnjyw8hkYJd+KZNNdSpyR4rVbwT
yc42AnuFcBBLesEBiKuFA0VNJC81uJimEhKL8pIHsLoV2BRKrc++IcS8IpBKdVFe
TlcUPgFRH5g7Ot6b+LACL0njFOTGQv+5t0vHu5buGdJNg1+X4HHNzhN9U5Vi0++h
+iJJJh/JP8vRqrARfusXUCir2+PJAY6RdGspNNydi1RNkfBpvTw3/jZlfXnY+QoD
GuKq7TuKVmcGMTT3oYGreJSqbeUbqRtN4c4XKFeOdM4FNGAaxwGv6QeHQJjW7pZE
x156Esw6o9KhPtBH3dlslGw3fScrbaHvzz5gMOux4fTmx6urDYjixxslkclmTaxc
6OnRgpNPiRT0l0+mF2VdJBcxglY0AQaL4MJJyqJDQvbFKuIa2tJWr6ru/nbabMc7
gR1JrzrhkVtAi9CoeC43R+ktSxG+Bzdz6O267/0iCIYHB7uU6RkOIT/AlNkKBpJE
POSjRNxAP/MTdeR8qdYNu0+YIS80Pr/I8AJA8LcbXIFLHQSvXhMSqh8Qxuy4yBef
tVFEugTm5l54NB1OOGMfbzJ1zzaGirp5eAjUYNEURfKcm7XEyiR6cMMFiL8c0k+Y
Qv8TVLmBhVGtQ0tAvdHlTX4m8t6pWat+622OCIhVZ928tkL+ZI0RNj2ro5vpsUve
PJinEk/ED7jUa+3sB9HA0AgBNAXHA/iyy9LnWDGE2u1MIj9ccX+CXmjdF95qVLx1
BOh/SR6E6+Zpa/zLrqbtck7TwfKLqGj03z4Cw504sf2ZAnw1v5b/eWuhgzJgGZOP
dAs1WxmbQv4q5U3ZAI6eJSttt1Ylk7TVzMxt95MuSZCqw3JAfRqBLM65uXt7mBUC
bisR74vxUUSmMr+YUpl5Pa0GpV/rL51Axxv069dp5ugaSV8YU6R3sI+fFj+nNwJx
MYWMuUnBnmbZva7H0rgBvXhsIq5it06bQOCoquV6f4DzQaYPSkGcD7a8KoWzaOhO
k/RI8lDavzKoJTDXILIUq7UFzrqup5QZYi2/CxUcxAB5eFDsKsaX1+rt06nqAU5t
rv+6lpLk0v/pEh1Z4Mo13l6SqJKU+x626DakV/WSZ/eX/JJ6otm4kCSEEtzfjHIC
tnlGeXDUAGNotCwKj0cJNzzvIC0shtY97VV5clsI97zjK3teUs8E85Sj0gkDYDx4
kx3kaa87u4JAPhqQnw1HBFFvz/WHLzDiUHe7mKY2Z90RBK5XiQd8j/77qfYFzpc/
Pu+/dOJLD1jaUoCIXQ35mzV+xoGWyTsfL+oBkJsBuc1BTJz+niAH88btQOzuWnLi
yTIVkDemPoKCW91UD5rKjfeErH5G+1CI17+G6D9d6NQPxQe/BGbILV7KWZOFRLHf
hOfB6MYqL5OTL71PPMJXz6w1DHa/KkqLMoTmK75fjjgL0R7PARDOVRm06gEYA34E
1MVcDqWq1vDIoPmqwgXEXGadkvmnbj9pj/RUnLw/gGyAg+wv0kSU9yCN9f/2bDWb
AzC2NhnhfaZoHkYCZpZokpNAvNJ/N6BXPeFDhecqdjvj21QX/wbfuDxCRkmXQIiQ
iqDjSAG1CJwXmCHGRNwjS20zYDL/yth913fryIK/4pBohIuw7bJc9beBWPfvXGOx
mI3WkmKrzzVlC+e7rJ7esuVsO4a1XiggXeJFGmJkz1XwGWyd5k18K/lG4MrxRKo0
LjWw2ij7aXmg3eUWpHqErgtwk4v3R2KcIh4C6BI2KFfVB999pNMQdPhYhd1LQBy2
S8Gpi1EdpSNb2q4tS6BLqi4IB0rOXNZNPW3lgV4aDmDj3ynqiDyYJDQqz3ISXyJh
rvFUft5i/W9aaq3VLSDQbXrte0mAaJPiPTChH4AaDpNxZrJwO9Nj6zDOOyP7DgvA
G0Adud370vggwwgUzWh8glmI/QviD+xEtiM4dn1WANm33A7LyuQ2ufc1wJQ5kTde
C49eQo3zfkTOScT4XAfJLLLELVMPM4DzdJd8NTrZpxpf5DCBZIfD73mytJrI46vp
rJBdVfbHVlj7ty3bRC05+6mk5k0mbJy1OQ7+H7hHIxlXVXteOd54rQW+za4tGlMo
Hg9Wv06y9Fc2mZDBSqs6TtXHNFC6fGI5uRXefHEeeAMRKbv+H5UYDptjbDldcGHs
FKXIk0ecQo35TstY6rI6oSm6rHBZeNi04uSFeCdeNxLf+xJARrmIpqcVLx5cBYHr
6lDmEBIKbQRpNs1XHwL5mtYFE/ucq9bw26WMWSbLxLoDhH+khos8FwHZBirMr6+2
4rYndX9me+DOpFbQaKhbtYsIyKx2S+pQxqVrolYfAt9QcRfIxSPnGPdO0QWDjwj6
CWHpzf4VjwTlr7Cy+vucfXLJ0SsKxQWOaPIhKyu5b7ywm1rx6rdXgqFUy89t/Rjc
LdB+lQZCx8CAwBMMqrtk2rXWxpFeCiufGW5N/mr/umt4mN4vc8Z8+cR40WwD05AF
djRX5FT01sz4ODrlV+t5pke+vXmcrOE5qUx5bnEtKVjR400Hromx4oGsDhR5w7kH
DptmpPT461MqPcNWDv8ehe51mXSnkUrSGdy/Afm/piV00GROrLHUK44kXg3kOrgV
lwN4NjwbLYIgsGcBmNc3/3NLmKrLXYAZWSDV2MCoPFA5ralYzIyvBk7ExA2lisls
TD8yV2n6353MTLsxS61rdmKVlZgU7I+oWCW2A1DQgoXT2S2KU3hJBu4f0qv5+Wvt
G22ThiokRWEATr5tpsQX+452n6CRUpn7UuyeqLqkIO8IeJVnzK3Kb1d9y1cL0/Nz
vWuRh5B+CDfOL/z3N1A9F1PTcr5eM4keb0mjyh4e29HA7GP4/JQrWKaNZM9jXTR6
OKQ+CllABc6XArZQo6gb4kL/ncuL8e+JUJypAVJqyoz2z/69WyuGFkFligT38i6A
46Bv5tvZsiqXybbOsw4NjQZefhy+U9ymP+jWgOfF57f1IOE0e1zGwdNpdEb4LxIF
Z1SwGTfreE/x+rTj5jYCR0MA42sC4lj2m8HS6DPWM8tKx7s+gmecxebUTLRDQHoe
a9qfI1ei55a6pCsScVWHLFFH5BMiK6l5Ppva48QEMTgUM2PjSQ5IX8zGzKnS6AOm
tKxGAQ1E0EJgI0WGEE477Sy7neiFy9qeQi+IE/mv1BAy3mhWar5FmvAkWnYqgQjS
Ap3sLKnRIwhzdpO+lZ3jG5XVq+wO1KPBQ7hUNEJ5OeOnT/GphBVZjsyggyf+VBeE
lHLTTVQgyvtGoitC71daKBNgy5rG69z51fuCH6qb63n77xXgAWuHriommUe5YdjF
fAMlx2Q0NAIDqdR+LRS3EyaFdsVp9uF2UKfF9kKwQY46oM2RgbTWloocm/tHVk/5
1vWMOH14SRZe7CYpPZdUsNNN0lOgZ4C8DeWxQD4KQHghPXsu9+IYsg42JDUnfJtT
/PA6i8xbRIVBTv8H6F+niU8gaEs0v05WWDRm+tpzXMStlsU9KyuQqyY2vzsGOhKd
5kKvx7zLB0NoXd1kbl6G5RQHyVItTAZx8q5XHai6ZQNXDGU+hzwoo/pQCu5jXB3u
NyD+CkbJLB4dOaL3/1oxvNl50PPZLEMKXqoeXk3FFv5ttFAkhBpIW2wgrhmwfxR9
g+y3mHj/B6VsOuYYr8SGaASapBytXAy9tjMfeHTTOkmx0vuzSuSz6L/ElfT+5ZxD
eztsBQUJu666hhbtP1FoT/JQdaRIgXCZuXu+gfrSfH9ejG+02XR2A318fUKSN5JO
1M+T0J19D52k29p9VrpdzYQpumCfpsyGCUNGz0DJnM/r/1caWUVWFYS545xoUGn8
v2rJWutGGDTgQoZcKLknxpMDOT2F5A2SE61Pz1KF/tD8m3x/HYDjnU3PZvQjrQZu
VIDN4TQHIPykwwzn5tUoTc342LlPW2vf6bwbWhK7pxpaPR5C3RO3Glp/biWFpMeX
l9nEjsBdl84Kx0ua087jBaTf4A/BWtzTdMbF6Mxh5wXZGrwFSJovrY+8Q+DfoeOR
1GbQMulBOJByvoEhndKB49+8T4Q0SupdOPgOgwlfWSp7BKaGuZnP0+U/ya/ZKXtY
wTns3QuOPc0DpAZQ1dtkn1SJJIe8cujJETOxNNz3Xh6M9hOR+UG9jKzZEg98bRtY
dPYYvv5mKHa9obnP2jeYkKZGDavu/qCYE6dFsqURJ8PMraFQYHhPeGJCk5QFcjdX
keexmSEwzShisGrBcUbAbAQdVyWbaco4Savx44NbrZ4PwHerEm7YVsUXmuyZZG4o
6G7jI5f8JZMtCVqAXvCWldC/OTFocG8oPqe5lX6hm7HA+78Nes/VJPm5R6QhiePF
KN3t6WifNrO8+4Q2cXGPEMkbrt0VS12ub1pw15tjy+V83Z6EiUO9k4eSW0mJoiFZ
MITjAZVYIh5IhXbfsfqbNvoxeASw6e2P45in+pUS/Q9oetYxZjrNPTU8b0Gu8368
ib/LYU197KzkxYGcmJmZHB8FDiL+UxgHdVQ92WB6k9Ta9BzfhwLZoamFq/B6s6Z5
k4vr8RhhvNI6kkOVwNyQKiU7o0/c82HX5HGbmEgbR6ZYHaLT+bsUGGuKhIV/hhmH
6BqmgqDMaozrJc43U3pSEivuvHDnfCgP9IoZmsPoQxzJVyaXPpBzqycLTNeTUoYM
rCejP2gITsmTntxnrCsQFPMBKDGylVSTaN3XJ2HNuPrJnypO2YIyMWQOg0XpspTU
R1tNqPkEbAtHOz/jnSPEx1/gVrkVk5L1V+ZUPU6vfxiNEw2mnWWo3cmEgx2w0EPW
v1Fc0uBY3O9BBhr5rWCDZ7/xZ17Ca5ZbeKf1sXKp4XUorc5IrvneInbTA1HJo1WM
m0ButTdReGdy+byOEHStofeiW5h8nlYvrQpVEirQMfXIxKGaYge9nelF18X5gQtt
5lD0+s+PZ8FiUO3Bap6aIlwyiiT2HJf0KayBk7SXC/9nc51nx5IOssI90ka3YycF
GRDRkJpOSAvXJTkURcOyk7k2chAMPhWjCCY1rnpyhhsQMSRn49HFdvad8Z/E4VdJ
wpKYyGKNVSCWJo6w1fCZ5TFJVuCPHfAZc+6ppTtkPGIrEUJwroM2mnk/L42vvMpG
xPkNpZCAUdYrxHHGo/9DV6kcdSCXW9Bhpfv/dQukJT/f4RFqKn/JTTGLp1TuO2Pz
ALP4ocV1FDk8pdqHJNabcVgL+FA4JnrI109WGZZ1TB+0h2hAiGW9/Q2vJi/2dCdl
JfZkrAtC5Evk4DoHoySuDmTJp6BeRlhuO7DiSWkmCXmOOupXrD4RuiWlHyBSW460
O5kxsK/L2ktVWZTWuKSQOljSn4DV1i2VSP6P4G8z8GKSBXNrmvE5iFew8hfWZsto
Wnwf9+cuB6O5W4Vk/0cFjkhchSbcHtYc6bQ8ZqrffeVI5BzWAduNYs9CU4OlGbrJ
BLD0tkwJBNmOIYEvuptZ0JW91CIrqll7d3yyO2EbDqypyyOcaMqYJSER5yvBtSrQ
VUfYNmpiczjzIV0mHHr2cizTIvFT4+B8QAfTzYn06SR0xlm/x/tPtKo1sFMz1oAL
5yKvtPGJNy7KBE0eWZ1YskScZgLc16D2U6qOHUl7o+XSnUZv0U8WlNgv+ja8IBz3
qz/TJ9dztaKf5eCKzIbSIRP9Z0V5I9/T18FE0j0mewlKgTI/qhPzzgHtJekYUObT
kpGXD8N9KX/33oGlvNbBaCyThobDM/chJPID+YRPghvZE5cVwEmrjBlx/OwUhxpu
/I6lPRUPIwV0Qa4XfHrkA5jGhOPPh6r4SuYT7yketeNKPJqS6DhZEdze0c+VG+X8
4rVf6WzyBBGRaQPNsj2wTL8K+ZbLm4BeFPnJdIgeoZW/McItnpJI4z/Wy93wAS92
U3WV2EEH7HR2+n3l6LHy/E/v854FXq+Lam6VN8yMyshoGYLVL2HClnuiw76ykFU2
Ks/8fOleACwYB4ejqzrjTHOq3+g44Dg6XTzaCB7GQ+APBixOrNd+9WPrXL2VSbC/
ewSfG88u5DWyrSEFU8x7/1us1dCIbp+s6j/DITbhkq73E4vqQZB9G+rcqLg1dXDs
eeqNQlYDbpruOhugsP5RCosgSpKA99egO5Iaqg/H7kq4Js9vm3lAQtqD4eLsom5H
XRjrWsvB3hdAre/pev87/66OqQiTHj3+SJtIFX9aMOMQkJbdwyijBvp1L+WdnQYp
QR3GOo7XIKF2DnrB54kNX+GGn+kcWTvF1wOEHpLnsNxy778zuWMQYCBItwI163Zg
uVeEvKDEf/sIUCC0w0tobwa3Vwbi+8Q049QIEJop+TjVai/GQU2hQ37b+5AoKbB5
fh60V/Y4PsdtNLvMNp3pOdBd+Kco8ZRNn29gL0+cFuntsiMs2MDHTGnJc+8E3HB/
B5srO4iy6PNcndyYCKfhEpAX/xOX/l3g9UjS7qeZfmmloZ7O2FnpFiadTi7cISqj
Rf9Ww4tT64amdbwxuG0dhBLITWXsljGkdmGOwmLClAAc4OdZ9wiAVHt6hgNZU7Ur
bECaibbvTNl+w7TrMu/tDQH+0bt5hADPDBEr1EKxT8gLKfcej+E4SCaCXLaCHgp3
al5oPprhDrBlwZqoR4JvPZleqPQS6Bh78YiZueDFbSPA7qIoIpN/DCRnLw3TX14H
o6DV1ajSMFQMXWPI2Ygoimb9kCE2zGorr/JMDljbkvkXvFD/YRvNKo0WRE+KxgjE
cwgUPyoPFweTHPUhkhNYxU3q0j5Kr5h2jzSOBpUlS1HGmjxNNGcNAjdNQkVqFMlG
fspHJ9/AiKVJX2iS7gbqY5x8/e6TbxzZ/pJ1xsD4qIe1Kp0/9FREMRbia8NkB97R
K05PygAKZJBaM3CMcGkJgrgAkbNaIrJ3nEJl+TmGiY7FBri3+0/LtYi9ulRe01+P
dyuODClAbNiwi5EbbdcOQrWj+Tep9j2DPj3BBPfG6NrYd/h5thtKatvGyuEMsqBa
ywUy2EanIbRHoRKx6lqWe6NyFHM8UnTmekQbhM+UfvFRII2TD4nF5f/+moExrfXY
M1kVUckNJBcGjJzoVssDECk64K2RYyiGixT0Hf/v2M8qfh+3iYknQJupTh1RW0/u
NNj80kFtlC2CFvUfsoESAfGr9nA67YAc5Vl+fuLtm74mhL2MtwHHQwmSo2mAQskk
k0wGHQ+0olemoc91fB4SsMowO201VtlhloxzioViNFD30mPrACV+W7ZWqw9n70N8
Dc68LK93sOhNWU+6f0HJEHpMzd6shcBmGVQ4546Oeti8L+nD0c9/74x3ipE3uuhX
GLxO820wNokwBe3xo8EMNJNYbKYBin5f9zPZLss5iQ1JjW/XxsejQZFwxgs+5T9W
cgAfZY5Z9EfSTYlDJ7Gi9egsDsSte2Fnfi/vGXgDARPhj367vtrZ3biI6lYsohYM
a4RN16+13XKjZI+s3LphEgBVGvPpeE96pm5NVVCFpLoX7HcVm+bhVJ8DjXhNw139
uOzRXChgQoeKwgz8teyp+hprAzqAF2xn08LYIps4dR/1G1ca88cnsgaLXW8ZipH8
XV3ZlCO+fWAnYpSxa5VK7wkDOHNTQz6/gAoiQx6bgwOQKxLb7pJqrOhubUOc9mmM
I+uCbaP9qY2Yk8XUOStjyfX3nQn00CUU+Yhx1zlUOv1StrO548hXgKiumXFZuDhc
y1CG09u6iNP4UpbEgazEf++a44BPzAS4pRdbyNeCo6mJxVnxhjPhv5xFm0+SW7UY
E8FqzbEuHLvC9890vef5ASiOmxHY3PXnmOx8SrA2Of9O6eAjUXp3pFFHlxqt2kcZ
robMAcIEV30GvfGKb1glvupYyinDHYzm5lC89gFx2NltDAbTuScYEnvB47ieMugR
lBF5ir/d9LYhomtUtZuxGaX3Hi/nK5g6bQKelVPrI0hdKyoYnoIyfOWGq45JYFiT
jd0m5Xn2zlj9I971i8Psiq/DJeHGKjzL8VVqB5BREXnTBTFsn17t3s+GajYNCNyx
Oqw92S4twPoKymxOhSL1F5RiNyCJLOckzLJkmF+gN+GNw/Zx6gFAvgTp+GeeQ3zE
gLB6c5dZqcrt+7WI2vdixU4MtOEPfZFbxlNAp/V2PGY9Oj6Brt4MZxQsYjaNu9TU
gRNNtLDlA37XCpZ7NRNhc2k8il1nd99E2mwNY8Bm1Zi0udHVN29vhqQaOlbcRTRZ
RM+LAMVZWsZfaOKE86zHWlSDKQnCpjYsWMqb5welPs7hlEc941mIor5tcxAi/7p1
pQJKK4TIpM7OpIbUrHhcCR3+uTTrCsItVYuhGIaq3RIqlYDgpUJ4nMLkT7UHzkm+
g0WW5ajRJHPoxSPH7QwducLqp3nQjONzNVWDHT8zhyxWKl7i10tb5V/pJWeJK9Ag
sRgjw63irt2H5yVM8e63b30qLR8SHjNs3DGgMJk2HGtO7CPoGb/ndwG/upJBHBLv
j0hRsio61ZEZTzNb8X8GZbFgQwz5NeXs+eyEb9kGsEyYWlux84N4NWetcTNftsVD
G4eZqf1ibOWeS1l4Nl4gu8uFXsyhH6M0AL/58t1fssAFKRgY4Rto8sXyR7t2HhJ8
/4tG+NF7rjJ7X6y4EtZQ1mxNdk2el1rp6G1kC+5Mj0UZZxtSQ9tbOZ876Zwwm3vo
ZyOOiJmYk6V57B3yxhggTnAbv15tCiDTmZXwY5WXSvwIGPjkCRHjrO4GRn4UnkrI
AuQPbbhppdGIwkFB52SRDpD6zrV75sAwxUhFOUYBU3K8oFDCp1xQR3qweYwg6kAp
TvCLdUKG17MGwebiPbvOHIrvN0jutrIE4rlc0Vd3WxLuhirWM4XqiFZdjMs/YwVj
dqaJzTgxNuyFLfyX0lrRcwlWi381fFjXtaDqg8pLtE30Qr1eQKpPxSRTwywLoliY
X7VZTqDkdcECo0qQNhA/o7HraKBsMXNhx6so9bqqLceO6pPzbPjjChg/CdPGGkFQ
V3TpHC9d5+7OPOoDTKc9+xT4nPBmC5RHdVYY3g7H4nzYDurbK/ycfrbrTbOfi9SX
w3nvBL9tsswYEGJEwBC2Ix3oEihpOodDsH8CpRc2SmebnNvvNkUmvuMsVPLGxAmr
+10Pbbagk+8FMeQMrTis1j69tnGTkrfK/dn1JVuyLP/PTRz+ythV08czW+b253ld
Dp9pfDjaPzOIOQAzE21ULnIeQskrhppKWev0d70K8gXKxOT4lfxfz/EBXCjhm+Vr
GW2q64tVYg7JdCmoBkROp2u/tuX5Dtu7jr0gG5lQHdDvbnJXPf5Pd5rAoT3TtcYG
IOsVauQ/Qovyph1HbL7klkn6/Cj2Ob/SOp6dIekImwLigbGdw9QrONMU5n+zeoyo
QIpI7aZ1KOdR2/Yu4p9zpi4Qv65yYKB1LJVS8uR3K/1QbIXCzpHWzVWp9fFDceB8
FrUQ+dwiEb3CowU5McF/Ozs0rUkXzfxdeN2a4bQ7aUTBOoYGFx2lJRTi0F+NY53t
LOFVFc1MLd6ksAMkZEQt024dQa5+Sqz3ZoYVM6YNFNR2mO7aH5ijy4EH7vY+ymok
IIZLgHrdbdOpJj/WtqHMqNzTXQemHUpw/xb3hiNEnRZxSBjZT84GdKruupYIPss5
ZovutfCtMOwUC615jekt53K6ESd0+H4hq/hj1Xm6DDlwwsYtq+gAlLLcAMBnAbTN
/suKteIli1hrNnPIK+zHfmNkrLoFAzU6jXWHKdr6//2+mxXOHAxINB3oOkbZCsGn
ZL69TqaGGPdqX5fmDa23cNtAE7ktc0kkHaWSQJCqh3mapKfyHL17YjaPHrUz0eou
rydWT0ojsEkA5YF7brr5/t7Ei0QgFVVIUTYoNI0Fz8F73al7vKrMYGB731Jui1Y6
L8on/4G7NGYJNQ5RfZHpTgKP70Qy3lQSbIbo4uvMDNVGQeL/6/7OKeF/+5p8QqCc
LQnQEF3bnRGx/rL/aa67TcAu2CIK83RBVgmvnViRwRJFaDSx1K00nEVnwYh4EFtv
F9uLoHfY8lFtFajSPgb6pswbFpyfAzjHuYC+YhCXi8h9cGkWkKWooU6Ik7he6LOH
3HK3pb0DI3OkfcoAKF8LbYUKfV7HdZMpwDL4ncTKTsAUV7eX8LEyDh8XlZlHeugq
LaZdQsUWuML+sFIhreHE/VVyyvaJWGY0Rwmcu2MjfKR0DpxrVwjvY/G7eUFV0Ti4
Ull2Ksh18Fy3i6JnUf6yEv6CY0zN0Mclk3ySIRPA6AoQ89bjn6hv/rJhlbXny1FG
SgBHw4yGIaby17JuFgzQ329GJaeKNSsQFw6WoEXR0s9xs9MrjT3x1eIozF9mSdAY
64S8iAjzrQXTnXb4ilzUwVp/2krzPnOggv7pjbRNvYJsdNGhxBcPQqz+PAFvRJXK
FUDUy4kSx50eoyIv9jZVuDDJ1cHvdI5BNNKt1LIg6dMmGi3oQKNKFKeq7kBermcw
ELMeAyyxAbmGlhNUUTpMZPV/sG65vaFjfuUY3YqXYnELn/AojuzQxmPC8zKw46B6
qDEUqFbtG05JddWRhBmODhZTGFcYECUZ0c0WvjJFF8c2U8MtO6nTLgrlFJCiYRAc
5xCKA4BzRN6PuWgNI3YI1KvVSXBeQUWwD6BgLBcehFAn+YfQuWgul8qDSt2mbn2v
Tl+WfxB9kul4UhMtnlv1ayA36Cj8hXBZ1Gkx/7SNmG6W/SwPqk+nOBQAKo7nklEx
ha6yrQz4PqNwBYOi8ZZgJDrhVC0eIhf19G/fF53hcjTiT3ynaOGlsQKoxbuVZiH7
Z7MaCY+bpG2tPtF40DOq9qe9nHUAZttVuNZ33BPmYpL5oJ5FQ9MqsWzpgwQnnNJh
0mhohO/YSLc3Pqt0aaHIUj7I9TLWtX62aDlz5ZgNnkUIjq3w4mttSzmo34vCHuOP
Jzc8nAUszjrfEkKwgxT1xILRa97zRlTn/sKQAFgqYH1UO034Uz0YFigIR0n0xI6c
wS80A6y3+6bEm7aB+0GzH5GVZlD8L4JuU0ufM1DbuSZKUokamlwZ6naRG2ZtVkv9
CdNWJDEeKiD8O/hcDXYXAHQZ3Cct64tkrGshIgHchQJLw8XS0VWQ6PGbs5aNf0be
wUZXgVZhAReL1zDfVxTMBSHpaeOqFDfhhi8GJa6wT2FSKRXHL92VYyJqvC1f//Cq
xSq9wPE6dvmBzxkHRahJCpslV84+E/w3lHtjXznyyDWCTYhNw5pIXoLC+7dg4lNv
Udl1rua1ezQGpIXWvHECQdE5JVaZvme7ZBCf/WmEep7UUgkC6Dtq1ljVlIUl9mZJ
oUEev2HGoAWT+ysJEmiUwX62z3mXeErcsNxLvtfyURNv26NYUWYELxURoXE3Nief
AHBGJbJW3WxjwE5CqNW4F4dg8MABPUZD+Sti9+zhQMzgaoi9uyyIOB1wMLUWEjz9
TeudwKUft5WwuEHvY/V5FSyhS7DU9JYZp23L7Dty1oQllKMA2ENGXr9oUcVCB3hR
XbrMO6wGQdXTr0u+n+0hhHjesY0bbVIXvp459jnjn5xcVAT3/s5u+klJ+WlTXGu8
0wF9YMsoA3/ilvTCCCHIWJGPvPstIwh/m7zNVRBEThpKDwxeh52fbnseoDWRVRUi
qrbOoGrY4G9yevuMPlcooX17R6lao9ofo9NsU9Qm1E64RVP1i7rCtNwiOvIlfPuo
kzr1rnVHPizfxLb9Qc55wSuUOba6EHTCWVUdeK3UeM2KnnZX7zNhZ6T8SvuMYLTs
eWsAEFb6IQbXS0UUaQc/CPQfEDj+Pb4uKGH2OJVJ4jDA2Y4CZFs1GdeYM9YwRwhj
iPnJ4c4IBsTP+8ELhAlMxQko7vMBj3WRT87czrUjMeoWt2D5Eryp0NUzjK1+NDEx
s9/95QdPPnzu1wyhRAtKO7N61BwidJ4/l8qPvAFi5VaMGEjb20o4OMZlEKPfasv/
ba5V6HLVrEbrd0+iTjkBlmsMWiGbrUVHDSoEzoap7IhuO3vYI4SEysyuNPoenzO1
qsbt633vwLTNIGRQXdkw8JX7ZM/EBOJl8MY7jgNDl9VxyCQ8+lR6m80PATSoOhSp
ELH1l6FQDz9RBN93e25I6Y0eMAHMwtj1XT9Ufq9OKDj2xBcX80hk4t0DKcOfhwE2
jJk1bEealkUBZ48NN7CE6qsk1rAzFpokRfJbB1GEEwhFHHXJu92cXoDhNy29fqkm
oZmxRZusvLdza9ZAuVhs8s74NAT8KEblpXDMVPMO859xRd+WbHHUxo/1+Y4IK58d
FV4qjpHf8y63vsbO9w6NGBqMWhdiye2dhOAZKBErhllnvSMhhahIyfIyEL19YaWj
WIppvRiWZIx7lhO7K1f27rTNswjDIn2Jm1HNY/KTPjXSanwjmBxXpTTRHgC1za9V
jJIYk+EKnPUI/LzNA3IB3LjDkRwr0tg2Odh+eExPot9CKFgxJVYMZgBiwKbEF8im
LjCFmmidYTVY0V+1FqRSB9TQ/tUNjSTkk1Nl68llCj9VsUlexVfv8vdxm/42+IZk
j4n5blf3G0ef3kp4xd9TzPKKN9sxIlsz1lMq5jo/l5Il1GpANyROAyNVGXgCm64l
qxZ1jKY0KfgMY8bzg2DL0dZv2HZDA3Hw+B9EtbT39WVL2+YqzcHo57tXkfYiTOhh
XD0kaC7vbLr50RWJYm4rPxNLAqTSDQ16heYmF0RGBdejCm0xaIRUe3Zi25b9K0C2
r6pnERLnOJVmXSudyxM/JnkpHat9CA4F5uwtdIxcvImLeT/Jat2rIuj0ZkNfoEQ/
P8/H/L4nMWXZXkUhyLmpcXdE9/Gq8umqz4irdZ14XbUWch3XsMxqYpRhd0hQ1v8B
efY2PbXVG+HHfZ3AZ5hvCHqx+enTe8X0flNs9wZW49UO7o1ytAw3Bkk9pJNar27h
QR3Wn4TVipNQ5Sqh59W0GJxt1MT07BdABKMrR/nLav7141S2O5wKyblYMBuO9OTx
cdKf43ULPeDYJyuRGzzMP1rEArlgB2d/eI2vVxLlSQ7wx1meUc7A+QeznDOHPuG7
pjgpy28I2+r4omhVjpRKuerBIkijVCIntTT7XVnt1gp6aYwuPuIRCOWlugDsboO7
O1m+b5bfjiUGgngbphNV1iGbRaIzfO452mic6CsiWP2ERflnJ7yE1vmyewWKTtqF
AL3kxwMT1e3XCPe1MHr8tcj1GP3JU4LCY+3FQA4kJFH4V4NssQIHMA49L+yBXZEw
O/tSnrSek/8L6UkVYC+qBMGwf0dNu5rw8YDuxbIDfF5d8xvIES679paunevu+RkW
2nAffSvp+R54Qcj+6HYJPFo+oqNheorw8U7C47b7Vc/F31G6LBqfI4AJXh0agSBP
EdeK0roOe8mJ2x1A0/Vx6whTTw/FQsyu9dslXWC/OWp4LETXSybTJH/7lCWZPvxv
62LECz+/QgWBGBhvMEFuUtYtceT3a6JGIek02zoal8ZOyjEHSVIwrpl74eIRgou1
qeeM0wvbaYMF/5TmmbbAuwcBVTXlNEaOAq1ucH30w7FMChK5Qg8qkp9I+TPJdcae
9qaOr41LgmVg3jTggUCR2Scull3ISb+6mBoX7zJGDWGdsEHjT1h9upM/9oWN8i9F
z+suvd8QupniFj+MY5rLfBWXdV4eaJtlZWkRvDN2nhJ8CKzbf1RRR9rUeiCg+xDx
+B6SEBOV5Qh2v1Zw7hAVrWQnaRoCNg8SrSasH1FQRhBFD1u3LNtVr1mvWIpVy4Vd
X3Qtl34TWyoNiIJ9sbAvXlsMzBRKMWOLqZwUxnWCqvLB9inGTSV9CY9nWg20p1GU
Nqe7PQoJHf3i3BOgF+cQsXc4GaiyQbBpPgi7mTxrJMtgmUov5wMcVG8WffXOBLKu
ugVmv1zoiFSNOvpoxzqwOO7vjaqndRi71wv0cAbmRx0sqBuoLMnz5J1QnWRBTEoP
VCn3svbO+GV8o6EZ1S1uOs23LhQyk3FrT9UBDp9f7jV6cEDaey6G3yDAe3O1A2Zf
poWoVRgO6BnSeqcYLhAEN5TMVmgD88l9FRTM3Wivi6yt+m1qk+Nw+orR6ZmEo1of
S5VWGckysw+FaZ5hzQ7Sp3Qx4gQiaUfH0/j1Ss0VEHbE+fzwR+YEz3FtoTylOxEP
OGHu5wCruKkhFTtd3dcRe0DVG1PtCzLDHz7YdByuoL0VJ5xUdy0BMujmSe9tcWkg
/bYrRsmlVxwkc3mC46pMFZxvQoeInGfXwd9sJZ3NIQdYpkXqEWbAyPmuJ3bxL3oH
0/7v3WQ1k3q/sxBQ19EZy7y2BLHRwtz556tXNJ/WF9RCDx/tY94lRcHJrNReu8Tr
Z2S6vg6JOqc/4sPzPGMi+95cDnAbnrLZcSzeGB/c/+ufeN4Vwsh0+MXCoEERfoYq
XiMqjagRje7CdKPU75JIaWHiZQ/80PS8P+tc26t7MmYKOcVmpqBHaqhw0yZCdR86
P4bDm8yzJYO4fOrvQliKcDxSLUkY+Lh3LnoPEgow9iNi8u2JWjfoqaDjFZ9Hajj7
asZyOyAixH7FtTAwrEdJKcoHGrkbgkMrzBMb2N6mRbzbXB1eLWAwLVmFBytHI+Mr
viyqroBmHbaqvJ7Axvoe71WskNitHX36SahgKbDQNYm+gIw1mHMo6zRP+LhXJXMJ
lQ7K9jcskizzlSw4qqzBK1E62XiB3sj8aSkYuNO2/KwPtC3uHz9i2R5nh1jy/ini
4KG+yfFpqcHpVmhNcFX3bqppq1ShAXm5J3u1eLsCVtRnqV95EOa21i8FnQb/Ug3L
QUzxmKYNXXlus+w8VbC2qiw2Ay9DAwuw5yrEFd855o3w6foKGiY4AYS3/1m5AQSB
vkyvWtnpmgJnEkusqvX3pVcWCtPreNsOeK1qRc8wM3ZXO7ftG7tQ/F5xk/9QAzgm
QE4D0VqEcZ+XomLIYFqjsN8jz6ZOBit+htauZQh6tDOHX7aCoBtRDsGGHKGjqkzT
Y7TXeny2H0bv2Ki3LZqlFqQVSJTfM9cQkIZ8EK3yxX4lXheHRBfo/UT8bevFd2C7
Ptz9D0dFV+0VyAnJ7wuv3za/+pbw2lhbjNIBo4Ys9nRoi8FHqx/WJmy5uFGO8NKY
2oLPvLgCqZa2WJCAhxot/koWWg8QRRQ73O0fM4uIAfH9stGiyg+bUclnDFlnASg8
M66oWxfBFFIscQtm00KKHVRzPj3nuT0tgDbYpmEtVGdV5hVm5977rMWcniX2wZXV
IAaflLDrkUNX/NUq4QPApNpyVkZKG/popwrmt2K1sS+qCaT+6tGzVYTaV1Dhm6sG
yOjPKo0yhQ6BUacPUztE6H0H+VcCmwpouIqxBJg+E6Urd7Q1eOrBssdORZYQBIzM
TNXsivRYiygI4AFkfx1VwhHwSY4twZreT8Ec27cvYouga5jzhkdXwrkL4ln72RWD
KrXcLEzGEh6iwrlkbNKXOO6SJbsNok9CqeOStdaKLyb8vS+50K5wr80/MsPP98R8
KUHayEIoyCsiSsNEQgw4s19fbhFzn2FS88Y/+CTwCHZmVFiGBHd1jEUoS/W7d2S+
aPS9OLOd+Pkyoz8ALEyHiforSu2XRaUwc8HPzr9iiG3mWgKCGbajHZLzNsL/lEZG
rt8d/85nn3PKq8CdRVvaXpAxGUeZQFCg8GPLeWigVXMDmOtmaKvM7Q2Fx4pXZ3Nc
eZkBtzmZGNGFsuwTrwxTQqIn2rsJjCoHiYhLKIXtMQmNQ5TVMb90YG+Juv/3iguC
XmXI5zKD7T0xtmeuduHDiRDunI8oPdV+r/pbWYDUl0TJBDW3vrTl7tehMOGF4QaI
TAEtRfaiOpNUYH1+DQriHZBwg/IyVhsqCRhEAeAuq6z7DkH+aQStkAuI0Ay+YEFX
DLacLtuQaLdGCbEjLH+Mfk81A4LPtPorQcumVP0eC4eWLUiKlShTorT71NvZcJVQ
iOoAzsHwZxGaoVEQdnods6Wgg4H1ERoTBtZwNdudc8EtKTCc/G8XtPdHTJ2tnrWQ
/Uo+pigBzYt+m+UJ5qlzw8yOw36XBqbwj2Ko2SEE+/IrgqLqCa/vXVdGyfitBoS+
66fMkFzP17zXTIlT8lrO7cB6MHRJck5tLcccK5oh7DWEkfKHFhHOgoVH52dtX2Fr
TtKv3e5oxa58N/8ukrB93ZPcVquAzH1StJVAD2W42yN5pDD7d+cCKzueIjYyRkea
V9o08WW9cHfe/hkhRb/0nzNaNW7TCgxooghFGBv7cowEE4yEkIpXlOtA4DlZ5azb
Lv5knAbAmZp1EyI/nDjI48N2Y0poH0Gud2UgO6i3zCdCYvImlhg1tEI74s5eibhf
u75ZVNeWF+C2wTwmBW70kLHY2rnCTbDYiECOMrqhFBQ0aNSEQdOkbpFnBzydGfq1
ALOsuFf87fbuknjRitixmgmqVVB5jr69DrEqhBFkS9phBVTyJaIbFYVKdLgH+0dp
9OI+hDIcJ+8lhjqz4MBl6WpMf6NC//21sOWJkcKFAfXrv1aLHAFF8uh/HHoTOLCE
bwTZYhCYOSiOKLI91NRJHmZbpHFhiOY7oEekyyKdlWvwTlXwdb3HizKrVWYGO5VL
EB0bc8vK7Eq/n05nwe5kBHP2En2bcVvuqNlc0hBpuGsAFbgjOc/ZNB2Utcs0qgQU
hrK4MVino+yql8wGiIFdR/SPZh06bM1iGz1sorVDh9kPQ/PLXzoFF9D+1Wxm8E1g
DNI7OHRf6CS0mfadL42f93cBIxfc2zeotIfcOBCF+2DDhfw68qPak1A45xf9iPT2
N/AVd0UbYCMyYHxbHNiAKhsWAyLeUSVYEiH2SueTQbkVjJnUxI9BekKXZ3JHSAHa
hmBApoekGI2MHPBxmpJzm2+XyWlLhyoue4Xup1YkqvQLj+vTcJzbqH3CaLF3cyPR
rZcktPUzjW1wYG9XjVcZsUQlUtMNqWKxoKMmVEvRyn3OttF0D36gbJ7UgU683TX7
bMmjT0XlGRJ4/K9hdC6lFUY8Zbc6lPokz4S3oVqmN6JBxDTo+fxQCyfnoiR+7TzQ
TtQn5+2hZ2eiS/wZ1r5Jcf1DvRt43qvNXGrkhxnSY2BJWkhLgumQpK8KijtliXAK
ev1M47uTozQpvpfTlsFhR1a1iQGrW7HtpUtEbQw4eSXc7uqSZ1xePCYexJeWY3Q3
am8dAszr1sYaFi/MOO9iV9X1XHlg8tDV8/HX+eZPXvVMEPVh97bkchce2QXzM0iI
dCkUYHr9oFRo0Jg/Bw6xM7fOLNSmZHKqCt7RoqY8WpCOdDlJnnthdbEmwxzR2WOX
PnijU7ohi0Nug1djp9RxN4Y6jmC9AYqoQspXTZkcOXEC2vyO1/BZA8JK8TF19mfO
8N3gO88IW9f5jNlLWRcQl3kb4HAeTLirSlRU22DfsbpmPFQmzKk71u/EpJrJJ8/f
bxRXwza83fJbvhyuFu2GXhOkJ1kvaeqwpadr8j6DtSkESff0No7aS2UJGyNR1Swk
RAOIN/s2APGVNoSMX5FWpT1KH85iTonYIgJJksJXm0ElTngieMlbdAgjVRPp8RPE
UADrKmkXg0fe8+/jTdzbn+hccfnt87fiSo6XKESHh7lKohlLdGMR+i7giEijdTjc
mhqkXi5LI+39t+EH82JmwNi6hDGgdUtgVWtMyrndY+TizYx/H4mMPxZpcd0SVgom
QCbQSvORiSsyyGrIEkJSBbnOiuT54vdsWU7LV8FLGCmw8heQx4KFc8vEs5gCRwyF
ByM5Kl/wRhv97+1mcDR1Plw27oqUwjxkwGdtDgST6YqMrD1Pm/3EZ7ONz9VMOG+h
j5JysHAwavbqgv9OPHt+RkU1Tr2kPoTHStf6pi/oQ5wDYNcQ0o9HT59iaLFwDQ7U
cRj6mLngUXjO4WduXlEDL3j9zeR8YeOTuUaO6OgswsRB57zMToL2F9tRbx2NPt8p
8qSolwyWTO4zxxJLTsd8pBWe70swkE+WTJX2vkoN+7fmPxznS/IjUTxUHlVULcqy
0BDlKBXnstLnPXIUGGYPvn+hGUKB7VvGHqtcCXGCAS0prGBjJ9dc0Ah/wccwRLfl
ZJig5zZ6iG1val2XXeCr81OWBBi4sfJV9OMQJxJbOT6WDRio9j8CIs2lzsC2tlUi
VPs95JPfYpKfFi2P+PlpcsDQRDaMp11ktDLH2tk6ikHYcAEigIpOEIP1WZ2UnM7c
Xd5Kc8MZuWuv12C9WcH1Cs/20zSbUf09yW7xjSiSnmWS4tyPFOCPi5B2Mq0NLJyF
ehyKnH4aLR42HnPi8X9e1P85AEh5jNH/evPnf9uyVWyBUuPE0cheoD9it5GS6nRF
EhKW+5xAQ71PKRXhZt5uHlaJm9DellJWUUBxBGNwykFz2Pdru6WFptah3PuShli/
YY6+n3bij1b6l8kq41gSY9ctG2xmm7yYbOqTwC0dLAfXj8Rr1eHN1G81KCUrpnSy
wMOZi+kI/HZKfdcErk7N/NmG8J2sE0yzDxzJkxu2bnPD+GDFfSAIOhsdNmPC04Ts
jTAVzLvtFTEYOPdgjCA2YyiQJts05VVJp+D+z5Z2i5iWUfkWdRN2PvleAudze97H
dC5OhnjlM4armjHc6iZgQYqGsKP8lk7WX1h0oOeF6vxI5DNmEcCwcekEnhdwVMyV
`pragma protect end_protected

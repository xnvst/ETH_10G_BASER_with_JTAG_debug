��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO�����l��X���e�~ͅ� ���!L����1n 0����t�<e�I)WƸ׮1�����,�>�u�G��eE��X5�-���4�_í�z���H��Ezߤj|)�J6�����=�{�s��Y������� �u�pA�g���k�C���o�|�}�f�������,�O�V3����;w��28����{�F^���������Afm�y"��&����h��T���M,�N4�����Q���g�Բ~b�J�nKf�Ȧw
�Q��+�ڻ���P#�n�vr<���g����F'\�
����M����7.�"��5ȼ���v���y�\�����rYN�r�V.��=��Z�H���.%{kF%�qR@�	<��y�ف݋����d�:�W6�Rs�y�Xh�hӪ,����ΫUw��ޜ_t�/Q��=�am���ܾ:;�����o���l@�Z}mU��Q� 2J͂��<;� hb�I7��lf�D]@���U���ҋJ]�d�t��rG/�;?ޫ�uS��5�6_�Y�q� �X{l��o�KN
�#����_��r�ʵ5�iӰ#�|u%9��a�e�� �<�pۘ���v��$��h#��Tf0��z bL���ޖ]A��1Fx#��b�e�N=�U;c����cj�X��u
	J��CW�:ux=r���V7 �V��r��{�'�u�/�h����� ���⽕P�P�e��	�`��_n���qP��P�%�V�Ί��\B��Ķ���Ϟ�$����bP���i��U�*}0Z�x�yHEM=��a��)��������'��h&�Kւx�D�Ǵ�F��K
�<#=N��MYo�Ӹ���۫:ӲRu&Ȏ�����7��b�G뜯`��F��S�:/�;N�F�&^ �|z$�r�b
�-�ڸ[ŝ��5㧧y�?B�E�$��ڽ4n<p��y�M��4.9��\os`I���g�g�Q1�<jy�U�xX�*S�F.�K��SV�@�6�0y<1�w���f�/(��?pm�H�FS�d��tޝ3��a/V����
?��%���MP;+K��JSB��Gá����Lϸ�^Yu9ur�:j�LO�c=�Vд�px�%]���Ti@j%�?�8�׊AlFXo��Az�$v�����L�K2�甡�oo���|��o�#A�� �l�)݊chf�ނ_	;� ��J>���[m���ʬ�7I��tm�F��*�hrvn��txV��:m��;���O�z,}��j:;IY��ڛF���U*�8�t�^�]��׹yO�_��6��IC��e-}!�1�����:�6�����G�Θ�׹WAF�w]����m�[�g7~�B�Z�3��n5��RX�)z�֏ْV��Nz��3]s�\���]*��V����J�#!�%� ,SPi2=�q��a��%����!�M�\Ζ!uLZ�jL��Un��qUG>�c�$�}p\�`:�Y��1!�^I�Sj! nSQk��`�h��W�����CJr���漒��}�՝�����J���\���Nf�� K�<*�G�mKv-}�����U�2!�^iC���x����5�r��E���$����X�Gu��MU�YE~0�1^���X1��F"�o����S�-݄\�J�w�hւ�"�󯧱�Q�I�M̻�?��W�P_�p܋���'5z�i��E����7|o|�tj!]����T�틆��x<lؐ�	��0O�Qm>���<�9[v�-6?�ˈj1��& �y��z���U��ԩ�������V+�A%����tUUg�;�k 39_�=�	+�]�#���ڧ�,�F���ӹ�_ 	#�M^�+|ނ}�9:Sҟ<f�KYg��H��&�wm�S�.��+�s�u�s`H�aD���d�u��>\l/�5��wZ-^�}��ބ�@v�;A0�2��Z+DwF"�BT4�����,��;�>��/l̾d���_�	Qp��4βf�HZ3h;���߆h,��p��J| jf��`}#��pm�Έ&�$��̩h�\��&A>!ccN-�ݵ�/��ǁ5��C=�^_��M�+���#��Ҍ����_�n*HR��kY9eZ�D�Hk�	���{�ζ�>í?t�P���'ʍ�����Y��h���?��J�ʻ�Z���3�o�ӵ�ХL��1�okz� /���P>j��I���
��.���'Y��M�@��[�{�?�e�X�\>d'����vV���2��*'�y~㾱��
��5F�M��'t[ށl���n^��4�-�ڵ$����1����Q��}�׻���<���ٔ�)�x!Tu��#��/��Y�rU�M�V	No��XE�a�wI�������~����a���0.�)@\ �����<-v��ڼ��"L�y#@�C�Ξ�Ne��Xb��M����Ae�짲��U8�Uldhk{�#�)��v�!�H
��&<��=s��U$�U��veÔN��NX�X������3�AAN�����ƣ3�}�S�l��wAD��n5�+�O6}KN����ݐ�x�`���gZ�	��ʯ�1�$��ء�l�~�I��0XX��u�[��4�3�ϴW��E�>V�zo]&2�OFC�$�Y�&^% �����>ܬ'�QgWZ��xt`=P7��EJ��xI�J��2�E4�	 A\�X�f&�7�R����믡ۣumpt���DJ��!* {��-���
� <ZG�n\����Э�Q�:�`P�l,Uz��vr4���:�'2(n���F��c؍���,_�G�B�O_�W�����>
��P��(���?F6&h�K�6����7�17m���m��$�,����"'Uk��&0��&M ^��&`ˠO��f����˒sIqT;B����$͑`G5BI�(�EɅG
����ګ���LP��b:פ�J�NЗHF�bG�TT��E�"^�h�QsR�'���A�4$� ?Z�R�V�5����#v���}���f���q?�y�U����θ r�����@�g�B[���-��7�_WT� A��7�
g>��tO���ڑ����}��ʇh�Cq��,����R^�m�ƴd���'d�&z0sMS� �m��<��Է�f}#
g	t�2'��g�����*xDc��l���C����	�Z��J=��㥪]ZJ�Y�䰔�������$7�''���X�Jo%����5�	U�p����^N�Y$��=A-}ī}�����PgF�Wc@ ����F��aS��F�ϸ���+���/�^�#�b���_�G+��-T��҉7>��z�|'���6JHhQ;��g)�Ձ��]7�l���B��^��M縝X�w�7����٢n����s8jXG��Gk���J0:�J�J�7�?s�G������W�E.S5#�ֻY��T%��L�-�T>�s�V8��A�-8��̩�#�F�MI	sM 3�8N��.���dJ��u�:��4k%Ix��ޟ��H���ټ�}�Ԡ�wNB�S���>3�3���P���N�I���5��)��#��A���ioeC~k���pt��f#��?�F6T�,;��o	T��s�b��x��*戂��^mt�=	V�X�[R[X�p���;qB{]ojD���G��n�K�PtBNEp�o�kcl����a�:�Et��������W�>Zlo6��x�N?f鐃P�}�Q��j���l���آgdX���kz
�3����m��;�d_D��驽����1�q8��K���U��l�5*+��Dl�D. �Tv�o�p��� ��y�^�R��lU�Y�Z@��� ,Wh�H��w�ٱs.�ByJ��듙�k.�'l2COv�JRI�"|E��SZ\�+^@�QG�^�ϰ�]��k�b���h��j/����3�)���W�U1;�_˞���N�{���%�52b֮+�Bt�C�~��U86�rD%���_ց���zq֏����P7k��솠�z�Jp)�6a�L]�2���m��Cbwkʹ���R�suD�����']���i�vn�Ғ��i5 	((/���zI?��N>/]W�ނ���اIF�SE��������G��RηY�sI�����!zУ�z�y��j�0�w%Py�MC�ʶ��Ȼʗ��JCp�DI��.�[�}އ&&^��9�ߏRw�y�~9�	mh��N��+���Ʌ��}���S��b}����_6��d9v�5re:�.�f �wජdL݇rZ3�\�ZW�c��ڟ�& �(v����ef�uT�#Ā�M�i!�8 h@�گ� \|!� ~�pQ�,-d�4��g	���댥)W�7�ӈ$5P�s9+�+6���a�� 0��?鿃�A��_�qx��b�y+hc�rZ�� �m�,Ӗ��_R�v3p!��!� E���w��d��y.4�e} ���y���L^��(�u .oL3
W�	���^�O���,"�c�1�>p_�OzuVs q������a�4�J���MP�j�O��!ف
�L&��L�u9N/�:P�ˁ��D>0��uf@F~|F�Q �<LH6�;��|d	�t�L��9�DjN;�Gh�6
=F�9�Qj�0���*l5�b���XQ�_USx�t*�^�u6s?�@wr��zp�ᆦ�w��m��o���w:���svmC��m�?F5��|�v���7�+�*�0h-�P��/�K����.b>���O=-$�P}��#����In�~��b�"�G��&�-N�)xTJ����;�O�82ie�%^ܙ�x:z��p|:"p��cP*�`C�+ϩ��mp�2K2��DRμ���Bέ'�g�g��?�$jv\<J���7�f"�G�L̦]J3ɕ��V��/M�׮�:.������gL@��U��V���d?8�q\y�3��焪*�k�MJ�P�e=Z�mk5W�1�'��Xo�%W���>vQW0*~���_W)�!G�N��A��!Wd�G"( ���~OR.�Ӧ)`�[}`��䈾p�iD��/ށ�O0�x�(+ƣf"�T_	��w�L�d3B�K@��/��9ELq��G'�OjV��ǈ�,��mavhY&�=�E���k��,�W9���(��W�ˋ��|c�k"����[���S&���6���i����9,� &	��wܚ� q1��o�Lﮞ*��a۫�
Q��Sd�`�PK������<Nll�i���_�T��e��;����+��	؋�[!�wJ	���c�� ?�H��|��t#w=�)��u�7��?�zLnD�6
��4q�aT(��g��E'��z��!H.��DE�j�ɧe_60u�UB��*�ݾ��:�+<>�u5ĉ���'B��Q����}���?<��[��o�}��x���o�'�ݗ������m��ɨFY�/��4o]�K� !\Z،,�'DP�A�x�tV�1�������/��0�����/��k� ��0�=�2����G
0����f[���>�D�E�"8�k؁h�&c	^H?�C�� ���Js�����M��Ԏ�{�k���[�h�Ǣ�S?��Xދ^�Mpe5��,g7JT�M�B?Z�%H���O©;�&hX1� �89}Dh�t�K�c�x�j} =>9ϣ�9X*Ti[@�<���d{e2훬uQ�c�(���/�����.NB�'v��ozT�/o�ʨ������=�����s+i�ke���:5��0�{^o�O��#�qeF�b�u�PL���:���������R�q��8d���%C�-7_�-���c>�[c��?)��lK���9i��f��\KH�L�f�E�˳������vf>��ʿk��Ĉ��H׼�_��m�f&����<i�A�a�[�|�S/���2gP�	���y�fjO�����8����q_�K�/5.�:�j�A�B6Ԁ "O}g�KI�k�\޽�T���f����]��ь��ˢ/�!5(�/�k ;��Q���%ul���f�򜩌��v'ּ��H�����_��cW�U����G��;9�j1�{�T���Ε�\�My:M@���Aˁx�G}IʑA�8����+���Lh�7Q,x=�Z�l�*>V��D��u?�Y�R���r�.�e?8]���)��h�m�I���~H��{hMZ@Dq}�ʕ�������*[�S�4>�bH����j(��Y��z@� ��� ����c��d��!5�T�T�o�x�	"��[i�]Ί�f�P}�C��V����'HBxf�%eF��.o)(��C�,jTMuj/�,�B,q��AP����}��7�x5�9��sq4�a����m�WY���8Ģ-�z0 ��͂�ܱ���Ekdj��{�`��Y��P���Rbc��/����T�b��&����]��޳�Y��������͔�T�6�>YЫ�����*i����Ø���5A�/|��8�IЗ��	�	F1�\����Wu(���K<�[��n������_%#ke��kL����h��C���6�B��p�Z2����X���O5���5.�Ά�? �ܻc��)��Y��M�i�����L]��*�,��Yt�;���Q�#���%�[Ѧ�������M4�N�h���^�4@MpF��!�>�(��s�����Z}�UW�P(<��vu�
�}��.wJ��Z1�\S�pS�,�SŜ�����E�_�OP�y���R��h�YY�.���ʾ��*���5õ�
w�/�Cʼ,-S�9e���ɜ�ay�=?�q��}��M��s��-��zR��~߰9�I��M�_)���e"�O�&�n�`��
ƷqL_�H�/�~��B�{�e�o}>NX_����L��Z[���`��E�v�-��v�[�?������N�3��p��{���˄�Y�sx~��˟Y궪k�U�h�T*g���i��w�O��[��k�4n�l������!�����.��h��!9��*V�Z��i�����7�G�q��#��[��t��@{���jbp9���_1��hO����ӱ��$�+�^G��K�ӣ�W������!��4{(V�yiP��C}Ƽ��EmX�64@M�t�s��
5�M��\����]�ɢ���'�hKj�+4*���^�DV���=�~���!�ԗ-����ݡ~3޶x�걚����Q�t�5NR`�Ws�`+�n�R��uU'�&�tiާ���i�����e��b���YBx4���]�4���?�b�"��^&� B;�rO�,��Ѣɶv�E[K���WF�ޅLw��Z���������/�k2���w�5>g���}�L��O�	��M��Y3~��\зȠQ��!��zP�<[�����H��b�<��k{j��U$�F��Y,�gv|=sY��ܬn��ǄP���۾��{�r矷7D|��1'�
// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:34 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rwJmoqmNebIjIh7/ZBOxV+VlPYooIHS2L/W8gw5fjbLl8Jkger8LgcA9WJ7HYMN8
O49vv2YDjpthlfbfSVPmm5XKO5cO0WrWNhcLwdKI1R0XgXdJw/xOb9zZ7N1gGwa5
QqC0a7V2t2hxxRlrrZFri6Gwba8zheZpd+g3fn4iROs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2480)
qLBokOpuJNcaVaxxaL+og9oNeZIHMCZwxeVnb4IfrbIkxWwI+FdZxPbhVcalak/A
7XJ+hcXPAiTOlRQ/a//yayDnHCof6ECKREuHpM4IGI2XiKkAqcMaXETvOU/HEsX+
adEREuoxue+rK2kXhOylstpso8cyMtjcwBZaxS1h4afwHE/eE5kBHY8EFyTWYM4q
YlGMgItBFetIhfoGycfOdTi3+umLwQieLpqJUMDSgYxNc/yTveUzgbsPAwnQN6kf
v0UzprkLtswVTE/WbI7yBGn1ld/xYU5OxM9mdiYUIUbLoFmp7db8Uexlf7ISxsrc
PoBG0ssiAtyt9h5WYMYfICvA8V0NkvczR+wiyGLnru6vSi1HkIgupfWqgY+AvCJV
PV1SEdWtw+bNlOHEaUzpKAUyoisNS7ji3TJN+FMhTYJ6zTDcQ1feTEbGc2iwmI1r
joMoFhxvBkXEReQ/Y9m1CnYvuSulj8Zs4Q5vr3kKJCym3PtBsmatZ8hEPn3fRlJU
pLNAcVUJvm1e712ML6NJfvYWu0L4YmbnKIDESOgkZE1rRfDnvmfX4N8GepEJXewV
ymEUcXliB8YCdrD/+rBCns6HbWTChwxZl3P0KvAhhJxo7dFeqMBSMa8PeKg9Tvxv
jbISZb6T/uZE7JHEGrcgYIiv9TC+Ts8aZxvT515xD8FBuGE+GmFXBqVoDeyc6TNP
u7wiaerLYMj72Gpn5xjot9tS6zsGcAZMWwad2hXR+n7s0DTLFnxBfQlxvcxDBXP2
675HbGZ8DY3xgHTlC/PHfyuy7ZiH5yOaG+eohX9o20qgRdk+ujyiQTK4bnwi0hi4
6+cYGQ9//ynchutb7v91DuD3J7TnFN6PfNTA13yL2cozf1RdSw0jgNuFJxU4uJxI
RZcLRJ0F/C9eF56YMcP4mMUpCPdcxOHMSeicOYfDck0bpXz9g/C1jDTFpEXiJ/0a
vPmHu6VNRnBF2MfuakZaUeU/PMoDTYyOKG2rJgawqTAhZB5kP5iCxgsW3j3UHnC9
TBFnX4CVKJqfAEMr+ZYrtrIf89SJQYr2Wgfqx7BuCF+kV8t1304InTyNcb0v271m
QlKWWfoJg5rFV8pM8IaQRdG1xBAtYjHjwQlCXWKQmeHpymmAYBtR8YvtMqVlbbDJ
OoKIWw5+E7H8iD/I3CDq42IExr58Hs4NxBpjyzFVROQJ0+C/aqy2dotHY9m4K8y1
ihtIshNQDFZkd8si4cwuX4ju76Ezhp2n1c60AUjaZU8/Ni2Hnt3X52C8acxIjjI0
nN+6Ba0XpYrL8t3vuJ1T/tsGzvfv9+GcA5pzouFq/XYag5mUYzTBPdkU2mBEbgRX
5DowQNMQJy67VDAD1PpX2Ym6w8NiWwA+BWJgA0/1g3MFvb3DYQulh3II4nZVITpV
EL1nFlEsDUPfrg1dLW9kr4WZZvhMFmPiSUyEl6HKUMpECttOQUwSvWpTpNU+F9K2
gIJ942sTF1eYYMa3oeD4GajdrXgYdvNL70/F6MZXHjykQtXUw/Z4WsNkFkKcUKEp
biEINpq8ZQrNwN+5Snngw/x84jBq1PD2jjBgxWhdnnVgjL3KsIcWG49baPdUv43Y
D0GgbLtSWMpjDnmuRhz4W1kLGTY8pUts+qqGNLsqVFinhc6vXe2AHbLnL/yF5vKy
vBphvvnnRcfQHqR2FPtnAHYNE+KhwIaUX+LvraH+XvHExF16Ar4AhAfA42geuJDs
z6d2C7OAZxc1GLfJ5ige3XKRACf2WAZwAOFXNkqlyqT8qtdOUd5LojC4UW2nXGlL
88D+vWDAYP4Ho0vpu/klBFthBDZ4xoowKydptmeRyh3ShmQ5CSK/cWWJRR/ncM5w
t1Ns9hPKDB43g7wDO338qNQ1CtKPouLMLKJHuGPogfHuSRzllfLTFRMhhuGPOhfX
VUalzQnTZWQ9KVT9DEnpptjvj5IH/Z2G0sAsXhDTLMCGsPvRLp9PkmO9x+yOMuWW
3ASAKTxqOeP3rxymP4tezYDadMi/s5krWv1/FFOqfDqsUGXWgR7vKR7zdIgnOeSE
kz5cGh5juxyzMeN0r94Keob9lXIYYT6+fDGai9JPyFjOQkLILkW3xr3rFEfra9to
jNyecq5ZkK1w9xTOORE1aHuAd2EFDY7vl6hS24qjawvxUu10lathamF4ByJUGlmy
bOjeFShOW/xh2FLHs88n7IngLuxSPx5Aq3liqmFTSoj2tJWpfk/Oa2IBQydnCNWY
9DldYxeIiJL+Z9H7wMBM0dhI4NtMVvxFU1L4YSK1OXK9RbgFUPC8j6fr24dSq/rp
Ws01JFdsoHpmhgj0SjLihVALmJjQlNem2s5BdDoTjkYZO3GGp1NJ/1SGR4drnGJ+
rmQvnsGU25hFhSfKAO4RDGBs7lGT886BPxJw973pw85AzmpFFjHzs8MUe59EEpfF
d21TtzK+jcX1MsyI7LyDTWaQgZ6vviieRkRiZ7bFKrd3F9Je7QyvrXBDfErdqAkI
C2SyOy9lXnjDXac7nPi2ZdnHDp1Af1UlF9mNiOgtL8b95NPS0QeGSfw2H6olB4SP
u7sZLh/xHHIuHqlTMnMgA/6vKiZdNjmcCgQ0L8YK8Zx5Yg99Nqm5CvottvW4sk9c
VKTHhWKsTb1kO042uqiUBpBj3tIO9t8Pc1JFDMHrCvekMiWKInu/RUggxrNMBKb2
NDfAh7EPK2r1VSWDBdqt9Ii+tmFdYDhJZUiIw8vHuLJqjaUzcRRLZv80IA0cIn48
l4QXLp7/y/0XibohrU6ysUy4A49+1hrVSkSK+8ABG9tvvQmwLvzDmix5xxxTNJ4s
/DvOu5kr2q6DpZmpNAcp/smS4psE4vIZyO3Ncgi/ZGarKo8mGusgsGW0wX9xqZod
uIR4zQQteEKEwWtz6nqzAC4scjtscecYyZD+beACcOHcSSkJIvvi8YQ1B0vbIIyM
gXYsUpZlQih5+cs6Svi1g94hr+VuZ0m9UzU0d8DBnCvZf/FpNmTuxtFly2LBZSQO
gnvs1zQ/f/+hj57IbMCn76LAOV6HjtcRiMDwynYOocFTXMyM37NYjHFqvNsSz3Hk
cVsx1WaaFeEzM9XeU6PbA2O10sW1V/LcRB4K7eZeHcD8yGKO09uXq52IoCcjG9kE
+Xvut8iGRMqGXhSFWE6O5sfGqi4Dxr68od2mP80heSj6RRAxRlPQJvZPQbVwsl7c
eCgYEdvTnUk7F77UoyUSDWHm1aG2PKRebKxJGe+rNV3sJIDZnCj+nE/jx4NcKGji
c8e4/m0Qhxd+mzvcqpfi+4KO7jb1Y/PlYGqjiUYoN1E=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:22:32 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NMmpvXWe+qFECABZXl/Csv1D1YA1/kZx5X1cnM8WmuIK9Gned1h113ZzgBFut/KB
iHrpeQhumSoC36NufdwAQVPCuB3WpH7XRMHBs8oi/7fe2d4q+LnRVHciiigwXeaM
lsM84U2BoIDF5guQ4sPmBtV5rthHgfrKvER6dx+3fQA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20176)
X0f1gMtM64hug9+rtU6r+VxDuEsS3RfBJ2yC+atX8z2tlpnKyAlgvfCPVj8zLV5P
Xt6mIs5XujHdEdyCb/TOwowFn5pyXa/LU35eAZUVkuQBpdDIGYeMrwsUTf+f8pr1
nzoWh4UsczSIbgEWVbEQBdp76AuURa7VCfMa6kkdqS9/zDf9H7Rx5SssPKOims1Z
MQh2mXOpSupOzdZUqgEbUEMNIbRvq5ng0c+6K7ie9wCVrxb4XyWI8r/bMvXXbpVC
uJ/ian1Jgj/a434kBr2mb2V2mk63m5guqERP25PbkWLCQxzQPWmwTslFiy93ggjm
cf52E9nbqHxM7fI0arowE7BmXE3QuFJnIWEuDNKBRJhceK8vs+dNitlDI2CNw32c
ZAl9OnA6lpjtcPzrqjDRC+KHS/TABBLKUHkJNwJ3IFYMCc5DKe3jtHXnUugr7IuG
jqYzXLpWtjipYKpEr+aT6genZB/N85ROmDEWLosYHaqIHiG25jbZ1elcou6jNERg
8StNid3lshNtoNcksiogQjYCCz4cpO6q3bNJ2mD3mJG0B3HIHmr35aRMuKBI9JLX
v3h8DHVJDUzTZ8Mgq7Kwi3vTbRXw+NvieUk7eccFOjKpoTLlRcNybqOZwsMfDfOc
KEREqo3M60GhhChlhrAs75mBOThByg9nJDXevw59fi4MKYRXMpguSs3eH6YHPeKv
PQgnqYot56wL9Ru1XLbjRPhN4uR9EhaTXPnHU50qUwm9HTbBNZvf0g4k33Zll+6R
jJSbmsXY1UtM8WizsiW6P7K9XuZdc1zOYxfZlvEJxNhv4wnGIWH6mh2G2EaRHGaK
lIpkR1wEEQsLu6fD5gBiwWFLmJW461HiGD0DL9/AAsI5McT/arPvhB2JWE020U/3
ZWNCcAfCU/WN+WXSDxQShG7w9xmS/bz3ppz3+dYXBSOxzpZqvMt9bF9j9rSU7T7J
SFrmwcWbWHzDkLDvHv5TSGZbkwCPOxo4S0W1CqcN59MV1k2p4xP3tpeKwa6CiNHg
i43QHBkE7VT77FbxRQ8RK/MTO9ZVnxhQwsxu6LiGrNt9qGvdjKWS25cVb8klejsG
hqJ4KEuZgWT3Yqc73xucvy3/xMxnsnJD+yHkZ15KPkPzwxuOobe770y0WUPeMJIx
+gj0VFcY6lYcUVs0SQXOHWslQS7FbjfPzq/Z5XF6MQjVy9nlDrNgQtiwB6KWjFcT
Yvs7mHHfNxtfkBy1FO7jmifhCtTB60HbzyFz6Kgh154n5gjk/p6rckwZ6PY4OLML
5YXyYsXZX9Nj60EIz4CcY9htf+LaQP34rEWDhjuPaMoJu2O/vCeKR+eQLPx0c2ZH
vO2PRKdD1fPaPrUhQW0JmPzbqL074nltfXnnYjo7mOtfqICaY/B8gc9aVTVWsTEo
BNKEBxmAXjtxm49P34bKz74AELAO0wWPcEWRHM01mJaP3J9gLqxMzxxMmeioxKUS
6GMK5my59xjeJCIOE68k8gg1yleV6a5uQ4qTq/U0fL7XuPi69vruqp07/nolj63V
6B6y6PMEI+SSTZDgzop/LWhh2xmeqpT5E5bPptdHXz33ZQP4p8rXtcZE1HSoSNdn
GMTlgfo0ws7ckAEBdvf2Ic9zuP3cC7IcWKk3bYljh6OWQZUcYHgwIuSVbK92nzyD
3vpy8e0c4s0FTMhXThPgiwouFrALmisv/KMt0O5wI8AyHexHf/4nknD1s0VLaKzF
U3yKBd0Lnjra76UBtQZxMH9MtWQ7XYXm4odgTSluqTlbGOfQx/GiIy1j++Z/YTNJ
+mUWt4fKFYN6q93P5+8BiQFsLCaX4QIEEpgJilWKbgYVDrbE1IMHVZvBHcqzeI12
3Lxj6Zz089AcdK+FJLfLoxHJzhoioK7n3AnEzH+IR/zelrEENAZg3elOlCt1cR0x
6O0sPqnHeDI+oAoup30WsUOqtAjSLGWPeq47Zs7yV4n8uIArjmPT+k3TpmFjSykM
xjQo0Dg86Ti74/6u9ZoUq+KpnMBwpgUmiZVwJLNkouDjuk4TYfhs5+BlPZt4h5mD
lcgQ8st5ueMzwKbzbz2EuoOsQDoStk3XVhqAB+ZzxcDu1SVoReRYU/7SIkSKfqh8
URxVl2pr/ku5+2TQeR68sMwJJdq+EKjKDPZ0D1z8tIjrzPid25Qtpn8FMCVp507q
Al4h/APBmlQgqQ+9zpZJVyJhgZxZdPRVT2tQqev2hZXV1V9sWTcc6unXQwVLlLl6
DCkzzzeByPEfriHUWchICeLKU41eyvGK5KO1modftwpIU8rgJOH1xu7XvH71iwe/
J481SAuEXZ0nlpn12whc0VjQY1L5b2GLTHDD4vp6i54231yesmqdN3iEHr4fdwQ5
WbrUmK7fBLlasegpC6dgUmKi7+e5ekwin0kUFOvVrk1fJbFCOf9EZOoEb8EYovd9
5Q09kiFaUviaKlSaPKIuK6ozsSxRYtZS6rVRR+ESYKr/SOp/0pzlDB6X4iUInBCm
KMHwRMYmYLxW5ZmXgnY1XZ8MZj2UJhv6hL3RdDuR0iqHI2WuolUwg+Q1HJ5AQ+fB
qO05hTwrT8qgksaRyRTG06Hok1+RsCfyF7dUaVqkFFFINZWNDbAQLqm1yZnjxR0A
J92QspQhSMVBZrmo+skqM5RrQnjG8U73Bk+3z3G0lq3lKsGMPtQuf0hcRcHQYO+V
qIrQDfhWqS+We9WOta6LB469i+t/TNIZhSKUcGFtCvR6Gd+HetDjAf5YwcjRo1Og
HfBNWaFkRzaDHsmAkLpW5ueSUumaaDqtYP9/9sOGcDXhiVo/LCYjxyfH4wY9qfyn
pfSZ+EV1YVLde1lXgtujkGid/eaNO/bE28XA37tWi6n2ZrL7OEtABbCzEzkrdn9B
9JcaKEvKH0fWzdk4AoOoD8lS2B52ymg+DK07ysU1LsVCj/wFDQ1Z9zVHy4MmSWWX
yy+/9z4XZB4Cjioma+73ZOz7dNwFLmJAtV5Vqj0MCNthaDcVnJr+Y6M3FSJx8/MM
LrevJ6aeqmqe1ySH9igGGTqAcYFr9aeiyI1PmWdIj57Q/esmCD2sFIRjJFprn4uV
IFPtjg8X2yVMkfWsmoFV1GPweu+3OMU0avDp53MFN0Jev5YYWwfRBYyX51lnZdzX
s2ESBzqMmoo/FgogIgq7IQ36jqkmjilCqbtrXAR3q/t13QwbST8gK4tLnar5slCg
Pojzl4c4EgdMwVdjkqH21vIP9n/wLlyW9u7bZUlbOd0OPvn9cZHrLImcET518lyv
J0sisUsOKNJC6EwW/44LaUF3iRjs5kYsCi7hYm+H5pdrKLX9+PEX7AglQ08mRnWw
c/C2a9e4PfVZFVoM0TSYW1KNIQjYIajI94ZG8eJlQwPuTy6hlzRo7tamta3hfDJ1
ZNS5olrlpyvGR/6KRNakZ0QBVzcc8jmdYnJibEG4zskC4MHK6kRBGL7spNweKI2N
BMyrSbY60ds2LaAD8hOSvs0h7g4B9PpsTYfk7W26j3jzqVJZxaGmS1OOcamFOMde
8P0FJdMe6eaL3wrprR3urRjs/7pQW0E6pE+lHYrVRG/58/XCxeniufCrp4ClxeME
ed/SnML3ysBPZmB4QdtLRPZhXi/a9Eg27KOG5+96IRq3o6LkSXEEfO+OTuE6WX5g
uasoDh6sMDgTNHOZhvKiRxsS/8ApUhGJmGmnrECP9+9I6LA+QKQdpKQtdbVjhr6s
R74qHZYcAEJ+3jwKfIaoukfGuf8r6+JC7bP48dMkxQf48mesaLegy4B/+MBiAgD1
yqSW6Q/nmMLDEhYvIdCFpcx3wOSyBOBJOID9OwoPftdBZtpRioc9VwbseK++gX9F
/IZJX0i4g7rIduKnVmKdxnEdra0SCiS96HU1BjUZM2MKuf4cBYsvhIcb6iuuWit0
bu+OuhtDuT9FN6wwYsaBuhS8ey6Dr8Ic6hpG7bKaGjgCqIX+KihVjfXGKVn7S+Ai
HhgM/t4FJoly6qPmOYjN8ztLhaasiYo7l/ABZzAzXGlYCXOVauYbWa+lgmrrvKiN
pmtdavht2MDtzX697j76EQ7NVqPgvMnQWM5mZTSudKyV2gIzpQ8NEs/Jv2XY/msT
cUdrOVDfPaXNABkZuflJT9qLTOZ778wTPkVnk0SWmToF+y1dYU0e9GrkGEhmTgc1
27JD+7NLukLiqv5bngFuRmBcP1LqeN2X9mC/6Kzv9Nmo6gDNmVWrH0WwULje2dgL
9iKg2mpu/frePKuRDXxbRsJjOELj42MYuf707sxe8SBGjvpFHMspBAFUsjEgNR4L
SV5PQWsBvRViNTsB9FgqDynF0v3OXSes1CxYc3DSOkY/46dYM+MLtY8kndWjfNwp
YCWaT96013ZuyNUSWJWt0E0o30CT7n/qutuHak35zAxBi2bvQ1jY9jeNSr4i64Ib
lHKEwYhqO2ES2m8tPayESrA+vCS9ZYZw4jAuxD912vLFaz9TVqN5vNMFe3MzZdLy
FV2FlPdNnXV4PLE7i1LBohgWON1XzDC4OBigbDN2cDdc5KO7COiMkZ89zVuwRQTf
wQu8MTCtCvjB4QC5OLwp4dpTE7ZiA6mwbXkllAUNKtdnrJeP3kD9VKIIsNGVVNuH
/053tyPG/W9RiprOIqvvYP3qDpwUuNsfMidmH3F5QJ1rhTNGbfA1LqbYWhfuj/3r
1I+AY2TvCHoSaW66ID50ex7I+XklsMNkdftPvM03VbyZ+7Yp1lu5MA0b9WfL7h+5
dTigUaGAWGX35etZxJQFwwXbXf3dry41tYKSgiD4OzXN6cezm4IDH8gyFXBbNOsW
6VOeopMNvUtzhUrPk1gRh4POADQYmiC4GBGijQenngpfyiyWY2y5TaoDf0V5wipi
hHDWPyLDvqyOkNJhQGFps7S89GgsP/KsGq6PJyWYzesg37uJ2n+UOA0Xgzp5ya6o
81x516bz0bEmPy/2pqTCDN9WAux8SJ+DC3LYdF+tjf+3114+5LNHXZEMlSHtbHbo
UwyRAsuBEvZo+TE6Fw86KMbJyhrX+JZHwYCWL05UQR/tLGJqHI0XoxdH1VOEElf8
L7NPLXtF956snZuCOq+TFMyL4smWZ+brYPeiEK3apciqcXkGI2u4PB4lXSlV5Ipt
FuUegKyg6fY/wcc02zFgMoo4QhpvqXTKwpGy1cavZDA78vcZEAPwPPio15pq5bs3
USGfvSuvOf3GiO/kXuMPvaIosntdSjB49uflPpKCyCfpo9UeVOgj80VftKOoB+WK
iPzi1w6vbg/ClIb5Pco6ixL+hif4Z+mPfF6zlvJ0lPlXxPqKMECK6/DXn+PoAucq
oXvdEtc8q+H0XN/IqKGw33J+q/ATtYJp/qRijEbdSv2ox1G+5YTIhkc/rJimWWWA
wvAY/jIHbHRoflh+LeIOo+Mi4XhAM0yThVM5sKgyGorrfOef6bZ6DI4e+GllUB4H
Qgc6X4LwfCKYM8h/gowjAJ6WxM+uq7g8Ub93znViFQvLXYGGG526uEvKmQQGz3XM
z3V1kptkI3vzKEzhRpKLYezd83lKCv0U5eoSyE9Xndq157FYXlrCb6Pl9QTeO8O9
3CgBxnePfpvkDuof76RocCv9N7alNQDhCS6gYAR4tWqT/j5halZ5UOsk2X1ggQLF
oAVFen0P25PUtmJxYlM19ytIMvo6CSDQrIgQSih7m36D4rSx8SukFkP7CZKhl1f8
C+D6B/r+hTCsnDXJwaujxSTtkNrdGsLNx143SApirU3nygWufHxUHwzv39gngruk
CdjIEq7cwzHdSuSusCyJScfWEwaJZc4llJYJnhJY7UyhDDudyaJhBR/gE6SdQmjw
SJsJzOqQ4CQ4DkqBrVldJA18jZXP5ZnqGGFbiNAecEsekpNlFDN+LWRrzGj+p9DR
3qcqx+AvBsnzMgQM2y0jhmvT8JcmjBu6xrrxFip3D3GvESpL+Y3wX/MqexzZdmlW
GAYeqfH4TSOh1ohV1MVyXNHf3dAw4UmFtF6T6E3RWdy+EK66XqxXjjIsMPy1jtqS
kx6sdoRJPNk/qt/LhaELJUKyhptujiLtYndavbld+kqe7gVFWEi7SXBsEUOKRRgS
1n788F54tgPhcmjC8NB4Hu2g4ohn0Ro3Q5KsDzjJ1WqZn8mQN0Db0uUY44MR84o+
v23lRooKQoM4WVTfKmrLboEVmCRXBG5MikR/qzPchbDKQL4LBbwAo/w7BU3Zu3p7
apDLbrkDeEdj+XBmo9J/t6044OnaV0XtnuJTu1u+BtUReL5ClTzV4yZkcgyXcLxf
eiMgUJkPkbcL+PMHCzbxxoIMg26hwDCfDm2TyHxmlbs/Y/+JF4D7qZzJqr290Rxa
Z23/EkHlfg+P2B16zh0ogaWiR9ivF25oevWuhZ5OgUDkfm7G1uHxgBUddbrPLMfo
4nlADf7alvgIsL4XkR70dU14x63AAzMrst1eP9IUNOiO4yQH4NPs40873Pz5WvA4
LUmhTDVxX3gjN52kMSosCeu21QBL8Leaf0oU2FhdlMqlUqbR4cqmFD+fkR/ftACR
XPQav1stQzMHz4DtcrHE4cXh5BycQsTkZQHWbOwRcx1Kop+h95+fyUy1GCjtuTWs
HEiA0Vg+v8LzOZxCIkvysQxqJApF1hEWJZmkzOsLuCYKh4f3o6AjUgt92gg+3hy9
44X3mACm4niN9JRG4nGRdZeEq0UIgeT82HXgoCWgEb5JjdnY+MrqP7pHDwIwYWgA
Riy0evvDkhNgT8jPgHIr/ikKYLrvBrSEHH0wwDxCLXIfTYHyYSp2lqe5ss3oVhi9
Bl+Y7RHOwhGx+1RFUbHjaYPLjIK63+6NH0Fm3bQbLa/YSFqVaXu7boInBAJXCGmv
wruOqV5keZ5nlQvOG5pKI0UvBjiWm9dLUchVrjrHiyEm5U+hURImOV0/qtI0Gv6Z
OBI8LJWV3RyaPfWK3YLzCoDpMlgmkfUcTGM3WKDEbuCr5MAQLjM693i0P0vPlRsX
B4Q3z8EDOeliraMNUqYdWyGVzZITZ8U2ERck081PbnMpIHh4xhNqLCLl3ov8K9q9
BOuamGD4193VXmsz40ZJ2K/HhtGepjNnSylfunw8mRhlfZDk8/4DNCP/DDzMArnm
NdyK0Rl/mwDIQ7486X4N2GtdKmgDxMyEOwvpTdLmOjZZJP29LbGMi60LBbjUiySW
Sxl/dCyF+u6R+H8d+jOb5Skw1c1BzYRIbCDCFQy0gxKAWaskIciJnFuIARFrxJRB
9cv6u26bRvOh0d2RLqb4OLxuGKmeb6t5Wpav4fpC6sNk4eSY9M7tShrb1oPqCHbx
2/7CbkZcgc5fKYICY1/n/Tw/ZMrTR3k7pt5ln6zeUIEaYiDKi+wXJSefJflTzCkZ
RbefxKgszEUDdYArNqtgCJeG0iDlBAixQJX0xz0Z3s3bxsGz/E+BZUSPLfDF5x+Z
bs+8PveUHxHBzcRX6g7x4eeQcxTiautUYUJT4hmOaB3Oxvw0t7cay5CO7ppK0dHx
oUK6NwoSC4ItO1zSfr0UKVDL7y6C6QLeapsoMtusRAVpktiwjO4tqXu0zd8kKna6
CNgo3mR//mpZJHoFp9jfwODREOmSKdRGoYV4elDXKzrzKpP2tEqSvuRaPO+F0JGz
z7GeU8Rdt91Atg+GuGASiBektBDNZ9ltd3aWlofWadWHell7XyZJM/LjqvD7I2Nd
tuloXXGC/rLvRn0S1kxy+YUlvoajSJVhNFBo+vgOwXeWPqOGAbokUrQV6vqi+GgQ
cqsqBuEB0z7tMzCv+2ZxYEK+FaJQUMDMIjLsGZRPjHaetDrRzoyrn0aui1O+DetL
ZDbCvLVC/XxI3aPGMNqcZurQp31OH/og21eJsUu/HC3tkl2NgoWPCbSpKjgvpjwq
/8qbFqeXBYJ2C2rA5YDZJrt+8NxihsdHHcg1HE6vtlaaICqUce3ZLNiiuUG7/OIT
MCs/NNTHUqpiy6b6HJ6TXVBUxevgex7UqDpemRpwQMgr051+VpLKOl6tuoSKESVJ
Rl0dxQCTg6eUo+cndweb7uSGn9+HWJvk8/mT7L+zb/vBytrhIs72CniNL62/KD3d
0RaMU2qHyLwuIrBkG1hvA+s9A5t0irkuzOv8TniJ5Yobc7g6Ad99bdxXzX8OoJWV
T8u/FtGuCslBX6FqqwrW3VKDkkzFxYrVQ9gHchQCyUORRJ5Ta9VHvMK/SuMHYRZ9
yRZqOcd2+Ro2n3Hc4MMXFINPnoVK+9t6BuO8UxAQP2dMtOlsp8UbMc0SR9eZx5fZ
skHdsvDsz0o5LcGmLILTTWJ3aVlvwMptdFCufMLYlvKcWgLMjP5e0kHgxFIwLaGT
iNuOb+cZvZINbjoJuHT79sucwhB2sr2QdqqQ+Jpx3ULF05JSRf8pXZFtA7+JkLkW
kxJ9eyfj+m/EIUh1cn6VrIWQtIZCUByvZgpN8sCO9JNouKe7OlO3aYKBMhfmVaZv
TsIc/CRfjwlNkTPGflDcdHn400swwV/p7viiKThf82+rpl2vHRX8NC3CyvAzFKbe
Ncb1yul6aM08i9I/MRNaGuszhydi/IkDqQLZRe4Cpo7U8Xx8ffm+piYBRinWZ137
7abg7lMd2xsJJWXnicOzlIXjePcT+A63iyt9mcTjGwid566v0Q8OTjoGZYzMa70r
pxKcm26c3VUVoY1kg3FZ+7sRG4fj2v33yTpNmE41SkGxhw+z0mG+B911rlhTycXB
q+hvLFoomkRMMPV2c+Oc0WdpLzaWkfDeafX1PWp55r65LIF8S0R9Ak42cVmzAOwK
GUPAdgRPzzaWa8QugpGThRu9eJ+YMbH/b5OjWOBWPHaTV0XNHkAuL4FEyjnovVoz
67uN0nlc060Uz8KN2keVVeWUgsnOGsS8tAdDy49hANr/rYSQ+tMT3XoKtCsER/tJ
NqAvNQbLNznCHAZ8UjU/dOetk6ZYuPZwMc9ENGQwrV/1KCS3LKDyzKnuKTf+QNTz
pJBrtclrrgyszmQExwHK4yYxUbiYZyQTJm5ULVggBf/Fvlc2weg55Mazg/VdkQqS
bQH3h/7nmiKNfDZAhd/yBG4DlOAyf0k/UNI/YuG/xYk/9EHrxXiwvcEmQHNyyzPU
n3BuW5mPM6O+HXEcaQR42Yrwly8KzQnZfPGkgtiyfC9OKHNByIKmzT/Og+/6IDHl
E4waZV+GFiUh7DrWD+1RsRVndizRY+5TXxDIX0aoPqzejpw9NXaUghc7h1u6Yu8j
vSkqEC3rFk/eE34CDTTh2fW3zEgh1rOn3c+5D33FW3n2lQTQTOJoX7hWkoKVdx0D
f2fZJ6PcBNL782nsHYex08PTxLdtAJLd509j71nLiCGKqDD8uW/v2g4yh1NGkwsE
LTmRgPcHRogVolnA80RFMkOC7xCAAQUz7G+mI6qYpgLz+eUGNMRVLLolAQ1+vb1/
IdwIO/nygzr5gCc94+3BEYlmsGJInNR1sIaAMeYyqCE0Hsi1EybR0TjGL8Cy3M3E
W5L1copcQ/UOJJsYH9k0a0wIoyCG8wUIkZiy5v03FA5orpIgsvPjRus0DIloQnC9
yQ5XltpvAcKfLfApjRMUvf6e/5f9O4kdaeaSniXMQmX53eE4LLOAvBtfQwgDRy8d
8/0dIWRz5CQcD8CKtTK3CwDaHAkuUFXoNF67GBNxJGGcZOuvp9mEeHu2j2zpDkxc
tUsjmPKU0SHdZguyopEM7SZxWs8G9izfrqBwxwlN1DExOP+TvhMji5e2Mgni0Xny
2RZrhvphYAOFXwDuvQb/vYugEdlr5bE7ln94OtMXU51DEf2VHDeele5f3/li4FyJ
dyKSuDnl5aPdDG082O6CiQ0Fow/WInME9X6DOx/IgVPN2nYNyjT6An5GKJz2YgrP
7U8AXwrmzkDf5aNHyKnj3pYv0vcCiC09UiTKf12ElY6Yj194Od46yqTrnM9L4Edp
EuDHxA4VrZP94S9rEdJKtvLx6ytf+o61LfacX61iIahp577EwXwQbRNtpl9BQy9v
rMxm8/IvmR9TvTjqoBZ1zGpVtGvF+7bXlX1xgqtNE7CbOAo/efXPjcAk5JjodLUB
nWeVVCZlBAjU/8+oEC8Rzf9APsJON8A41T/S+cqYw0DfgG1ipM9BehD9rMpbkWUk
MhREwwLOgLPCyUs2JsyVEe1Gycsj6mgXbb+nl6/VCeJ1Hq3KbwkUOysI+0xoNnKi
D2TfXttZE9uVIaWqOF0JwXzCQ1BOdjEeO8FCcSmgpbM17sHGsBTCPaSagRbXGrD2
ZGi5ZJb1uFhnpWrsdr+vK3dVR/HHltPn6Zk4b1+orDl5YbEeAlMXZC1ZZ1pQjZEb
nHwFHN++D4wadZEMP7e/8KmbFe0IVLTzSTutKkpL7Ult3GCSODs+3p9/YrpkAdMi
4YwDaws+0O8sl09Tj+zumFT4Na+MC6tlYGgUIyae9y1DcrrrFRA0jSnaO1Bdu9T1
PAXFwxx6HMh7O5BzK6/WXuH5arlaRQ3BpdbUGimQGiqh0OQAV40z1A7hjxDxmi5d
mSh/wXfL+lVm0fpxKYBSKB5m+kDX2nnZ3ZdIn//JWA++IKd37owEgXWhbaWOLYUR
EoSxL9W97m2HQnmezRQtjTMC6iqbGFMFx4RfpJRl6rPwjlJKQigOqnv6xWjyfyXn
mQlv36Apu+hO6QqxvaW2u30PgUM9AaaSH7XsIqMBcq7MYe1nxeBH4x6NMKuueBUM
WbMl2D+p9WLckAiPsLM1KkziIuLJQzmrKvxFKGSvnzYjo0XRKgsZD8Qs9+FOFEf2
5b1FRsv4NmqQqwgJ/bIXZedZEC0Ow2WV5xkA98y0DGuM2xk9zavaJU7gUClUkodL
FisrKgo1/eXMCJD7jrJJ/GswlQQS83g5qCIRSEocHRTm6CNkm6/XiSOHu/BaxzME
/wgbx3ypfxHZYiOXC5X9ogudYfl8dyVSowAtmDvvruVmLulxdT+HtAsRJ7GjryK6
XdDPXIURFp0NGygh7gfQF48931ThAygiMZkBtaCRyH0G+T72oLcHynvchsLZGHeB
bJfm7ylqUzye5Q2k9oDcK3QtuYFdN4rEPmEY6HA+aACUk01UDzNJOP2Jl6e/sLLJ
rpGIfrl3bCeHuTd5FpQXPTtIeo2Gsrqbndhe2vud0dK2lb6s5WlWDfWzEJUOZlf2
xLCekMCtqz1V4KqWI3TtZ6Zvfc3EZKKPMF2qbWdvOIQD2l51IASDPl6DQS54m/Gf
9XBg+4F2yoEh4Pbsewles5Y7Bb5qzf7j34Qd+5IOm9oq9o9szr+pkXUU4OMWWjvW
RHqGK+f4maLK3HEcLiInE7NERZUV3qxgkqzB8Krd+RXjnyg6J+wPjyassx50g9Gp
H+bwbThPPK9+CL/SaaQ1KrAKOHwTp00WpNxJ84KkSG3SAHulUEZJAIrg3Rnysash
+Z37TbKUQ5Hi9qZzWcLpd7YierPY3DoDND3WvdRl4xuD7SOKA7qIMuyFpZD0dC+g
zUxbmucY6ebj2Xq46yaRW3T7tAWcSQvm/STlCHI/dWWKBY3/YWE98gyzHgrZAaWs
f0R+A64dgWxNePcDFNUwQP+KdaYhguVsGdYxxwfqgIyVswgjUo65cH+nj7rtqaH2
zo7AZW/kISmJxU8BT5PPw/i84l51Q1LV3oPTtPfTmZwVw9EvJA0LtfC5lozca0uH
3NRsgfjnGoOLzz7dWkP+GBMqx7gD1ngH88c6VBGszJRZ4BKEjKhCYOOqBBeyCnd8
Cjn3J+YExaJbolHTKRFcS2oEq8Ss+CghbuZDNqFmsb15IEkGvbNtFcj1TSBYR9hA
ttNAz8ky1+DNJ224Kanq7zuCwojGHtRD/8+TQ6U/CvL3H9rRLfrIbnI207Y4tRE1
sfYFnOZ8BpO5WWlliNDIzyLFofqeDHhUSCfpN5DaZySEj6Jb7MrRM8Uxv99Q8u8z
EiPw/ZUm+bMQL20sIq65qkcFXkACSGOjkPvTaLqE5P7/3ZA5ilpcZw3+/AFEECmh
3AqdE6DcgvuwjW8atDHaKJqA4ibU2Y1V9s4IuWZYnGSUrSAeeGvXkUI9QxawRXG7
I3vtH6tlhsVc9CqNP1Epx0KV/E6rPoO5iE3GxQqUEnTodgJDeG8eW/0IuaYR8fOW
Psg0J6zMRvbvclGxHs2ypLFL0fHQSisMT9vkePEPQQOapxNB7XAIwGiC/OJIAxvH
0i+d2Y70sWqUj9nuglN2ZKKel6yhIlQFk5s8OkTs2stZWTQV8pFnkSPLvy+UP4l6
Mclo1Vi9Rne8mjJo8Xww6tVBWI+8DhzHN37YBqmj6+GMVnYkEMbFGfhOI0rgMyMI
Kl1Bcw+abioLOAUx29b59Cvq4rhIj9LJCogVp7UjlsvMG7dhAIMHZWd7fIhp/bnU
vjsFQf/Wj8XgacoLyRWcqJxe3TZ+fVckuSusl9VgvQK4znBKtnvXGIW28fuqb0xE
g+qCcCF22YfyoS58XVgeBrTY/x8OaMX77a7l0PjKokAwRk0F/r/RmzAbBEIZbQ7T
c87VSiKwZ0LXvAkZN44O4vWp3/P28+yADiLo2rWcrnwFJZ53uKDKOErVAL8XJpau
AYfnfpkdiv7H0eqlreauMK0d8Jkhrf9bK62hOCLxggEIna3kr0R/DOYW+83ygGN3
Bb8eaAaWiOu0HkmPqtopq+1IngSZm3qDRYtYeRME14b3Baqe2lTTpcy0M+0TYupi
7XIPMN524mbqjfRiIMu+L0SCWsZGIr+nhAsuRB82g2pl9cYZEt7/0dIqGTyye+nY
STok7rPQiiW4+X7w4vIIDIikXhG2Yn6DW30XnwDXdGgCLW7j1HLSswIQ3HJW1lai
opHlOI5Uq+ad6DUvCNzUkiSNGJj9ERa4vd58+C+0B8VBlI029KO27ZUjKTvkiAaA
pDP/ERZPADks3G+xmj/VL0EpV4ECjzdblydzWRAFCoY0xl2OEZlWFHZP6KS/1Amc
t1HrX3bp1txG9ahPYK5B616E1F2RToo3dnc0I3f5Y5PQ4mKuBpIjKOFajL1YVeZW
C6cV5u+FYuHhXLBkwbWTORPkpZTtapcteT7g5vQ0uXu3IpW0SGI8i/NkTZ807+Q5
8MUH3Qxfvxo1U7nG1WWT8b/mZEp5riQoGGmCg+hPfUZ54x9jdBi/3dr9dmHOsmqm
N/0YEQqFEBEzFUfLiXJQVrGW+hVt99Qclab0DOymvGamqq3H+AKNtAoKjXmVTpCi
OYHa8dSOo3+GSG2DnG8mGylSCt5Cptqq7i1jTU4bkVhS64ZGgrG/ncPXdPGLq11G
BA0RJT3SWK3ZBNPkUyeOdMOkPqBupXPGVARm281BQS6ndvLVDO+6KvMDEdkqOe00
bAufet87pTDw5J9G49uDCtNH8PFmY02rgGOTLbaa5NNlK99UNae/BhHpgpvYK4as
8omE+bs+0P8SYJQ14+OMfhl09x9gH1jqWqVCRGg3+rWDu9cV+tJ2SPZKXdeXXEoy
dmpjByRKo73xIxTkYevgWMxVE2L36unbdqcVkD6MTUE8E5J1DgJZWMO4eCbTYuCB
3yn0KwaouDkCsrmT3csC0RFtY3Zt5mq9YkJg9SuV8U6KBcxT4DxL3dup5qMqz9Y4
MhCxexvAvf4hJzwFDHX70xQLxqkeFI9zliSJpiWg63uBsywOMroleiMNG5+yVzzh
VnI0YZHU+SIuNrOSKVFAfBniZlm5KvgPpTeitCR/S4h/g+lHJyaN/9VvW4y4UR61
wcQTQOo3Svv7thyTrIrMoi14iZb3iWYExUX/YB+qHMH1CwUB9p7GnI0EA18iDIM2
XjrX4BPcvxYp355DG3afsQ9aAFYmfe1eGlwydI0lQV8xD1vM3paFXwXv1xlxEZuZ
dQnKA+FxHKMNomIsoLUuHBJR6PjYxmZNsAURjABPvnkXuqE+z7YoTbm4kMqwji6I
OgehaF+gdfr69hDaWnuFi3jRIVdppmlhIoIeN9TtRryy7LYTYuJLqRCJlgv+jp3z
BPATEWkZ0XEleWmlS6Q7jzN+Get/GxRbP0tCBtNkDxllDv2Kfea8xMvAi9UJl0ZA
DWvet2Y3AMijQCvSYqQndOTpkS8SFQBionvSL20xLl6YqXWV7KgfmQY5hzSn1Wy4
7bB8nj5tk7aE3QLERWeq4p8rlnWFaC2tMLeJ+n/r2hN/byjwmswPDB7G2x4/hVyi
8+KcgrHXyx7WNIxNK1iK4D3dKZly319EhVASXVp5v2/ka1ECnlhkqlga10MOg1sw
zpEf4Jzz6gl/rNLyCOY9lz6YvbeEb5ojVhfyKQQCp1wA/d/WnEY9QBy3cCHFKiWz
NUqSE5hvujaduCOyYGeuiiyuZn/GGUM8MraKVvgMeV271u2V2mVDVo6seSiFQk45
Q6xpEluhIjBj5nY76aGykgvhYW0qqAuHEw6aoVGz85bfLntHzClFfEfmnhQFoRA/
fqRApZDLP/2VywWelIE9X9KdoKHu8ai8vCAuJBKk06QgBBAMk56AmhAUOdWabqN5
piEV2pR5nUcMUEnR+Yu3K2nKgBCuH8L0VhCMXagoLHHWJymmz8Sd3VCw+UbxV3st
PvmdZeT40meGrKbUPqiVjRIo8taOsMoXHwFHRZGqTIPov2qZs8OoutcxgCz1TyAG
YsBqZ+Ng0uigG2Dyhl/JwXLJde0R5992lW/cojgqpAf742flEQV1W9m6PUZ/QUyu
wJfadpp7ZY/FjV7pntGg97CjiFDAlKi5KfpCC233/jp9sffJk5B1nHnKwgzr7hPN
cuq6pKCdrjSAc59S8le4VsNnqxROh8hJH4qOt79Nx9sILSFSupRP9zgRxgPHyFk0
hbO3xFWiXSy02RP9ZdV2USVOtuOiD7uCtHYwGyzjbIcJvxtFTl8y5WCfZcY+saNW
Vj1lwkLK89HApuc/3NLZpFaUYQXGotkT07OoVgdZjkgZEHFjdk9tJxeY++uFEWus
XXTtsCRQ09MHIrvxBc11XcboL8yjEFemD9HF/aq53E4zWbJ0CNf6h6Ut9MeZ2UF2
2F1WKzfZA+rlKkN1nuzF2cSQug+3WyV+7q3n3QKCtwbddsJ1vq+Mgi0jlacjiLOE
wk3nEBb1YhP/tJKbdZyA915lc555lkRYppYxwb8BJc6eD0MZJWWeJt6Cm5TvNWZA
xzS/GVq22+bxN1TLaT3OTYc+68MjAFc/0sIO1NjF0M6fjJQ6Jvhe+6CGM2JFs6Wo
KuIFYC53dR3Cpa2Qv+blZYlBq3I753alUzrdWzb0M8CeH3IU1h33lT+lTmC4WTLR
LxNAlQ5Kktg/+4s+nFqqdZ41eO1JCGTfhplnAHoSXC/0AxXPJwfu/msnJwQeW09R
z+/bnksGFsAIqmzULs1rLweOxarwaLC9+bipK5ntXhF8MKKlaPHYWcQgwnSbHVBe
zF+lekKN4ncV89dafP9oRINNurGOigY6Er5HXkD+v7d14gxItw/Ug0e+/D79cSp2
yOZLiORRfPy8R2txULkKjF+TNRlbcyfCe++vsB+nd2Hie0XIJnB/ht/a9VooZxzO
K3H6eqlK43sYcBMw8zKdCkAu4PskMvZiRVFX31iv/k57vR1VZmh3baxEcDneTWGg
N4sNQqHB2TtB4YS4wwMpvF7f0Cf5razvHIW7tlA+uocWAsO+a2Vt5tmuB2DJhgTN
dfIlNcUnCzbs6PKij2O1Ddy0uvBlnmjak4sSmeUiiBkTRlZKf5Ta57ZnRIO0lUBO
L7RbfutxLiIVw7shhFx+nb5wqiUFOhminPX1oEvKtkeh0DURppHFdJGio8FiGbVU
CorZvIoqNDpCvtiZWAzcZHGq/90zqW5EUlx715yUA9j+OmvOBq5irM1CQIpbMJCm
6LAcBzj1sqDXFxiLfImW7CZ9U/cE94FDDzCIFMWeh7eE5ZT6hmzYVER5VxNjdLMO
rDnrpA00Cjc9WMELpyK7Gz7u8x1L9HJLd+8Ak4d7JJTw+KmYwnaG9FB8TcWS7Kji
lglk2JYYViX/zk+hTzlvWMjrGiIbPokFzBl8uSed1vNhsFlxXTHExhMX4kF5vSju
AJ1U28BIeQQm0++JB+KvrsDdp54NseBzXuAUsgBYA83i6cf+EfkCa1eFvdb4nFIm
aL+RO4VCLC0AqevdoubKRAQEvaiVLZgOYhs9TEo6rTen/YAPjBEE+Ac8sCLRtE59
DrnSo0ByZ1FHzr+nl0erHJQJnMDrNUaYOeQFZ5AkrWrItzQoC9UkbEJOgJe6cHHA
SGvQCLB9ItZGfmcdS47Oc+yOPlPDmuOiYF5dpU44ijmw8d7bdKNdzN0HQK0hbM56
iXNb5zVM9YFhzZ9ozuUWwKh6ZENbfFDdUAuUg3Lt72Jpm8AMApgzQsgdwVI2frZu
eKvUiJuZlvoYCAPPOWDEizMcWK1tZDHnJPbx8VtegxT2jYVGmektwMidK/M8B+pm
NmWnVNA5kfkr5lDbE1t8xz2kvJ/cou+UMOQyCr8w9lOnDRnHApfOcv3gmuhRHtyh
5XG+48nL+0CJnIiq2abR6s5ZK6kGkTrYAuhNnLLKuayy3EaUMMX4NyKwG/JUFsWb
oVRQ0qKb3rBdalmM+sNhojDdmd8JginKAhYjWozaXPWA02ruGHb/GOpBrUz63cDz
5lLCCC8uWGw0WJ8+hpFD3rtDUf7Mak7sZnVm2XkRrQMiJACP5JLyzTqTs5ui8cg/
O2Iw0uVH6dCmlrRXWps7UO/TCcwVXXVO1EJpodaigDtPln7yzztb4xNxumjJCjPt
0H6RUjC3x1KGckycUAMA5VZmRW/NzMY5TZnm6IYMiypuTUrLu2EkIQSbP3tetzza
7Yek8cxDavAJpnIFXBQPTCNkhBK9Ibcfa8Sk0VQ7zN3GgPCl6Gy5gHV1XJ9KPN4U
K0yejHzTdG6ES8BROcdyQShwxG9pC4mkM1Ig2jai6+kwY3NpbPxBPY5kfYJfEY1i
3bV+AUsbDjIdh0TdU/rI8MDE1ECdh+n2U6+el8almX3cbIqcUyIEGQHJrkqdbQWe
2eS9PnSgVi58USewF1rZex2TmAr1yBM/MoO12WMgKGFweeisFZvDX5TmjuUwKaeD
WsvPXQj4bBnKltVn1j4wnWsx6caFUOThR3aiO0dQsMz+ZuLwma4/0bgA5uy6BRgL
+g1uJmpxHpKiDm/FrdR21vnmrMaGYSg+7FkKnlnfc/TLj2eLhx90weAUPB4QO5xl
d2ZqDD46ZfJ+y1In7vrfA5ObdvP9fDR0CcplVf3pqZgrx3hzg5hkux7sM8Ol/via
swHejd2XNXj/xxhis48lQsxdTiouXzyQ/HdOClqRfvGcD9On0RscPmNFhiLUIpUi
BED6XlPhvz8iBngRDtRte5zO2Vz8eGFUQDvCzNw0OwAs9vxSKu7vUUMYS7KxTGzb
JmKsovI59axgOlPqjLfmPYoiXL9wHyAbAVuWTHv7sDQNM7Di33d3JDpDczLVcN53
YdoOOjaY7QsgXt/GAH14+m76UYczMVTw+v887aJ1RuhDrgLVnloQsNhQ4SSPpSbq
MNjjru3c5pZBZKrEBBr7Fr49HkrN45xr4saAq06lJP5kGE2UJkG2pYS7hH2RT6A/
fDDshc326W/Pq5y7xjDNhlcaRmqlkp1ToTGD5QnPf5A0+giXZ2aKWaW82HJ35Jl+
Dl9brohx993yq3YacSbNmRZhNzkheTsfAGuDWckTHtWldzyts9+mTima12/xLvch
eaW4DkFwX6hXSARKHiIaFhZtOxZ92ke5rLw6HHcIrQxbuTZEqkSIBq92NCrd+P0Y
SS9Mh5JoRlxdXqdgJifTJMc6G2Uu0htM4DizUVOA9Mhis1gRDVq7/E0LscVBigsb
3IMIcCi8sCHFqpP0F77/b9ZpXILWJsJPwstnv+N29AJvL7dG8S2CTSVnDONsgAEl
Y+KTJiDh2LyL0K6ytf21YeQCncACIZa9vKgy0C9+ZU9z0a+s1mW1QQcg6nQtEoX4
+MJxJUEJdUZySPh8yXnniFgZlr9Zh4oJUa6nIguBgXzN/uzJWaCuqGHftU3JVP3O
NVNK52qnwD1iIjCyc40nGtNrUxJnoDdCBHyuh9uB+0sMACWQXzdB0Xrd31iHz26V
P4uqULk4aD/m8i0iXwuofH/A/p5g7CL8UL/u2iKY6w2qTK5PF2MQ1clQDU0NR1Sy
OjI6WSh8tKeIR8wgqzl63sxINz4fVt8tl9rR8JqqJ9/x+6JUDUhteYwJy34eEoZj
uRBPq84vo5pwJAUdaNkIOSzhqeKN6z/LFkJBfS9ee7jWVA9kWvbQOPWfVSbfOwJ4
ozPGrG+pPwsKB4/49Bpgisc6wdPm5q8FmyOHuCqILuAR6MqJWW9y02AqAE7SQkWb
4e8aYbJvyiNQpQyw8xMnDTg6elTmUWEcgiOYcTxAVY+fYcwqypCe5fPqDO/SLe6V
0cGpeSHJvlN8oJM/Ugyd+VkomLGfVirNDoOm7uwz0oJvEEp/vz1SWb+u43WRAsMX
g4zluSxNyOSqcWTWd03GKjxO2hRdWCZO1yQCSi0QglznlfptNEGTR/48dDFOCeAH
yY4eH7OyfVRqceROb3sHT0crIxo/siVlili+i1g1qVZqLx7kkXQHEcbBrLmpiPqd
feKaNLAw/lTga/Cao5ghop/EhwzcttYZyHhypA3yVpK2vc/1KLbfuAARnQpeySTP
KoKEObT1wk+wVbHNjhPBiLJWqXLgp8AZCB297JrkdIJscsFVfu78LdSQ9Xf2fatu
B2aARDzDzT1pmFQM8r7GKnTlYaAnOIlRgb3r6kLuOXzt4Lwh/4f7YW9FmmwjmtSW
jzQAgGI0nwGjHDZkrTx3tEnkY1fUNYpVj/tQ4Kfm5iX8+hwlziItXI7J+lGiEhTG
b4umw/jaCJAFSoLF4FiiOIn9Tj1of3xK2P6LooZvgTLkMtMQLau1GF3vJpiZ+81p
duWRgoA7NMeYZeyZyMkyR7teNBU1uqYXaPdAVlqp8UeDedLPXWsV7L/czAMwYC2B
VwGGPyb6mD8W4e45Ii9n1CNrNrp2SkvrSL6FBW0YjXQR3ObDlB9FPS9TpR9eiJr8
wvA0CBinTSnsW1hxpQKzuSdvMMAy40o01zT5ohZ94ncWMlWoK4qkcdlI62HY+6G5
Zk8cqS4sK7NP5/IztOTzfhAq+DSF+W0H4TZ7qmDd9cQmNaVyN1g+Nibl4WBlq9wO
/zl/5n20rX+CIG82+Ylqz4CpUKf8ZfaiOdL1iklfOEfpP5oC8sruXJnI5KKA4CZI
wzxVL7hMOIJQ6ZAHvN/9B1W8GsVxmS3xrTMj5SqpBSeGHJvrWR6OuMO7NUNwgKCB
/gKNYxYMpuDHjLgFAzSsQE1JGRJAgWvyuDG1mmyOJL4QC0H4jk8vJAdZ+2GpBdNO
cE87WeAohcntxpV6SxSP69qPoaiDZHVQnPYYwq3U1m9EOZBfu0aU4gcpQJoUc3Xa
Dti9CR+LeQ73LrAE1a8HsktXcwpHv1i1Cy9DypGuO4zR8zaMpWpH3wtS/AMXxegf
QpeRsVRgGLrQ8aYnOApqRJfgyGIcJSHb9wCfzI9IbUoxdn9AFyQdMLhQa1SBgCHe
SAW438mVezjyNIN+jAFXOFHt9TMiwDIOwaaTkVuZAC9Hswyy03Vicwu6m0WrkUTl
R43G17dSF/FlX17nOubwyLVoisdkl2dFsHnqBIzRHfG+Jie4JoUWPlDtlzNdD2mA
UKAWhJPILZDdWEwq5fr307tHOV22Xh8Kd008vSJ2WVvtGBwW3aWveZW6JyroySa1
bJIprBX08KLQX+42GtfN3/O8Bvu1AUAF8kSSCa5tdUSWF3LCUmg/2T7nZLUMaHOi
GPGYHrXaf0aQBMeM91MFv2PEWqPmLmKfs3lKNR2IyTiIOmsCBy7aQ2rxBIqjD0UV
B+azzt03VPDcHjXqN4PLbnyTKqXhDFahIRzkE3TL8Va1fdFlfTiyYZkdgHLYgFAO
zwHfIpiCYKPte0vGd/qXni+8bW2AZyK+8PDGDYdPB/xJzJGvP3O1qes6HcTI7uXD
v2QOoyx6Asl96E9S2dr1rJlDz9MBaJe7gPJ0IZeC/UxCsz2p+IIWaWFol2/t+fyg
OBD8atUypPUl+uoFXzk4/Zg71oK65Yum4+SR9a2BsCHqUp/qCG6GuduZ4bD/Jsbh
BAqa+eNV9ZCTo0G20gft7dOwIcOSZYBMM3FsjganH6uuFpmFR0/LPw3hcGa16FlF
m8EEDzVlyDuzoaP57xQG8A/sLC84Pd6HKn26dytEldzt/A074v28anlfX2EqdPvZ
6RD46Ag80DCxeWk6k1TThkCW8e92flnKpNqkkuOw9picGrIhK7LeZEryhI41t27u
Hl6BXtfyqg0F0KQoa8HJMx5joaduHLtyDmEthqIodVB6lKuqFiHBoHKtaRyLn+VH
cg1DFRufy06cVeHltJvMbZcAWi5cfEl3apWy6w0leshVHZ3+RcQUUbczeCdriDRv
+v3/aX3lWh/XlHZw2GWhgEPqNvIGDWWGbZJW79OK1i+QXeUQVCPT510XljZ+aktb
ikXRNrvkchpQX8EqMkWwJPOuWVHbYFzF3yyBNGTkgXFJv7/rPFY/mtBdc7ekVEz7
OTrTlRotakNmPl/NGZZfpOX7zvYcv8k0Sgba522To+sgjbnTBx0kGYbZXnRsta2d
bR7SuDbzF2PRiARcLuvuB19YWVUs2KQuCAD8ic3C4O7ZA/wb1wxYKzsEC7gkzex0
9QDeoAdSSvjG9aUY1gawWfmT1VGDkt0jyd8OJPlVYy4axmNPCIGuqoPZ5hBxAWbe
rVaRejcNklvjrPYt5Vh18kSzE1TRTbTcvS4pmnyeHfw/kccIMuk9iuXDMfIi74Ke
NFM1hxNR8gms3stJFk//EXdmmFc0U25IXDHQk0JrsQz/9G2TOo35ALQZcpRwMzv6
JIFoQRCTIRL8Q6G+w6meeOKe8NS5RCiZpUPOp8KdUQDhS5PbDduxuCBH5Q0apAYs
Y5QhovLf+Kp61Qun75UKwBDKR48lM3TBbFq8LPU7lwHA3pOq3bhbIFpQlKlK0sFN
fUzyVPWsLDbQKA+Xq762+h9ijIBd/XCdcMmwZJeuGx0IbdV+ez3uyc/CFu3Eodsk
SN4HmkA7PGlxohpZZNLODYchC7VmnxaJEfu6SpPCPneaqjIveRQzQ0RSaGjKYpBm
tQFxBRCKgc8Kw+e1jbJVuvPCHGTB3EpoomD8UMbwEUgZOqAofVv++IbuQFaFIzr3
wEe2H2W1rzX1CS6f+7/zLseGc1ve0fVlhLDMIh6IBYCZhCZUZ26JFy8zelGca8tk
64OUoiBaPPnUqIRLM+Xl6nJAa/5OAKMmU8s+ZAorOnxRo7FbCyePV6tzMwsVJL7+
BphkLBGA6llLU3gRxooAxb9uWMYEvC7sZCAiPYY2v9gD/F6fuPIWAYUHdCQer+X6
+nbRRbPbOldUunJGl4gyir8TFyztXutmV0GIE9cit/pnRAqoYmhqTyD3nPGovRWK
QwUu1tfHVbKVHpnoeFLn9vOJ8Ises8hS2J3ozullfBBFNCmnYsMSWbSZuPVkBjfl
oa4TMMzZKzJb9E/2Cm9dXanwgvXt8YGqDocAOkX6JLqAQ82pmvEsiAQm3SUU3vlt
7BlBrkxWJWbtb9jqf+E0FA3E77NMv7aUiUk5Xem25oST6H7qNAhMqTu6xu+PiDJ+
4mlnbVC43Orz68JU9QpFzV8Zn42lWdF/2N0Asye/AmS+Jq1LuJLn2KUSiK/ZhC+d
fBwHhH5bZ9IklUfvCSQkqeQsosAwjZwNj9hqjrblb5m6eKx3Xs2qnT62nqNicVQt
jyjXn7Rx+AfFkbZrngGfrRpXI/AnawfdsDdl/FryjhOM9l6gBUS8Nct7iUsC0+wu
Wxl9naiEEYMDSXVXghtLoa98ttcMHfeBZqwxO1Fxb+g7Aq0j2CMAKrhwkgEvxmxC
UQPg6606lWUBlCCH6h7SbMxTdKBE95zabO1LaacGKt+Mmz64V48dRxpbkMrTprFh
on154BcQfcLNEUsMGrnAO/E3z7gb2SjT4d2sd3NqWFJC0h+oFz/1jd2S62AMfX02
ktofyjVygyhBB6/Wi1kuyed0Yx9ey6JHqWVTmYA+q0vlKpIzWWLjrtTDiGoj3apT
pkl4NJD0bSDlUyCcPZWxHEMq26gIPqEZIzLQsK0By3+nSQXHf65pANnKW319e7XM
XvywGFjJqiL36teuXgOxvHXuaxL8RWypECpsqPKUvYGpNOwAsQlDW1LXKAx5jNy0
8E3RTOoGyIP5g/PJvKIp/8bsWoEMxa33sUQc/3zyShi9qOamJaB8xNGcxNPN7z56
tEukmqtTV7JWMY7pDSrqLfBvbsab7awSJp+5HXcoxYmMaICzHarBJsmKl4zJ+ZAN
w1X62JGn+uJgf5poLXEq7nzF58ocaICtk6kg/S9a/7RpehYB0sgdEdkrQ5O/aD/n
oMgvwo5G+pqCvtCWzQFZwpsrNwam0w2lOE645GbrNaV/09MJ9XvIc9vSt1TT6y7s
8J7XRiHsmoJBTL+5W3CvY/0X1Y6qPfJQgiKnX3hvm14FggJcBqo2F1xzD8r93qMF
1swkh79AcjB2qMJiduGSJqEUrwnLTSHcrC4bRxRFBfIjXjcQj7BRpgLV+AX3X2l0
KEzBQh0gemzVTPKV/meHYrMtBC55L00dhVw418ytWtPQLIUTAGZhNNDeGESFXsFr
thK2B+x8YT8ZF4vPqZixl8Ymh8ucBhrEZ9UsIrGQuQrxtPjSSRLyWy5UXfrKxVl6
R6x3eAmFFWAy5eNL8kyk4ZXiW6ixJvQWq0grAwqyE/QodsyV321ULBXSLza14Ge9
T5h0UP0mzsmiFwNE43fvQvW2c4LtMaZBKAsftNMirKXgcmyAF8Z2nVLh5yvnyZlV
yvCQe1jobIXCK1k1Woanl/VMAaLQ+wDDWmIVsKSRn5zB6FKQrivzwjEG/QHb0WDl
3hTqZ3EFV6qItw+rAyZBuJ+9e9Jb81Bue6FVbiSG/Ik+4BeiuQ6zjtK484qG/rWZ
nD4X7aqa2YAVF9dct0N1yrdY4i1gqwhTBs6NAaIQt+4hxa/GgcYgp1LTSly8KRhW
utwL4bJ0cb8CPaMXxTe3T+fxFW/HmrLnRYmA8f4z7s6PK7lGx5Kssnv+0rDM4vsn
FUb33IqeoGlKjYct8LiU/MzyOAHl2hIyzgsa6tq2ZPWhLGXz1fa9KwMBMDMDY9LO
5/UXFuNjNLYkS2ZaMIkbjU4kYOI5qMYPEpjiKslMvhjq0kI8OWQJRejyrb8bLNSY
NrxIM/7M4yrxV74ugGH4oMx22q3EZL87Q4h2Hbz29l78BtalzsFu98moRDZ7+hHW
raHUzGs9lJ8JGzuTzNMOk4Jmw+3dPjs39xB2lrWL8yPXovuXTGkyoZK0uqkHsx4z
LPYuxyaNQ3CYEXBJA16otrr86+Eil3jHa18uXIfGKHyHoLas8RCSUh/a50X+N0oY
24nKZjxTje0TQQSxJO6qA1BpG3zXCG8nUPaX3OYFVRBvrT1fJRP4/rR4ik1LlWKx
W7L+0fyzu1g2ggg1BisYIvFZmxd5sOvO6KSBYFqvqP0bc+BtZkHIpLvooZAJV+Qg
Bj/RVF8CRvnbiKLA9K3L/4JQIUYGbjGrLW2rj8+OIdpVSzWztbAyFf7ZUhb/1/tg
oJdtNX6fjar0RJfCpNH1DS4U2pHXGiFh17upKz7wdNvmopMLbshIUjv0FU+LEbh2
+/HqZ8SO275RBPjIzEzC9CFRmMPfRId0rwZ7BoY9d4yAf870el8Nu2lrAjrdKU2f
E+k5RU2lTWeOhvMilI1AOUKbErUGu30tLFbP3ZmSH0RYiyiwrtJEvbGzMutz8l1u
+smjkg9qaUHqFYPU2n9Rl4SBspE7Hvuyit4C8ePymSG8sx1zIkm3ejI0+NI5R5D0
Ii5rGlmX0Ryg4PgAE14siGvgUbMAGlmMc6P6DEdrFHFZqcEbnAfu98LeXpOsFxCd
TTOWxD5i3qp6wibg8LlkP5waij9fPVOVd3uSu5Ux0zQ4YCj9H0/Y6t8SgeI17uwz
VLbOTNEi8Dfzv6atYQqnkXpBE90DK5TFSakI9YRG8l1xnA9+8TH4ezcTF1Y4awG1
lEaJulR362285WAWfJL4FEUArtiisOuzZNSxOR/P+CV1hlGy06QDqeHAs5kLL2PX
poGv6kVZ871L22HdvlVIlJMEMYCZsZE8hrIYzLbj/CYCuX9B+NBONZsdui6NMXcY
MdK+TovwscWDTSZb+xoma2kCrx5drBCqS+4DrlkuHBqcb5WM9PcBoTeNS2bNlaIE
5AuYPp0MVnZsR+94looUtGFIf05+LgfpKc+LTIVprGbnmBhIIndz2wySGY1PmOkj
GMICEc6VKN3hMe6BJlXCOp75zGegpFgNX0u6CcOmeHw56yoQH4wV8JOGM+PWSWi1
ZLnK70yfmnmPZKj2/rVGf281kSW23380OaB1pC/ABBrgK9x7kQ1K681qmL1OEaJq
CGgyaO7QAeoml5uXmRNLokda/e8XGmskyrXsP99ANYtLyoaVNDK8pFjoRycf4OMT
SdDfYmUCaWHeUZbQE8NhCZynof1QgSbEW7LnfmA+oXV3b0BV8GZfFC0kluS4UGJv
wCIvbIpEFpbMK465UCmsr/K0yLW7AjGzjKOa6DwRVGql+vY/7bTOV4AJG8vfG4oB
W2qlw1CT/lhCi4zu99zkEVbw9mScNZ8v68jNg9xaN/zZMDe3xgI8Y7EMlnSiu6dj
s/7JsaYB3NUA+fU2uuLWeF0Rr3yYpoS1JJcuGsdXPXKMrDsALC9Zk9oFiRNk+0/9
rs28IgWsd0SMCrVn88eSsR7kWxpnasQnDSBZhkgrMpCGqsmZ1VEu4cyo18PcWcSt
y+guyPJCIS0N7WxOqXkoLDqHKmWefgNq6MIzaNSDyYrBtNbj5zDLGdfLg2+2TPqX
MEA0GLAJ7uHon8V5rT4v/TD/AruIeihr4XRtZ/0yemckodcOkbxRYnyky2fM/0Mc
YjajSkK4pij/4ww91t910jBTL7srYvMAaFnG+KvH/QvJuG0Z4RvvBijosGhwmBrA
WBtVEYT7fcz36bsYh9Nwt2WGSZkSfcsrqOgqxRODGU1i9i90EaoN/kRINbq1Xcvg
hRrBngxKAKj9Wgo8iDLkWJbRhtq5VvjfZcDYs9YtW8eEWTOoni4luX99CFx/RVC7
fgS9WbMXRt1rtgXA5PwXZb2umRVyeygmvXYWurwYtMORNsHmUKnJLYuO0/t1mh8c
toqsCdVh44Vov0Bokq7z6Vwiv7c4QJ0dRAexyevoHtE3qzw9baBoXaWApbGPaTpZ
uYr/4sSoX8ijnZqcjhLbZcDCgfGi69Lm4APiR3fY8m9GfL0g76UDhzoTi6T36xD9
RCFTWTJexinV4ucO7CJkv10SIi6pjKGI2i16DgRkoANLPBzx8xag+8g3Bs2O96Y0
7ZnwpzC/R6jn+ZA2w8gd4lAclEeIrX/s84yiprCYgaZVKhGEuJmh3tis9oMWU0Re
aLWWV3l8286RgMWitPUXUYeDFQC0OIrpiII8SmmrFFOIj5cQur0jiF5vwpEBDAyd
nfDjRhb6BRhOHZ5jrKWS8NICoOuo1j2i7KaBdLkL2aisxe6ljZGURu3/xFeR1UpZ
iPpKBR5mtB4JnUXlbUx7/lagLExSVB9sMwcbuOFvQiafIH2t6elQuZmj1P9vAdQe
7wlvWgWcUyQ7/wXw4ZL1pAYBGD8t3VRQIzvOCZAHElRYPGleEDQW4axe7qbeEFIB
L47xtfhSAmGzvcoSE5grKCquTWB+UJl84lr8oFGQ71kd1i3c4KB03KFaxFuk15pl
EB6FOZ4a77u8/GiG71oxO3a2VnZir4dGQEEuGbTYSL98d+pCRiTPDcMnUL9zr53b
teCJov1tJTFxGd8aBeoDE5cDTSD6NoIr5bhDf48kXlCYjnb789c1He31/YmkKRra
E1USqgjSLULUSTyuynoMuh+2Xbw74sI/bzvUW7K064Kdp1uphpH7SORS+NgyeBUK
JtUpEvo8XLBkrYrrA81yfRTLpIlx2fql7DLcdVev9CZdf02ApDkNnkxn+RBPx9TX
p4yGBjYD5sHw6Ln8qZK4fUxvk3OHg81GI72u9ktYFjuaOzib+rJhU3W8oR/ByTQf
5f44LJWf87yitlgXQhtzquNtb4L0u7EZST+OpvIlkmlxEeeqTmVgjhlARlkr1Qj+
eGYvlXr00dHHhvIV3Z16E7U79dQpTnzzAPjtCmUCZtoZ1qpXvXTvuZoCjUWQ6xTj
9sMGMpwRqgDWbDggRTrsNDmg1nTfj9qUAGIYEgaUu+R9pwa39Rnj0c/k4/HdVCUv
8t/j34pkxKV++D8PXT3PHTKix1LK8V7TUraobYILGirTqUCvxd6VIMyq/9a7iem6
vxbrNeC07g+JOs9Q2cdwkjOtWS1TNhBoDll53FOiMddaElTR/sjHY80d9hUhwAv/
JbbuNtW6+dlH1+a1Xqkb0OlKYFYeNbsTa2CV5bLrcUvX+SPledhsLph/DhSn+PlG
obFHoTrm9gxBWziEGdiSLUl7UzYWUF2VAE69JiXHD6GrhvCoqBJaiR7hCEyn9HtS
zM07hQ9DsBbnYF6SBC8yQlFnQUMKSNYY/tXB+RWJ2CkbsdqJX1YXBmfzN81KPFvY
+OL5wMxbcWu55qa7M1t0IGpQNforX3K7PrK8SE5EAH38EJZJv1ZdCOiKT0t+VgB9
AX4Q9Abp5UGUJOaqxtrkqSCEaBF8O2Aju4NDkqcWlUqV8MhToqkxGFJZB9QWPGWd
Xh9slUItNxTE31ZkIIwOKW25rrwnSaELOGU2si3tx4HbWvD67nxXWZuRe93OYeA8
8TtL89mQAmVSFGJPe/MTy2YibXQ2hLo8V0Uk5/PxJa8XHKEaUtO/4Gl8Yl4GNugz
zf4A/KQgJTWHtRDnP6A9ow==
`pragma protect end_protected

// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
cDnvk+kXublSoVaorAFjiSt3cFsfcIIfKDpUBAt3cSTbUbixTaQYfneD8lpJ4cUFVkxk/x5ybyMc
bC0jqr/opnkF9j3/1+qNbL333tCrY0rId+BaLs0wSXKoT3ykyn7Hw3d/1VYhmXsaI1p2X2ZC7hYX
Wx1gQ/fnIJgNVm2DPSZBAc+bnfnLTueV5DDsI2xVstFf3v7cbnsoySAEniiZZ8/lXP/AjS+peU/b
HeBZqYoS72DeICK5BXJ4cJlpJPIsu9lur/dmve0oDQzAt8YWGTIU2tc6DCiKRt1e5x80gCHImDzT
Y5/As3wsKAS7UsQX5QlScHg+JrRhgF2G5j0vQA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6xlPC09QQhsbPshyFn+eEJl/brs4Y/Zz1njBwjaaOtetEnwlT3h5zR3+y1YwIt5J9Ad6g2HxX+w4
hBeLlbrmfToyxX63DeGriWHDUQBsHW48BIzvIkdKOSz1MRYPnWFD6tlfDjRX160GGLS7YVVro0sb
TlYwme1cQZQBNPP84F2hDNt1UPwHH6YASBQOMbqAL9Thp8CXUStupYcXtECUvd0Ac2PzwLrtN8Cf
4LTn77oqHZrDgmtL14jdg8G5Tn4ohzElhrwNSiiE9Ct3LoDTU0GikSLipLqrA9/yjXCrz7fT2xpt
cRY9rXBnPtRZj1thvLyZR3KHjx2uLqP7LrNUbS3oXheiu8/fCi7kqciv2r9wJ03kYrwh/MDYULFc
jz6M8uOEiQXdwi+bgeb2qFkuM+7plVvqtaq1vgnYpaH+YOSSWMuRskg6fAYD3oKDvIuzQ9B3TDRX
UW3vXye5zS/YNnlQ1QDWK6DzyUHr8wb40AcNkbgmmY4D/xoSGYmJCouT3Z5/j4Gq6E6HMa3LJmsv
NUfcmPw4Quxx/aOjyBKT7D7xghbO0M2zcVw2ATDDxDl+7lGHw2/aFcbJkZrvk8qZzcYeeBHnopb9
dYf5yj14tvVqKoac8cLmRsEamWvZhu3kboFtPv+K2aoHKTZPCNNf09MRpyezWh0npIqJ+94V/F7L
KK7X/gi3OkdfK7QMsjo/CC99f4QCvLVHvjbfEEHMZauBlFECAhuwaNyHrr5XaFgfaqOe2nsHh94k
NrVTBmx+JWfN+3MjFyhlRfgv64qRGPdsDi9xbq29WY3c6HlGVoZcgike7HcEeyPVqHGfjOS78D30
13OGWTyANtI4AwTqqz3johKhUSzoRrVYo6aiIBs2JaZkJw6aLtTKZSkuJblrlRi8Vo2vrZhX0Wdf
FTBVQ1yoMdViXCCxs7Pa+VpXVdbm2+IocVJ8FjvEY/EwphCQAPbXTfbFzA+ByO7qES8M/Ifyt1bw
zvShRn9ednWnrsMJj0/9qEkVD/4OXngrffatquXSbgWKjoHXaEhjcjCFv40SnWtYZzJOSFtvG1LT
vBrFvlosW7roiKaDvutTmdih6i9m424yXHveYvJsIghuiN53o7Vgo2xhw6AuUuUMaQ/j3IGOzwU8
elnE6tWGddE9wKEtspIDWq/tTJdrVbj5a0jLjj7TjmN4dphCj51X9RcHJ8qi4Y2KICbhMv8bHjAv
7f6l7pHBrFyhPt5qbDRzxNkTU5TXyDheZcFuxUHur2fS2DNnJg2x0M23eFfQvv68rADPK5yirRHe
WvMTTBD3DIwYZzK+nX1pWRzcK5c0xQsP+/cwYou6KJNSNG1fZKRWq+3qUmpmuWJ9Pwp+2er0jypA
37QzW/jzQitcFWFLNjmSJhYkGgdHv5R6H3H1+qpCoDtyj+Xo/UoF2VTsWUvIRgGwi/I3g7m2Kjoe
XA5wUUP0mabsy6G0RliRMQyIx4uGdrpdctWDKnA1UaUSmp19cpp55IwsZfMZ8l84Rc1LLvOxOgnD
ZeQ1NNWKzUMujkj6T+Lt8xQX0Z/xWmb2JTOnLjBXJc6mH0Yt0xyAnQe2Cby2e8l27uEFVkDR9s2C
XMH/asvIlS9j1vvR751ZjtcxFDqq72uUsoCPT+ORWoppaM3QHBvWSH/8hF6+m04XwrYdnZDDKacc
xC+7o3Njqx8qv5NhnqgtbYtOQZD2FDHFaG/vIqKnEY0r0VlYGBbvrpzLi6EzfzJaR/OM7mfuSVbw
d4e26Cb1oMpO1cuot5OQZj5iXaalirezfxMgGMvdUrMjA4DVpHn8yg3+94XKDQfgORity+dPf/a2
NKs495qEVEIj4SpfpQnqYf7yQYm7kJvx5hdhKLdLgrdcBP21yGxzMvRy3uAmjiLLfvyjfIdPo10J
1DZLIvzD2xC9SWdXarI7XI6RsPTobm4aO1+yU5tQ6xmB5cfSjsUpEWIIjp3MpyyhMhwP7Hsseyye
U6XZ23JboNUF4xRX96FDMhTrTmWnGCt6exfNXa+hXrhFBD52ziHDZEDJTHQ8lWSE+F86sBdc3PVb
RyUMxu46ubP18TN9uP8AIhd7HFfCM4+MIrbU36/lzALLoU64EI2QMCP4weh05cI3pASs/yuDQQnJ
b4zln7NmMQIDVslOf2ZPol/n/+h0+lWGt2UNxLFTZ57Oz+S+W69Q+2plPt6i+O3i/Xv4h7OY5Tes
LBYRPvWB+LgyE3Av2eXsHEDZ0Z8B69xXB30wTqwwnn8mYIs3VTaA+qQsm1f2butgFekDYVYmb474
MSAHREnf1+KMw+JLKBXhSA71335Olu6glI0DH1RT5jF5OzunT3zsJlqZ5xbgXCG7VzQiGI7c/ZQA
23DdeOkuamKETjw+Vk16IgmhqLvDPJRkv/z1smMHLGSDOKoOzIx/ZzYEXmlESSqxiHjPcqfMNP0H
n4YM+CCBf0UZFIJTnG4ht47P+SuaLUWOS96RVSDlDW3eoHFq/3k3t+dfuicplMC6qGJt5wnm6uaO
yiT4gA/GBHjiW+u9gUqCOVcLSdU2cOML69U+K/VQq+Gmn2CIEdnsJKQIU8LPAgBjudj6jmwlyMnG
46DQ7BYY0xvuCD/dtSks7yKxTLPjJkEVv5cjFPrAI1Gq0ujARW2msAZAevxT+ikHo44FxcnWM5Jt
EZLNCqNPYiTMCCdVgDVu34X7XCQV1NT2xwlHVN0k8NeaOxSnBFBTZHe4yK8fTZc4s0dMfWElzKPH
IlVKmINjTmd5l9AmJhcSlfftpZEXl7GgisJtQNsOYPn99nSAjiM55T7f3iDRQx9L6VxmkD8Vvibr
6IEvD95d4rlDgFf+Cp5afYLEe7CZpVQ7wyrsnnMKqVRxAvm/0THg9U126KeSokJw+wjXYEv7lQCU
JbXTjjpaGxRljNUwOUHXUm+p4af+G/SzZK20zVuKipwHYrkABaeSZOYmeV9tBGjJuk5vGsqHAfgb
Mf9JkGUoCguYLv/EKQ6DbeXndAer5MhwRQWx3iFSk0PiQ+tyv3vaQYvzGBMc43P6bkp9PvbmBi2T
GWp8AXmwUjzsXpo/4kcRTk4gWVFxfUZO8HVkPiKKqX1R+yL2R9WSlHheBV6TvadXfsUy6w4LUguP
c3f5+os9nk4z8mLq2LV+NIsaDnsj4Mal/05TIRmkt7S0AZZNzcc84CUu1Nte5iNFBk+R0vVmL5Zv
RSHbXoo5rD07BIp9a/rJ/nGV+y1PAEIQcP2g5/17/fc7OFWrsq7xx1gVYfzWtG01RL/HweczIOg5
wZFKp1jfTChEmYKTIO5Gsrm4nkEUXnKj8qr2QMMZ2KaM412rdOSXNKDl4zkGmjlqYqZij/ecCKFp
CrkKMIRZfwuUFXEL7Wrvtcyt7JOg0BwKtNyL6HeU3sUK1vQuh8/P7A9GcVHJ7qeCKiG/g+XfRM8v
dNhLOgQbXvLgrMKZe0HBfWMs29MdTEo7Sh8HcfSnKo1YjAdFI5R8Wn+1DfnkOkfE2fMEpVy2Mqu2
Gm+88gvBeDHbOStpyb4AHBunCmJo+LSM0UtEZD/9y2SRyLp5/OjXyzN0teX7PMuN+ui6S5Tf5TKr
+qkQOhbYQyCgwaVU1py16YZIa+brmKmLispV1i5g52bjNEl4uE8gi4ZQOShQTfyE8OR6aiWxdIJZ
xZkCln464/El1/dKRKXT7hPi64HqEqMuPt8KrSlvaXCIa53YwFGMPquJrO0FOmEnlkX89dB+BH2h
ATO+p/z8xMig0Vu3c6/ZWAtOnh/IEyss5bj6MZd0Ms+yHB+DwlK8qdsfM2qaYUMVIKH2YmejQlgd
tizudMCAVTpYITmkb3KSznFKBZ1afccm5+hFiFdwT1uh+P3Rl6MyYttZwVV5WafCHspBlvzMkxm5
6IshsxyiMbeP0QLTa4s3X1KEAM5TbOuV8UdlwPwGsDbV7+pJs9HdfbKmGLap58i+bYcs4Xk3Amih
S5VO7sAoyB135WVF36DyDBT6T2NDTsxCAoofpUtWaMdDDmMm2IcrmoIsi4L4JZq2Gtbf3IE2vw/o
ZHx4VXcKufrD7NkpFPpyHJBeljhFt6BHUOWSVquarUhEZUreO0YsCy27IWfZQ6dE6RYTSKDL49et
80ndRD1J0ZZWaNNVlUJMInrqUQApqMw7GrY9ou09vSH0Mv3nRplgKpcG+4umlmTR/J5vNqbjC1eT
HlNh4kNuthPUqbMoBGnwP7mtjZRvkNPjhwhjVm+nJkT1YWotiW/lc9gnqzfy4ORuhXP1llg6mI4I
TG7tP7LucPI2ox7yTBvVUuFZvK6OxxaLxHcloQjnFtDHOTwSt9yHD3SW8Ol9bjvsdLb+RXvGb1jC
Nqb9t6Yyyb3siLkl6z9Sax/vv4AhlAZumVuIPJOVx7pBcTHsuVjzJBNySBUzpOM63HN8ctBsRT/F
xJ1b3qVnxv5wms+iacG2Bxabgm7U55DGzJTM3Ss5BWgn3r0+wsQt4ttza8LHoxAeKHXeysRL+EME
ayl2ThEzkX7gRe9R+gb/NvkCEJnCsb08HSCOi7SW6rYSW9ZwG04HbeRY4sPdBVmu7jzZ2xyw4mFn
4NWYxDD5zTLDfB/SBxCc3+JxGAncoMJsWJS6hvNregxyQ4wlUcYMAinhOQt6JQjJagD3/ZhADWUW
aCOQahzu/EhW+4FzOkRyl9f6XQS5Z83RNyP1V0splIBuhRS3BXiMHl+tB9Gjb1V4jLSivWkCaA20
fmsbg67jkZBYmPum7oS7zAHtXIgwGk1cDZ44QUkVg+K7AQBcdaIzZOq4gtLOU50M/9XpVSbEP38j
MF4q4+fRI8hPcgYXGnQdNlXZWTycanT9krqPw5CawVQ9zOxooknbJemIUCYmcxNpU+WIl7vP3Frm
GT9Rka1nOqxweGnY02ZXmTRrzauuyseuEvnYbeK/06eQuJwiWBU+uSTCk4w5ricHtkpY8liAbRfm
QVz2Z9I2JP9QNlLfRG68ui153W5HcWCQMWQhiLg9GUEM3rFnQK3T5nNWjxwZZP+RZ5+P2fEys5WQ
A68h1TSyYG5uPyTB2h7DSTH1EpAqYaKW5Iz8h/QZOvfMGIlBaiiSR/kON4JqNdxLrHx5u8922BVW
F7KnaEBL/yTYeARphXaF2a4wvEv7ARuXy15KZHHCzD33QtmTK6rHTgifDgGIW8e8PPijAVOJAKhl
WlCr5rrnHZC2D92h0drlZrnI72pVYWWRZkNGv2kmrQ1EQVAJ+QMTZ4dIyv3z2V8l27mZ3Mv5s8xm
33EhzgQ1VEL6w3zLXnv3i50ZuqmR2G8yXVfSHMMf63fUG43phyL5qD48M5Hps8LUEkbm7Ew92Oee
WkM3jhNqkDeqeFfnSK89bE2W3ukOKKRVoJxiHF6jyA07wTDirczWrtXX9bia3fEsUQMHGGI6/G2A
8HqAp5w35YD8TcvJS+kjQVXrL/ifBxGjMZwyNuNUwxTRJyRcHV6ktyON4j8nuEmfkg6o0iYDsdzd
qMl3XKMgKjK1+ZHjTLd4ch+/dI4pQbu45TKG9gvo2+tM+GWnaAtmiBuxFkhyYA26KBA0A0EezHGT
ybCd5SnBAh5tehA+dVSsE9qnxb7aYPfwVEAAIVQ6BU2VAGiRgLPMA+tWgvPGmz9GulkjHxB95eMI
gI1pPmxi/BuYNrIb6SsUa9DaumFHUlAK1fe/GaNKTXyzfqugctrr4yM/WNY0MWCxlFXHZKqgeKE2
kRcCwGfv+D5Lwm9rdnjhwfVHFVmv4Awgh665S0gZbjDRQIdQxx9jdsAtykD+8mERuvn1vht7vP5B
0lji5+Gpkc7A/5w5mGrcIMpgknKrZ4F09Vyh1mmjlCxWWh9EM9MnRBnQvrVe5UJCvzS/z/47aZhI
ZC9vnwG4B7aibYYrhAudL7SXLGglTOEdjqLcrqJyz5mhH+811a+n5yfj4s0TVq9C/w8Vuif8rYbv
Lb30qKZDaqc/bSoM5XxNM0VlmtCINsq1HurPa/qWCbGgkkcHJz7pfXTN1bkq8Gma8hXNSm5i1CQA
5n+oEh10o4CecKFAUhc4ZLuU727efU8Gh/8cdt7egfqSDDPtxu7WKiBzAGG7NWXMmSNCy/W+bXwj
RwrMJtrtSps+AZ+UYDmYpFg5WU/p/iXYID0hJddivLfUkloDnRCAhn/v0QykmKgoxVI16TpMRBEu
jGJ5CmhQYmpL5vD0pL5MHNrEDEbr7bGpXveeplE/vx6wqdPacGtimrSmQKL8XF9+xC/G3+2rhdi/
vVbOrOutp4l0jmu0CvGYTNn01cr8vNPgKTEuBI6SiIQCs9nLs1W3PYCxQI1SvkIdyTVFODWazmPh
m9LncUtRmrWeIbb1/K9NN1lFDbSSUW/FOBeBQ2b0KXJ7EiVTuQT+nad4zTLVqXLU40AKX1ABz7T6
hdTaASDMQhkN5bB+vvw/SBYaCjsS6N9Qc1uhwgnY7MH/t6J2Neb9wFxQiHXzcGnGSiY5Sanq5oXO
phSeagVuDCo0Nfow/fmF37FW5lNiHETRif+Oo5grigsJWSoitMIzrjLi9pKAn1o0cr5Wx5VfeQVA
isVakajlNSQwwd8K2aBUo0Yysb6+MzrrEBBBph9zYDr+EmLVcAt1J5QXHlXtsdtQlTVISq865qhJ
tXyIHsxLSDEOSyO1Z9NMNDgBjnLqBFoplcRvK0EafRiWpSOuV50r6OS35tF0mCfp2tC+MYxmf3Zl
bpH/6JiirxRTUFpBv90Bb2TG3FEDF1R5WF1Got/1syJjEEV7r6NT2UAvCb2mCcNmFhJ2tDU2u6je
RNtPTsGJmqTwjN4a/V/GJhCYHhpl4XhTAtIC95m4aJcO47bAdEZfinRxgP0qoePaLfk1+a+NqO62
FYoNJd+evwkcPSLW4R1y0rVSg21n2ShTmzm1/2lINrhgdc7IoHAcs5KuqpOZu+5F0Mku15tflyAE
m02BXDJNJ++jdK4BeOKA4nqgUv1XOM3f7pOn/vIslr/LIOFGOHlYcQGwa7YUOxgAcda6gGkoGCSa
tmaZo8vCk7vv/IGLZSd5LbVPNhv+675z2g0+nnBqYhWmdr0CLDVBQ8ewTbyzeu6kezYWf7f6+oaU
fB9mScX3xHrEb77/5h23MhH6dJ/mCYOXdo1PSMKmOO6eiqkdP2zJds+4CoOmtbx2qwcNrayYDVtD
rw4SGbiOiIAaZDhyzwmXEr4tnJbg0YeXu92P/QqgiPOQLMZ+kw8D0nEnPrFyvgfwnACyNaXWjLi+
pNvMRIO5NbCNEsvIFXtVSU8Dphu3bYBpJjtLV5gulNfhhndmM7r3zDxt24VmgMqMXs956miR1QBt
Q7RLlzD1vce+Uon3kuVSB70vdrPXEubgqjysXGftKYJO0b28pkgA7VH1XiLpDBFRzNYiemCWtBwt
myqwISQPmOwt6ob4D4AqvGg6fBj6FV2lOnxLyqRzCuKSJM0q1jqYr6GM8nHtOlaaBGRNY1dL+BT5
ShHkCOUkKNcp60pzqDavCEzUGxX5svsdm9s/0yEeZrVGr2JQ0j4WfoBk6pr+LkKCLLXi3vlluq6s
2AgMD2hxFA8dxgcY/7nDOvDvHPj7D5SdR3K+BSj0/9fz+KWC91UKNlQ/X2gynHv4GX05hcxTrTRm
45U4IfB5Qhm8wjsIxaPmPIJPes7uY+TRIPuE+bqr/3wxAZaKmw2jhArzUBG7m93CRyjl7oLfzhdC
rIRlLu0qL3q62iG+jB23kkXAqYzGQbHSPVjHTwOmZg/q6qbffVajhpRC+5scNbcdM7wxclIeB+f+
Ftzw+d/hcYzxqX98MSHPrRN6hPxbfYkAr+BieidnC4a+XVz16czyoFftrY68rQfaACR0I+lRyeUE
+Mgme+qbvV/OMAz+e6IHv1eh40pYesA8EnPcZiOIlfRE6e6Z6PHBIPIY3S2Qmu4wnYKKK2P8Z3K5
uxqij4aC9I5TYClK6BaMHVRqzMiPR9GvGG/vy8R0t+Sd52T0+HaaAfmVIXM8zB/sl3vnS/Y0XnCp
ajHVSnaR+HUTD74YcH9XfgTccOhCYm+mCVbiae5GZoGnC3vZF9HS9rjkHbDXICw8Ic8m+1/lKDeX
HapwC+rSwdcHmDzIgCug41KSfOBzlQjF9DRdT7YBHnQZsrsxIpNyCDppISHiSoctV87/upqmrq5g
rY13LLGXp1SRRRXbI7qBCcPA2fPi2J29WDi5lzzRyUfQmfY2bwn7oE1BMQgQhgjqYbddFFMVwDX9
s31aybP/1ReTJBeYwezejiUNdJAIM40lW/IOZ7T5tjxFKMFrYU9mlMup3UvAcoCNAkdk5GgR6Dot
akwJhp7R46ljccNE3F//6+OnRffDtVifyJmpnEXuC+gFFModab8WiSZIvUFCQZ2UyfIsmxfmCYmh
ouwcF+USplFjZw3kKV3eb10W/H3ZZIzfoYods+/CgAOkRPXa9Oxdugsb7R7JFsuaS5HZhn3t1yGM
uG4h1hQF4yWQvgD84m0gJILmXd7tU8hZq3pPhuGJo08V+QzePxegJk0ob+vpbU5vFsqHbztjZmRL
FN1rgnouYa+cCKVmAi4sfSDsFJ0JUzkXQgXrJEfhHoAifmlHtTNXMoaZ78paa1HuKNULNeD/U2DJ
d2aH4Hgba2nTFzVA88qFm0H0BZJAoYPqg8mIqUuRKWe0wHwqhkiytoTUpbybWaAOuEFNawMMM/ml
6hyhFweIarwppEJt/PslZUwKX75m9VFY03AdR6OhlcjSfPyzLBqq6kEpOxQ7KxUJBf/ajW8Dchb+
y/7uVdLweQWl7M6kjzkpuyowDxLv/CxKFt3FsbyJqEtQA6WcNJwJkamtQKzBzWhohTeFYRlkGK6W
qnbEOdQwBaw8pnG5mqn+4ZUN5GfVRf72gJRFGng5K86vPPXvOyHeAGPJ5LeEw6ZKBnNZfrOMJqka
x5IrxA0jImDCxRXU3sx0W6No6Q1w445fLlMmGxkDT15oEKKmG2chgUOzipN4kn0o9DHwScW36nA/
7RBEcgHBMVya/9h6Zyz7fupi28JyTTTtyxAmpvAukB+SwsbVnG83wSZOWb80haqjYcfhVTHPM0ck
kFEPsOIEttOV5wp5kq7sgjKu2rmRZn6yE/s85Ag/JngNpt5K5x+E/2rnZh8xw+J6vDhFcFh9OZ3Z
hjd5OlpgcSveO+mrTNRqt9wDx5cBqHRzEYoC3uPBR0PwSnGyANdWIumBBjbhdJFvRFzmcmpDNfWC
k0QK9xwbWtfsn8yeueIDdmkwNSlvmYCvoMORtmd35zqVzBfK1InwqW43ZB8CqZDGq/aRB0Hst2/3
ICckEcZxl2gqlOenAyeUgQlVOB2vJDDyXRK+uBO/wBvO5cNO/sQioauJlcNE3Jf/VeS7jCygjLdG
45saX8EkmRR9qmvN7yQAop+aUo6MXBQqkC+tz4M1ncTbAv8N8fO7PilJCHhjm/VlT+e8Q/aWYd0y
cwL3N6P34rG67sVKu1uM0PidoQhwO1Qu8I5MzXc5BZavNIHy0ZtJlWk974ufGR1zNsyQTZn/N9ls
cE0Q+rOiX86o1FhlSbK43VQV6eKita1Mi2IQuT5tmWgy9I3fUHiImBklP/IY5sIUpp294BoJ/dmV
3srnFz2lLhhen8VHZx8F8D9xOAgRUxB37+2bJOGk5ktv5MMk30ag+P7aRPFeNv3SiI3gKvNxH1Ae
rQGRi2f6StOSSKnUI8DdijiGUZ4iux6avMRCA8Sl0z5FzGgcCR6r7NkgVuKv/T4G3VdWiErwdmWU
R0cEwlNT2MWCSXuSwX2Sohe0OyajAki99rXDRoUJ/3i0CkvNBAwzFX3ie8vVUKUFDaY3kzygtjyq
N8Jcsqg2+pcDXxKlfWn71agmftYvDUlqvcaClGgY/d7IpjBVjQydedHxFyCSpAeEvzE8DpXHTa9V
lrMEttS+MX00EE2mEtIIuw53aWVjxrGkYFS0K9AcpXHM7sqH1SiesfAFtsl18sGqhkQGEOtHf1Hn
KWrvbXkOeQPWm1RukQjrgZnnVIXGLoyqTKAWxK+kmHDk5TYBCxUioDcl10bna1O/pVselgUYonsy
b4ooOP6EkiRghaW0wvC4AdUXcKedbLRIQOLpu39otn6bJVfSp+enIMfLeM0H4QJfr97fGeEkdE9K
yor/Di2dr0IfYXyAjZzT4ZzT27PtljpphB8l6jGkCOf6uqjl4yF27YOItpDW0Kt/njRl3I/Jayrv
tGw4f0qlkdoKK6g9yn2PtbuFZBw3+RVhBzweiIoSBrLUMrQCJNItkAZ++97cPoS3MXYJHSuX6wd3
Vm/jLt38K8Bxd7oE6uBLgubXjXphAG3zVFS4GU4fwakYnciKD+Xy8y4DOKmIjKxLhEu6USkdkCYO
EWJs4tA3Bzb+9oBW6YdLJeJ1o3UDocpJmuiEHIiYwIis3hkOmOijEN7B3QQNLYiFv2BdaKZv7o45
DYZQ+t78umZoN+cJh1j2LTFC5T87bAhcZTeiBd6qRaUtFk4ZBXen51y6PSct4arDwboKLnhPYz89
GqwQKyTrhy9Q1FtRORDotzSUNOU0fsjlN61Om0cunKJ1W10rKAYTuvdFjgLGxMvqY98j2AT4ukJf
1A15HuM+di8PQBg/DFa6XVxuvlqicLZSfzijlkdLk+wvnAcXbBriY6vP8JFUEKljYBFSTAjYHi/I
14ouCZ/BBb6hmayf2mj+GLdgrnQvUkcskW5KHccNtq+jVYAK3LETNx3j/K15chziQirNbebswJhd
6s2v2MdJAtqpvRWT6zQ+ZwxWrzpvHPpo6wXNO1Z6+LT/QdGNaqDaVs1l3ywts6ObrEnYE6v2L4K/
TZjaU9Vyu1CcaHGB/7sOEVWZsYjwojyPzsNnTAUA9di+EG6pUrjHaDaVSXj5O9tBRSduDBEQiFKZ
0ulm3M64S8/Sid/hrmvU1UPsd4ALbklnSpWgYqj+ubRoh3OHebTiY9cM29Sds6sxba2fElPLHyFB
f1eotPF+WSbmchVSj5yMBfpONtyQS1QcwzGrS4xVKfFdoI7GvMc7C9NNFKSjjbVj2Swn5nAT06gj
GmR9RUqf0PV6/2cfg/CcsU8nBM6zh5qjrryGeeVds28/nDk4c/bKhFV1lxI5A9H0l8FzDPWAkPia
VbBXI/qD7shPd0PiOynOX+pZNV1PkwHYDd9OGxiSlJ8mbkE65pi4m2QhVL8whPeirpetGdGUimL0
YCzCy7P4VzCpw7IDfU0fAPG5DJxDiLgkKp+0x4DFGQkxSTB1JiSJMb1IJRLgSlYkmQ2PzZrygmZb
bKrJZElVtQsOI4yzhZTThVLEZtiMyPFbc03oKL/wGcZbY/ViQNjuUjRk3ueuQLs0LilgB+1zbKJI
n4fGe1Mn2wtUpQKv92uboVD35Hg4oucxqlkX7X+F9lB4JaPf5w7hoBoPFFG5/s7SNnTF9ylKs8i4
MIkekQVTs/PqRG4rXEXYrRgBsTnun1WY/H9Ze+VdjCKEgyrm+5nhdnyH9Zac5mFDemJk19DNEHXd
1Ukh3lH4gOeorhZzqRBGguW9AkrcdnaXNa3kIax3cimU+oft/zpnz0iDS2LZRcM/sKWstzSmBcDv
OdCPKQ16TqjrwEV7H1KkpIXC0v0ff12gH4WXo14bmLBvnRsaouE3Xn5QmdjszJYIsiVLAidrfSfY
ninnYSfh37n4TOVLpExMrZcCoHFQ1tJkXyHMLoX5CyixsuANggMYuLklvWopVTUZQ2ESHzAy3/ah
8H5lYo1+lx23FlK042zcLwsa1W2vXtXrmwDlH/oWgOju8f5oHUAFMUEsSQDZJLOmygDcWz0PXn7M
pQwFMTDgiE5OP3nJbPEUmJqYwENRpF2NiJoLz1jCp+LDL9/4RESWKnLk3T5cS6srB3CtO0Z02bXL
z/Wq8KTeY4tgRVGFS4LRbJ5RxiFTXJqW+1BQ4oIQhYypa+es+Fw2pAsnHp8pzIOxHNYxd2oKjGko
j9anSciZ7/TAb5o0vo97H8Fx39vfxAJ6kUsbOaW9rKxr4rmjrG/jnEF6+GzVURMxwu1EOTFiLWyw
J6xCHnTFe13vdQIh0jrZAP+dlXdYgXcWcp1B83qImKYwbxyQJYeS8HZS9uH+O29nQoNLd8v1k2oZ
isirnBIlU/zO9cHn+LjTQmiBta600Q2C0WA+47yGfkVIJQlEfN9Egj3MgiiGPWSTBCMBVQ3HoB5G
oy+zm7Ov5U3AwOTP11g6dZEVov7lOdJ4+yt0JRfLb48tT6CTAbF22/IP6x90nqxKi5Jt5u57jyFq
W1c7a0o/ugFJEdOCIZz060XPt5KzKR+FRDbGNg/bqy86Vy9IauG4KCVml43Pv8GdI7DpLHEtgwMG
On7dM9lsHVN+fR7R7pqMgSZe372XeszgV1FoYR3TWRJEHYSN8hF032VkOlHDp31/Xs3/89CiIaBv
+1DrXRhUytewlqSHDLCQaW5cghATXDZrwyPh7DYKXNhhn8iLWrg5Y6fCXoTpdzWOx7tbYdBqq1Po
yrCjiu1/IUra8fDlwr7bsNCOB3cIlDYHf1Kxmt9jxVa0tZWL9bqnGICoK5+Ht72M5A2e+MY/EXoj
1x/33lrLwEwjMIlDTjoAMOH6oVH3fYJ+QNpl3vhrK1XQbHPR7XFQ6iu9TykyOvaVPXtYPInG3Oqv
tCZNjSIn6XL2UYkgNPPru60FDDEsCXvP7t3zTUwYgZ0zOPceT/8xPr5ODHnvE2ChSB4PafE7yCXv
GRYQsIVqCYtBxX9PwY6lpCpUeG0jsBdFlEqJkH4u/bXpct61aZwhmqmjjWV1tnUX6CjDfY0pMV+e
s1UETQH6FKMTOQZ0iyXS7M4cPyMJBjPwYkd2P9AKbBLv51u7pFUKV4lWwPiiAg5KSOPvrvsOU869
T+ECa8CSMuw/Gz5aAP978WAUdqfld8/vySMT5igWqrb0bhWGk/ENpji4sc1ELe0rpwGUPLTw9UtZ
Op8mYQ7+2vuFMxUAYVPOmNgCF/i6WpEgDKBfm3nfM7+pkqLRvDWgSB8AKRk+mkE+GpY4HyZfGeWI
iFgMOXFBt/iAZbNLvY6CW5OERHGDU6k5glkE84cfUVCP3FU3rA+Q0EOJ4Bnb8ia2+2kYHhcXQMYp
VQTX5U9zuKHZAeVC5GQtjGGXH8dGGZil3X+Da4q5TDMN/PQFReNttLnKPHZVSJPwq9oNXtKcOHuf
OrYmvXmFek3Lfijs3iE1UgxKz1XrWC3ThiKAMpCfT5kQExsHfjG+kvSzYNfwnm+zr7n4C/FMWFO3
Nz2McCSejwUeCDBHMTQJj3w/bxT5HTpUo34WVBPUO+iKVW6fBUf+DSmppzNjY5YXSeEqMGrUc+Q5
rx+51qBf7fMFR3obgVE7xQofXKgp25Vonv6y0Fjd4+h7h4U+3TY0gbZ+xmoh+bCwW98g3uLQ2hdp
9UO8G3SqjzFDN6zSK/2a909s6x5gHfgOkPo2vwSxuJ3mn80Y7bMdBZ1/XRoDox2nd/t126nKyIkl
vlvnlX/EZqI8b+yjtD3zYgYNmptBQ4+xAnOIrbTbnPrpBsoDA84N6XlhG18hbepdOFxHI6OG4ebT
AcETMWyC81mIMtNpfAehm3KxMUcDhAcVHhYtLC+vThG20eI/lwurPVBf/z0IlbcbVot6x05NoaAd
yi5Ye8rAorOHb8RQDS+1+zLJNAdXQeOMpS0O0ihHZZeDHaYBm2zGHXmfDJW27Fqo3x9ja9M8huYg
BnhYq8pEZlbx4XsZ19S7k3zubmSoD6+GI2ZrlZLJlLpxRQAt/bmYD1n41pHEflRYf0Wlcp9OUIW3
Eh9jZ54Jz2w0Brau34WSFTqvC5nodVLwXWbYMpQpKIG706ZrT6NxA4Dj+SLgadX57+kPmISyW76K
AujGen3QwLEX1EXX7EBsJINQQ91QG09eDQaKdrugWlHCezMBVj1Y35LTbmyHVythgTUvh2SgRgCH
/Tnpe7B73MlfmzoI0actLh0MMKeO+lpBP+/+T4MgxXlgnZQrq3HrRFCODtjoAVn81veSEpWzOECs
+XN4i4ZKkQ5SKAIqTMnHNp/loaQKViKglBTijnNTygGEK4surjzvACNVTWLsE9oF0MPr7qCwZxN8
DUTugfv3gxAXK5A3tgp64a1ZhrG+SC14CJZDfQr7KnfKyEbBL0Bsyx/58YKryE3czDE26DDzCRL/
9qm4CP4ZOJ3cDjxx90ZZYZ2KYpJRF/0YEpVQ61ZyxIHauOk1XMB5TB31EIlrcAINPNNjCPr5UOz+
rfREjgrwsrCU7Hj5TLMPsT0j44byqfvv/oKsDjP1rEuSJ0Esb7F+BUl2Dd+9B0I/4iHixItoB9PJ
UlrncT7RaiegNyoRfHjxl0E3TqVboAYOViDim9b/EWBl7yXukfzvyDYgIYw6gTypEhI82/tFyBXG
SjM7GQOGgg/ehSFV+bLR/Tysjto5Q7nptaP1mJvfa8zHjUolC+h/GXTN4ON6Qi74SxvxubrPfYsg
QT8fRe56oOVD5ji9bQGQCLLKaFPuC1sxtxVxLYCS6uMQ+qsYlbFQbRat0lemKJ4v9+1DLOuoGjWp
5Dm9Iz74t2NMDMinbcDT7Z/b9KNyHr8net/RotcFbxFazFBfDIWy08iPTSJ8u0P1erl8zbXhX82w
pa1iuZtMB8mbxWp4ktr1o0nRsHKFFoA/RAci0mQHP3Q58OZY5j/ALjCOw67zMXiGr0tbJYDrBWmn
ewoP/qs7yi3EXiTs8jJRBhp8j7so7jYeWyiC9nLvDrg694ULE1UytAP/PdIXyMQ6U0u8f5syskDV
LxpfI4u4P7QWIAyGRMIwWf8IZ5vLnZg2tMhPcN1ZL/f/N9W4L2iarbF1HVBshksgOsv+BZ8Wfpxx
n2InfghloXsGWXuNJE+69viANSNf7EGRSqfAq3wrEp4NfQ8Ho87CYGpylNXRusl121cqUNQEXliX
IG10r5YwpfXJRAlJszBrDFHHL9N5W8bGfAsur8iuLNLor3zmbiQLenk2DTdsUs57ljvCPda5aU5z
Hi1vJVqsFIP/vYr0/0wKRteD4BTHWUfm9vPRvZMnTJNi/T3Nm6DzVnXFcb6kC1iy65cDwB6KujpB
RtQWIpn5tTcp6qbLnrrXMW+EKNWJxKtfIRfUStdaqKbm/Mf+K/bXScC1zT7rJzpHn5EnR2HeV2OI
8se0wembO6EYugI8XlsX/13A1T57Ukuk/T1o6oXKWnKJD8+cG9V4tbobHeWS2H4Bfl/tiXKDnA8U
qE5D9pKwikFd4UgX3EIJimAtCpeFmgsTY6aC1HJIkH3mT+XyuKVNJzIfXBquSSj2d/Rz6d4ZM1UL
4t6wBzD48sF4JzxQedE2MtWIynIzQbTxSIe4nB0iDnSzFWw4EB1W79hmizLYgYKWMnp70ZfS70bw
VwAxe0KclYrtivzfRbF43xFpvJbiaT13Y0omUl2pGkFYWQJW8+e9ViK6Q02UDk0aTNe2tlESjM6w
W7rCJbvQQhn9GiJ1acjlrVwUbrIPuhN2EuoxeSKuaT+G00o2Kw1ZuYHVaLuWdA43RmMhlvMTjiNR
O8db79Bw8LJJbQMP0dFWrK1m0MhKRPPQIavQSFwH1FoSWO7bW8kR3NEOOE7z5ltszrS5OuMBkA05
VePh6XTFZOmyvaOWJVo8ju+LCt9aLhjWmp8c8sz2rogzkzSvbKVyEDbTSNfsajIHZVHBwCIfPnyG
atBaLbt6xKol+xLag8D1jhh0kqMICo1zQqiEq0HswM30NWjxlDMfsxfU7+3FFo2T/BkcT4jvj5gH
OWTXPlRN/wZNUsuolJeN4K7E0Ffrl5pqrebH6pSuut+/oYiw1MQ08SZxzvnNlrQQGl3AZF1SjtGU
mM5Sa2jtV9Xj6DmOTdf494Xt0ljBwgjGnh6D0TtOnAfais/zWE2lRxvxSw1yx4M7ZhUYm43GX8tf
hrttejcGqHgJGE1AKwDKKZIa9anta8nZ8flECgR0nQEizfxwl87aoHSXR24wYxSzXY8hmpzefVb9
tgwChG9TyKg1KmOGLrs+watkHBNBiE6FIRffIs34QTCfsl/RWRE6VVPqj8syp3Q1ug8DAL/gTKw2
zmtoETNAHsYdeQeIeZAVLAygj/eDE63hXAuxRhvfTCpHTiYptpxnlcKDJUv1uU5JcVGsuz9SbWCy
gOEc2GhW+7UUVKBB4cAt1xn8qxER42smVg+2n+uEBZhrbzk3ypgH4q7FIQScoEukHgwoRRtr8Gdi
nOx1rcJ9LfvDAIFAmMk4AWWcMDLwxSs+fUOHKINRHTPxaoss1CzwVKKqTvt44KvCAPEZPl02nDBY
gtFPqiSh0CETw5GkwpMu/arG5JlSx17lrnxcS8nXOhNCGQ1XUX2sYpKUCcm0DdkbImnfPCtKr/1m
G0lL70Yb4I7dMQZYRRYEwanehOexmlKoBdla9cW3weezYmQ40128L8+mmc+Xv4Czazf9FZr9uQex
r5CFH+suDsdEDvE8qiG84MS6a1Nn+C8L77/m6cwDoWVe5IEroRWYqfKt0QffpmVa4JEAStvwmDpw
BhQFkWLDwpwUgkBzbaF6PhVXXhimeNQ/Aj9CWHCJgXSgG20swKwpzrM6kw7A6CApv2irmRM370cL
EOWL2ELSNt6+rg+CVD5N4AdxLE3mI8WRCz63J9Glbn5CxmqcxJ0q1/o/Jku32BgA7gGgBuPk71uV
ebzHjd3Ye97kuYmuD05z3I2qfpyjn3K1lSvHLVS2ky7o5dgDzo4Ry+aOgibs5qWY3bJ918KQXZN5
BqskfHWdACN9AUBzHtr8FXfaAjrMbqWUUojX9joALWpUxzsiC5qZzuPY3iqIBgGB9RB3CiNAJfhD
XzAX8u3XMehhNEXu2Q7QfQzzos3w3fbTiDfHhn42ZSy5XXVon7ZtbJRSFASEXDRn9/6apynFlJtP
r/BjgguAn7VZXu7dSdBX1Mo5esS3d77qxTH3sE9GW7Nqh9uROndIu+3Mh7X+A/X8jsAmdZr0OmAV
Gr9Yr9tjyTdU24GZrMpCOco7Sq3zGV+bWMMqQQudvnga9O6Pj/SLTwwEY4tBj87Z7/2DseM9qopH
stXu97t+hIOjLqHEKXg1/2LbISjiQGA5c2sYmqF/Z2uT0Q3s+me5/dvm3qSQ+OPD5LPP4qO8cmX1
XsN8uOPL0jWeXSh738iW6DqoxSlZey0fR4Uv9ipAh0lTj0Rls9ljI/Rpe6TVt8OtT51t6rvNcxcj
eELlGjsEvJ6vNd+Rg3DB4AkotYFTrxFc9YK4cowh/bf1+WKl0WPzMqpes5wxMmID7LTNKg/B/VPF
74/TLnXvMF3cmaWb1q+JmN89SYUPEeg9B2rZOFD9Zmops/TQnuEFedGbr2H6doadIdhXyXZy5nbi
uEEI+bhbBXXQPsdEaKvrSCZVbSIVCnZ8byoBUm9hR3JpFDYHeP9424uFKkq16Wlg1gD6FkTWesQL
bLdZSA9n3GWXDqv69aZh+fUaBYAfq8QTUSmo2HLwW7CleIKRgCPAmn+TD8z7Z3UdG43jKoPMsEJR
Co25xiB8lUgeExThUrFLU2q+sEFWqg2tUvpxc4jLZuvAYdBTFpgYtxB7jeusUB4oLex/PsTQd5wA
LA1ef6j5AS2vM++MtjYSkV5x1UycOHtkA/f9sKLymAu+Io/aPOukNAvZp7vd9WwqH9zgpSTRNNj9
vKveEAc2Sc2IxCWPoqWcuYIPRqhNJWrqe6q9bRs5GS/AJi8VLyXTi2YxXH7qi/CbSHFfoDfqb0So
yxxSpEDRV14SydtumMR1zeF/nTDnIYfPQKEiEjfrbg+cfTk/t38eFQw+BarO+8W4jkEjEkQXcdLH
aaqTxR1Ek942sD9LOOoSKwqnaEihCkzrbeVriFY4t9gMyak+nuYrOq36oFUUauepl8rR1zdXPLO3
7Pt4sdejrxRAycK4rd2iQBu89t2dxb/J9hdcDSeJPQfBTdsaDI1ZCRUUUQZ9RU0vIDIiQH/Hxj85
CxBy6MhR5lPDEvbqP6/10Ec4w0pXWZ7miM1HwFTLCEAa/Uhwv0ZF2L+TKkMS4i63RH71gd0AY8QP
P+TPlcF496WFb1wIiK6TEYruUY5LjzRzcKXS3FXKbcfnwkjhAQExx9xXAZXScEdPTuPAWWQStEKC
BUF3rlEYK3UiQAIXdKvqkgS/ur3J2sHLOeRUs0QtGvJRhrePBliS2TErx5cuecXLggKNcy4PC6af
qHbU7kWIpEGALaG9D+4GlLIP2BBuYVuYc84JU1QdYPHMXqDfXNz3Xb6lFWRJUvH58Xc8UMm7rogX
uvUtXqVCozNPLKTOE6nYhNao349iS0x6FMpqVGtHYIt/NKDpqw4eeXznXFdIqxyIJH6zOgbzOb+h
yUC35MHDRmrIBbtSpDYevs3htTLuu995Deb35TVKvwLoNmyOjiL+HAJ3388R15deHrbWpBKLF+y7
NJknF9/ZMBjVhJCrJhs9lyx778DeSwCkffpn0fCeOczGj56D2xJMPm/XxYwFdBQGy4Wzm7Y5WJCj
nPXD65EgK/lMxPSgxIMggqiUEpMpfu66gingw1zdH7mBzLEpU+A5hHjf9vHybGdbDfwgjfJe3V58
TAF76S4pMqVuvvIQIufJBdmr2bm43rvjUUZs3cSe6i3cdLvy+MpERK26wYqjldBQA0l3XE50780+
sdOe9Enkbbxd8xWtS3Cr3CnIkJmPy/E8EuKstjMcOzf10d5zIFg1405wI9S4pY9liIDMGY27dAFb
ghdX8lRguyq7PgbV7zmFTw5GPU7ojwVUIbZFIe5wDexQUsgk8azUhaHeIVBW8ZIEYdX4d4mSYlV6
FG2LxVFButbHvjGx06SQdb7Ajdqj2b0Hada2dSSIVz+7Blsc9IAXIcVHowCC2yJHO8XyZg8BpZvq
/9cEr4wX3yI6/4Wa2HRH/5hMdCnVMKvxCcsl+6h/ezjeBRUTt9Nnj2Poq9bNQwgLDxXBD3lVIMBT
9qd+fuTcmP+Zq3x4R4LVrUK/4mAMGwZE6W06UaC3qkeG1KxR/+j1WngBu/Iw0voZqalrS/nUsWrK
h+oX7TtXDdBv/PuObCzvlTt/EDJXzv5lkCwZ4o1OWRRUrPIr75TENU4EKFgQxdXurHLj96gmgXiz
QbPgQSunyD0iY5RZej1XWGuATCzhjPfmQiNoqMpOScVO5wGQGQRaWQ5rh0JLtkq2ZjZsMDTyZW92
JPTeWX0OvOMMFE0diEJtpgrQA+ArI7TnJl5bmsJeQgmKTZ88MDKT4SINa1lvCxMnuJORmWYGQK95
xJ4i3wjylxPU7Ni6Xs+hXOqF8wIJP6MAe4B30+/2kwQ9u5EvBpSEaiQOPOlEzJhOfzYq0MyJKfSK
8wNxUfZoCEQlzU5fg/GIUeEefVJ4AYUZCK2tFsTp4pQ1YvPEt8eVPpfWZpAC2fkRWMK1LbM84WfP
jqgPOcl3Umuab6CVbmBcsGYOwg9k5kQiJXg1qRNgE1/G14+ms9q6/0rjWlflDVv3/56Tr40hzDSD
RJ+iFCowYorqglPyazX6M0QYxMJ1VpMy6FDeBGi3f3MsnPHEi7y7A+7J5/vPzG3H7AHF2KioORtN
6/uXFQRTG+K2H+1eRL30r/gSeZN3mIq8AEhm/ROnF2y5FRpT8h7X0mz9TEa3I0SRMZUbBP9wZ8rA
9fUF8qgl3O7b4K3SvjdqCMHHiU6/FQuqgikC0KeWRLA5XRQe2eBt+UX1aa90v/c+Yv8V0DW/aLxD
22q7YZfMCt5CIMhTrvqF+5aVOuMTCbWb9kOvooiFYp9LYRely9JdR9OLdlb/s2+w93Ifjwl4cf/y
24p06dBPHiGyRObx1gkCqO0Wlrm5L4IqU08z5wo863hKQgCF/QS6Vpwc5vb3W+Gbs4Did1hT5Vwl
xawj8ybHcRQKRFbC3JzpuKiIUg6ZlhOCjdSqFyY9/EakQr7wW3YSrBiAEKDCERZ3MuopM08/jRKW
a0iChIVJCh7RXnjAPvGT+Z3kXu7wWEc0tispn7pL4+QrsOQdAKhtKy/94TiSOacRWkXL1DWyD6vv
rVw6VEeUkhWkGXgrCYh+zeZyzaCjVE5LeeepaBpC9511V6Lo6IYxVj3TQwDt2ALzRkT0muhnhegX
12X8U2blhZ2Nfi1K2eLV2l3TXW+XQ1w6DjrH9OGXyQN+gDC4HXPXacrTrthS9uIDXanKuxUX6FVM
WYdM1GHc5XRRfBjiPbooymPiZR8YaO58G3gvaQ+abzrrl91jA9myMFgTKY8vB7MxNfCTL7dKYAiN
LRChlbTeAdpSC+5EqZ6O4M8cowL95/7O0jROqZMq4IE9+0VpWPvyrwrxiqFOR8RP2Hc8urttYMXV
pBafTvgXi9OL/FEntZmZwnhSpundoTjl1IhaOiDinEVubgZ3eeyg50oZEmu4b4DmbdD4XwIJlHQK
1kHSCsk5GIBE6UmH/kPh9Yxby2ZR803qtPSFtBFgpdDtngLWtGCMO7xmRodfb/TYjtl5gUXvNXg/
+jY3Sz3CTEiZqgDAoFaMzNY2N/3qqwa8PfRsHsWIin4v2MKGFcFV/H4t7saLNFombtIdwPnsha17
gf3IxH0NDROJ9get3RA2lNyVvW0zyEGfm4gnh9q2kTTaqD2yhz6JDBJUXIaSZdquZ8C70tzIF6Ax
8UV/qJR90HjoWPrjQ+wLKWjMgB0QcSESi75mSWCl0rAOs+RLFJ5E5Mpo0bZAryEpWYw/2bJh6xz0
tMk/2C5mnebZxFcP11i9UVXy3q1cGF06VVff4P58gwmbloH/MvIMk0JHWtdevYf3s5OaPR/Sznuo
RJRgqGL1OZwHkzhmS1hqxS48nTRaCWnZo3saTu8HlEmViOQIaqAsmda6ZHI/vUpzKhmD7GoxNORr
6m4IB6SM5fWoDbpLTQ0j9p9An+JnrPrMcwBJdb/pBlmKsMhhYD03CcVhP1TaRcIoA4/d41ZmW/QN
5G7I/gXs5Athws9eYXtSeHGzCOic0TEY3bUj1Gie6GFkB2EKMsOWJH6pbP8fEgztJiUwLjpTUK2y
9XI6Bc+RIenrdpbuBPDYYTspjx3zziwy3HCR4rMxyyiqAhliLmNYv8xYxF3MNHoNV7K+OghBB3Vw
Mu/yEzr5MP47TsGYNZWSoYL3Xsv09vW803HQZcMv/J1MpjASNCYfxNHSTxTvXBCm/glRejw5SQoJ
j0Soi/edwyLx1hTzjilDyb0TvxJI14aGWDT2N9dM3HaAIbj1RApIbyrh3oF4S/7nG+KzhOZVPP1c
c8N/ol7lwwEyWJ5Gxs1KyzSHGrBiaoug95/teeq6VOfhDWzPo4DT0Ws89LEA6f6ZGIuob7JHKzr2
eTCm1WIxzMvmWO2FvZCE96KKHZ6JxFIOkRD382C6wgQZi+fSlFziPUKx15sk7y1Y5OhudDRLDBAZ
DktG/DicUldH+lE3joYOcgZMLS9GJexiz/sbDpkf9mLTXrWeUcuYtUZPmB8I44KMJjYC0sKIll0b
BX7UZDGYxW0706JFQktZr+AVe2m59ymjJEgCt56DlQldl63XCcZibYnSo99/FCNu8662mKZ1mbTU
N/9DV7fOqHBwdhDHxehgo//jihrMtNS/eTGvoSWmPFgdfkg+JbeM0wMDBTic1oxE51yO6ty/yp3O
FTf0BKPmqPHkJl7x7MgbmmIP6FaUxElWZyZbRuCxkKwSC7ZXkx4rbZ4NaU9bnAH/g6Ooc5ReMyZu
F4g0dpq2XUq4hufd0K3jBagGCaz7I/54k381WvO94jTpnyMz0JdcQBH61x92TSY24H4fdMitLcEL
r+x7L2aTdUWtudNRyKGBjhs0F/wJ3R0s99wRBPh6WlrroD1cT4jRHZHrhPt+HmOwDQ5wdQw95gsY
lWDA2g+7JT+iL/OJz2tzPEtpLM7goKIgxrCzBR2Qz7UzGlWbshTU09Acx98I5jt6+6UJX5Fiy1r+
iWwUD6GyP1wvFEspAyBy86rfimrF2oqCmbMlr+m5w1pY2h0y+ARGWmrB6d/DC5DC79uxDgDCCxp2
Qa/TGcU5am1F+gh/PG3HxLrbePfSBGp79Mh3BYvQU//9ApZirYsWdM6083c7vhim3pxiHkvYQB77
f4c+G6J8K9D3P8HZ+SSIX9PmnWLIyf1GH+d6Qz4mHIo7us9Pa8sZKJgH0vYMxPsQzH+Loo+t+6y+
WHidZlGlOaeMepjHZHxGelGxf9wiN0ELRxpRaRQKLaynvTW2mTyMQorl+pdCF1Akn0d6ZaQonhbM
LwbYQQwXJeKGCYyiEuNZLBJuNr4LyXUQ7pc4z/TZlun7fmyiIOVUJEvdMcuYNyRX9nY3AZOhWshM
jvACS4TIuSLq6563zxzCdQSqzUNNKdbE9ZZ2p4TUZ8AsTes6K1nIU9SdESXkXvo8JDFjYB9KPqOS
Z6Fb2nGhZm5eRidCHQGxCnmVBSyVQREh/TBEjvtpzIUFy1GCd1pEtCfCj9AEhA1wVkaQSVILiini
U9UY+D5g1xf6Paggr8QvONmzfG5uWBA149QW9pay4PixiI+2varN3b842qmg7teaNq4R8bHO6OKP
SyZWcg4rN/2r0C8jYi/huKrwW6RCTBvO7fBvUWgLnhgx7XPegcAYB3nIUW55EXSfZeJrsq/jzRRW
baBEKvFjMfiycE/bCIZahbmKk7yvyEMALsn/nOhD3xRh2Xp6JpYZ1oaNxlV80Fk11lhIw55pwlO2
zwutO+WDp9adatNIu7HtbqHYWX37AjXENOsemIu0eXkeGbfwLczFRSBaiiFNQcfepQze6vz4JL/C
Lunk1suH7uhT7okwe7Lsnhs6bPAOutFKd8UYYqSHO+X8wjDZSgIEdWUQwpPEd5Zrkut9xUIKJtnT
TY1+9Hp+HlPcc6KTjlyv88jrcERLgwsZe+eoOu7qSTuNSTiP+wFRHelWHfT+845K7yfaY2nhOTHL
ivH/ZgY/LW35LeClTBOWF4GBdZnQtbUJIrrrEx/gEaVV2+jQDQ/gMPcl34VgM/1DSBChGtWIk9sq
bs73OFdLn4PJ1WmYIRJUxtShYeZEDQARs1m8gfbSQhwnmPfMrOPZb0yXzn+oXZNuV8zR2VBdwrA6
8X9LWDsMOGs5Hf8VQvHcVk4Qd/S6qaFVNrLG81MKWr2H1CEcxTrArVtQa4LdUVTIQtbQofkZZ327
aJJXW43sdIrts90Q4Reoln2b4ixE7gPR11Wuw9bR8DUHgk3093mV3xPrXfTUeBYM5Db+eIaetWFG
LCH9ZPWylSSwpmzsF2yh5YGfGdwWUhoJNr9YRcRU34L50iezNxN2n7o6ZoNZkM4azcvBq9QrRY2k
37PDc9Cn4GUXc9iZsiIQ6axyCLmx1iIu8/YzM7i7bOH/pE/slVwamb/KMQgG0GrFXVe7dX5JjslB
Uwi2b2DQU6g2GP0IeWRBxe3BiibWAnm0eSrCNnrsLea6NqHj1k9cJzXLy0XcqjcEkEHZdICCeyLt
ih5iKlcLJvhB9xlBEf+cD8ZZ0Z7Y4md7ruJn8fPTMO7CQdm5zutTqv2nfWhrGekxnXQS/ikq+Ijz
5UUMwmVyzGd+rCJ7QYijGO3FlofTU5+aSxsDMG5SmyoBzmN4HH+QULNnPeF1OPK8jo3QeT94A0Tm
rbbHriVeFpuMNThOa7InIpsUJ4AmBJYN75V1/jCAO0DAXr7RXjW1tNSGDwvWIAQXub5bBMv9tCQg
2KBJCvwM0BX0ZuDDFesbzSGvLzfkOb4oWxbgi237HrTVZJoB4VAviyUmCoq7fJBboaFVv55aqajv
si64i4K1TYwH+Otvjlna3gVIR3gA8xPSK66a8i6VjELaBzE4a0z8ltWUWtK4mP3h6Gu5iDHR69oB
aLsuq/GM2yr9a/OgkplRwCRSCgMLDcLMrSvB6Z1JYxjvnOlctTc6DDmfAe7V3Zr9s2q46OKiDsam
qfgARNPusDizp+rYDUENsSGv3wAdaEyOhlMe43RBLrkcJtZm31KWRpF16RGP7oARZny9YwSR5qGk
4yjQwFS8ydfpchV+alzKMOqU4XbXZ5WeORCI33Tg6x5PYNIx5OfnShMTsbGTX27luLFnMNmL9c4G
/TZj9MVZSmUdI95Gk0obDS9BeAY9VAY9aReEK2ouenx4TzRsilRalB5aiYW+YfYMQa44JOi6021o
3/hwkFeQGNN2HqKM6PhNtaNPIIf9V7NYAy+RYMAANWZ+YOq40LnSBEDvleFRpn3mWj2Rpx8zlC0i
skRnJB899y6IC9lUZ3xqXL53aHgFtbtsZRovUZwobhay8IpRXGm287dgiZg7U2yCgwK6juhFDaqH
FCe5iVnhheNelijgUWNnCCITsmlqnhwA7jpmPVnuALnWjOcK3FKyT8Erfncxzy2TB85qt2wOyXGe
3s82bXku2gsgDcTF++V2S5c6bN3HRO8lmV97RRMwwKfjfPnh3CcE06l1kaHJyydSUdGMvSyCy7pj
Tie9M+kMyY6QNgJ83TpOwN/kRXDs7qOOilXCGNAmG9o9Fdm4tSZyHRU9NCwZVWIrq5S2L1m0udQI
XM1AFc7qVFcN/d01WHuquVXlBweu7cJNok2nfS8xSKZYbfkNLqFXnzED38Jw5zOlKpFQH/BU02vM
iUh0Os/ol05yne+R+dG7s2bhpWpSTAEe44fT+K39UIq4I2FVzb5QBA9st+wMFBsaGjOiM7cuhSkj
QG6N0JqJDRzufDmHVBfuuXgjaJJNBXzZpHJGumOvHj6RgdCI8kddD7gFNvu9eQpjLcePxtBwc/O9
de70uRT03qfh5SF63obTF4XBrOKRLPxWRD3iqozi3Oculb8lgDir9PF/Zj60zb9lIRpQnKQisTwx
YD8fiQI1/BsSKT0x5sgjnjiHHbWSpamg5279Wx1fX9OquEn+yyArSrS8h39wL3EMJh69SQb1YHp2
cdhV3GdzX3XNO0Gp2aECkGKSgyGGGmwh56dBm1g4bVRMSdqDA2YbgzBXdFy9ZaPMnZlls5bqC0tE
O7LF53h+Yr0m76pav/AUtlhO6ufU49tRDvQNdwUTYxcb60j+aSGIhkU2NTn8OZfM/+v3R0WufbDA
10sH79oB/zYppRM25ClQM+saZxBjFEtgrlJTKpjyrDfUeagbPnjqeTibxlH+VIHlURTdl0Z0SKBn
kkcVE+63xMOTm03DZw678CkUP1WOJ++i3zDqxJyKyoeX0v4MQykPYneS8vPgqnx2Qjvx7EidEe5a
XAb5gykqtp7X7ov5GHXhcP+soo2Sd0PZ8gCxrTcMPTBIm6yZtpRKaCZn0ni+o+G9/rlQuubWRTK2
iz7Df40ZpeLsMkXwhwvil5Yfv/dqno8a3MbIFQfp5G8o8ClTKXMfZHW1VYfh4T4IRZ+JgmqznALt
N9/43nkFGA2rxHA952sbFv2292ll9RScEpJ2cScsCSsHeJf/kwoamtsrAtY2qDcktRKV3hYjw/Dc
KYqrY29SX0hKodoexfml6/d2GFXVwsqpR5Bn8Tm3xKKO+JQSI16pLIsxdpMCc6HhkZNn+sEfEdbl
b3bZHrnN631GCoJI5nTpYLHxPTPDK62d5a405rVVVLyEY3ln/iqgMUYrBTq6xQxH3g1z3ZG8n+vT
a72Eu50WqsULbaZ8b2eRr8ae2XQBQvBM1W0EC3kP1EBnPY1bm97w++EIzpPnpVkqAdnr1yEfVyHm
aZtVZ9Uo8NAXAG5WkJ1x7IHExGtmGrM0QHS51Tky6ZSy6voZEYEy2itq9Jdw9MnN1GyV9Sm4QzS1
R56LgXX7qTtLJxTkw46IbFdo3zxq6XGEj7EDSILiJZOb6a/MP5rN0a3VOp1PbV8VX+XJU47eMJeu
dPFMmIQGQIr6xpLvsxP0I9AkrctxcANIl3v+MdbLCdgyLIwcJreqptqpYDv3/K4YNFohVMh1uzqa
OwWV4esn5zaun9/r27xDj0JhPqDWU1CF0O8E2xSOeQy5J0rJIwgbQx2LQiWzSE4dzUamKrjnjF2r
bV8xkFXhoIj4vAUFPP4cDPgRA+nAtd4E/FpmBohRcJC0zphAE37BFrNkD7rYjuPcKfT+k5Epp2wQ
cRpbQEOMiiYpGqgMmM2BRWyKE3uJExUjMps7ndEWsEPE/QoZcWPabOSwd+tNZ5G959+37AZxb4KW
q6KmUsW7XssCOImBGmbkNYjBLfw6l3khfjRBk5Jg90iTzPN2HDPMRNiL7Zp54DWkutJnGmHl9Tlu
N5h0qlK6u0JNZ12AJQdDKvTmOWPSQqHAiAwzTUujALq+eScAyDRicZzB71ZDK8hroPIlIQTqa3YP
HSmcbSC98bcHM4tELDNWIofDbOK0kaH/lKJk4C3yfOgLzMKeKP0i4Iwfvoh+jUDROFCtUToJy8Xi
zqR7flh2bEX15AtXIX+lBwnUmgkmWZytbCTtBXy2UhLILR3lDW7CAzb+FJEgfWan/nvUUwBKaBlo
NDgVkxEEDu+olNUDUHtPwbow9C5AbVqPeKt/lbJWuPKMO5aeAKVaJeyeAeS4Pyg4lnsVIPgikuCK
cyXL3aXYxgsfglHEAqTeOMD0tWWcxYP3Pr5at1kJpuyrF92Lsm8YEe/0VyoUdF1xRjNc6nF1LZVK
PbBR5t+JlP0oVtba+p/fo8Mu5IJdsBMh/B0Hn9Bo1wZF4gj6urcKNNPMn9806jnQqpU5VeW/wO77
g6ZI9bplustpsaJOyT/fHNjOxPcLDiBCLhls09VBzlhA/XWrX6ssk5NH3aSjOkt5oJtSLsXG4nQT
6FvyjLs0Kp1bYQkM2XyNiOtF1rhY1gm+mtZVNmXoSi+TGN7Q72mS7aQNDDG4M8zp1ZUdoZnZtPqZ
rq+PbeQtSJOV6wjJvNXr7dgUIbg+9BbFnMcq8Vlu3OcnnS2dp2j16AD5SRdWd6GY8ghiFsSYIOtL
2K/9/ZJwZbeEfV+/lzmrUsP60eHLXaO5O7csc/OVtaM+Tb+TIDTCj0ZvXO6FTmICdrOK0Jbg6PcA
v/VVYxtYXQTmCP1GeRHtZp+XtHtbBF0CN2pjromRBzOcsZoUuDMzMBT3Gmdq4YDYquOGjezOi8sw
766cllNFRU3oin7BdQ2+8vAYXNXr5NXCAbPC/D4hHYCM9xk2lJkOaHWrRg5pGTKRKM5p04ICFFY9
JPKXzfWhbCmWJbFbiBWHyvx+fnILg5Tx+KPBty1OpPjBS98Z6X5WlgQpvs3dnP4wnZq0SyXaR2xo
E37nt++i/ELFYndxHOm9MEIWb9Sj4KSOgfFhsYzGTIfu2kW24HG0xzBaRii25Tarwsns3+vFoYJE
aMEwy5rHMNSAUFegrvpfbaCyqP7lnnMR2chEhNBN0PwwRjD67tknNBvE1PMF4bKgkeqWOc14Kjly
eMTrZMuEhToVUTPzZbOOp09SKnnBIwyrCr3GqbJoMwDkGxQlUx5sMyPMRbS1KCTXEWs4L71PNk4A
mXD7yO2tSrNKB6xc8N93Is+BmXXotAsLgCl9IE+vZg1o2dHFdRdsjWRwna5CMgmgCee2Fy6B4Lg3
G4BDgDsiGL2oztfH1UIInGNn/tuSFQ5NGtDIOIPtBdzTDD5QhFyWba0e3ykAyi9Ng9mRTPl1NOMA
aXzUDyS5IuGXqJcHM9GkuylFN+tpvWCLdELHyyZRZNXjiK2ToHzQY66ikvqORQcyRx3DRxCvm04i
xPtID7iWEHu3LLmHortuI+Lw2vHBXnHlKcCA3C7+oc73e27NtOAXHj2IpXI8+1tZ39vGcuoEi9Vt
bs/6ZgpaDvFZWQBS3SIWURTGVPqjE7JWRd2nICEFZMCKYwS9OHXR3t4fiOVcvS6p8twED7IAZm+j
z6DX6KrxAoPlkN6x+RSkkrMTAyyE+KeugO1xlYgyQOHW6hGTVi9i1akZ8xyzMAz2tT5dEfUjfEAm
yj+An5OgmUfa3znOG4dm5YfFrultSxefWyccrXYuu/23muYgYJgtICj2tIRIyfBSgohawRN2f9g5
X9i+FfcK/6RxnGxWgsdsh9Fbpe2K7TIbToMbHZSRRrwVCic9J4QJIDIl6131KNME7eOVOclgLJI5
hQd7GfrzXIbaZaPFHjQIFtCWtevcMm6FbYuiD1MtfloZKjjOvEQMMCsmV+kzEeg+X7qqM/nA/Pgz
VGa2cqPmu3ikpqp3L4wbI/adylBSxbsrX9bfMGy5yXBhRZHkQVtt8xo6ZXV6M2GupEmaYFSGKNX2
uOHfiM9PnQBKgQ7Bim7n8X9KwX8lvhTmb+fYII8qj9TjSwJKNT1+jXCK459ITn86sfLK8ukY+Y9z
ojmkj6R8+Tkng4mCsO9+8AHnkCbemgcHLPacHrKSTqBk9FiS4Zj0s0fphy6OfuwmOjLBrUIMVV8V
uV0eM7bZzReuW6O7Xde9ZJoBSpo9tG7fDZrL6ihpD8vQaxe+lsl6kccJIXyZOSg+Ee+x56GoS2Yh
ux4/uup1Q/sZmcfbPMVN2Pkt8a5exfa13Me07C+oePnfCIjzJHJW7aQpm9G/GQxTIHPiqytk61kG
iKjO6VHReCW0dkb+nKZzck2q0UZRZ+aluWHrYMfR+L4K6/k0Z8QH8XLTwUyxycbBo7XcxE3Qq4F+
auTJNqyUk4Kj+7lZGli5AyGmLlCj655TTzUF3lK5APE6rM7W9p5+qDseElaZLHZZhkIVTRIAjJx2
yqRVNrGUOoRq0DmMfPhmwne+k+2BHJpwyZtl+MTVyJN8scY/HbEwwVY1J4CMrrqGVYobspcvWGck
Mvzkwjfuc08HHDTmVL7bmvBSVPp48i6X1bdHtXMaMx9L3smkxvM6daktrgKCvSLXxbhQ0ZtKl8zI
Mh+Bf6hXfvxGlbS9tgEeHApl2UPsr6uC8feq3GcNJes8vZ3HHvoGykBs8GkLWU6IWqOwkiT42oHr
7fZ4CCnImePzuTmfNf1Gr1xsJqe/WmAYgfBAhKlv1TOMUDFfksOMnHoRktPx11I6l2Ft6Hw7jbYS
NYhLPE2CqJznYYec+1luG1RlLUocdzGS5kPYopdxvnMY1kg657y4we/55J4S8fe9S6eX4glGD9J7
CrRraruN00XAPfgnHeO8TzTFuyYvgnshAtXqT6HdegnqJcS2zbM8kmR2xs4XiHOni2vb2AVvciS8
/ZRRk9GR4ifH+VmCDABPAHYjE35yPcGSJ7twGFgWbZuMMezGQWRsPH//4GsCFTQI7FQZ+XC0FSNT
N02QNjVoxSW+c3BuGTaDz06N9x8SaNd8x1h4Zpi7V6mQWqfujMoas3iFsE2Zxa5omE878Dx8JsMD
+55XbzUVi6WbBSflRP6CWTSXQidbDN3BBadF5Y60y52noznWdoIBus8hgyzykUW+ewVK/bhSMJr7
Rf3Y1hL+8G5MSGz5jLqKoWlI1OPV+aLRljAgBmckDtUr1SavrK5tOd3LbefPeSsVi+hMoUXEOc5k
zdOxN6aV9QvjVOH3x34L48YYFoGIkcp0pzrUQf1/UlWQDndRx52NUunvIZMwM7ac7lWwPhFTpLZ3
ZiYGKA7VMT/aucwxHYETiXriYuLwQW4sCMZ20RlRPeDfT0yXHgBLRwxhMTHpdxBQIGi1nez7FHt2
P3lUQqugg8/xnzmnJWEF9TJoB7wDPZYE7XbwlnL0x6kZysHHCGEt6qtgHHEh7ymhzpaAbTNKJV1w
WftidwQW+BTSCSDpd+r9USWfEqCdhmuHlXigkrh40f9JSL6PcjEoIdHAH68UIDs9Qoc1TOz++3/c
Hl/bCpH/g9AapW7W3TA5u5hSnhprDGMa+ZHgnsAWLYq5Q7PWXrwV7XC9B9u/nnyhR/5UdJl6GEDY
+IQZoeaMQ+esMUTweyicrIF4MZL00Urua94E1diI+jgH/wcmTtmfXCe1xaubVf7nQfZlwtNUOKTy
c3J9izw9nY/kw6JpF+m5NZBRpel2iAOzbEQil0nbGHsdrkDCu3HqmubDbYhwURlUli++O19TxJdZ
zaCGFHXwI7Z2SWW2uz5yLk5a3ZztEuJZO3k1mYGvW+RkE+JIIkY8YhulbnadXVX0DUNgE3+Sldmd
0P/b/oE9kv2kQeg1EcN90jqWJJi5aurERMPi/plUgqQ4UKsSDWq1Hy4pAnH6C0cKoqk64CltqwbQ
7Czl0gIQw4AouHqkzcrDmwA0DpbQ1VIniXbK8oqYY6KtgFopb+7PJn6frZIyD0phD+7U15u6RnUJ
Rg/XZIH6GoCt6/jzB/o4UF8o0ibAmx7SVs9cVLxcw3YUSCk36zFvfb1nxy4IgKvPwWatGtsBKfB/
D5g6PQG9hzS5qdRMWfEUlKT4LFPFx//5dVF7GVAY9glL1uTQ+5nqZ5XU/VPGUDqQCHxzb2pRbGdX
1nVO5XNAffSR8l9o73eDT3y94bR5kP9EaCFvDsvn6Hk5EoapGJ+NnKbi/J9FEgIVylM+WzdJitu7
b/kCFc1igj7B0Q5VA/f+ISGS7bM7oxSsgrsHpgz6tcgKNE5iwymc7zCfDuQgJEmYfg7uDQGOjYbO
67F664rj/UC9VupV4al6PM81o0NRn6olq3G/zseogoo6JdaRmxFMemmaaOHQGjnIZ31a76bXyGTv
STkxa4Bjf35kfyYLivexBxPa3565PRMnmGMca9wtsDwSIJlTvq/4yemUwN+vxK757sYFiwLETfuC
lAMS5GqUVwpXvP9s45Qa1KJfDOfW/JOlpchWo7ZLYjAXW7AHs/PFfQpYxPA3CKdKHm5xYLM9iJPR
owU1ePz/S9Z0b6gvkmh4j2xtKuNOdKSzI6drwKqyarSke+6dhFrSF7BGT0jmf+DXLmAmREId4ALc
G0O+u3Bg6n50IWCTKdVqTk+uU7/XMNvyWynGs6WlcX7OXoo55FbtIdE0DFXbBUAJWp22RXMqivfK
yGUHg/V+Ix/lsaER/Wb/z4Iy41+5jDF4WMZ7+RUT/3Zn87t2ucP5tRLrVia2fYiw44Se7Mocs7os
Hj1ln6IdEyVh/xk5/P1pqGGelHUAiEATYCBtA2OOGhGo6uve1uOAEHKZDFMJJYkn2zopJ5/tNF+o
vvOfOMV9wKBbqNC51GLB1SkXzdy7gB9kF2sg7JkCzMXZrD+tfsJKwzlmOxzP7Ob43+LQ/kJRjiJs
rHzDuHoiEqTopsNRmn3tu9g4gBVLU5vAyJ6IpasB35jW91rRCBc1G/UBj/slp9hhitX8erWsRM31
PyelWW72FDj3q0DzS4hJJtIkikeUD+/Zsby7S4gCdVpWueLj1nORQt+a4aC5FWEcDGbAUZGB0Rn/
5hpDEXPRL4uO84lFp4QKDnGSDPFUHfFjotx2H248V52p1df1U2eZG5rMfl2FnhI8wd6qTtoKhRBk
PK/tTg6u7e7uXslu+CvIAtkwesdFARRJhSSdiC5fYi54p5bsBiFZX3IVGhW7wsv+p85rGTb9wJlL
MQvEECz4VCtOyQBIecG6Q7xajlBdjc0/oP4py0GPmImkTQbpSdwv9H8ffQGOQpeVudknWdAJIEdV
Q706Mu0ECMzkMsANp5B4yPQ3JIKyuB9qloVQxCknAYUyxmwXOAVLMnGrQNttMfxZnuS0etS8fQGH
Gc76tVwSGUANfadaoPuHwKzwMUnewCbMueMWm5W+KYzmBVhLSrcvF0niPH7dBh8+lw4LFxUNcJDD
vHkKc9cO/QFPqocXfHig1ZAVwUjsBaYkDtDZZ0eDjd+K38ak+pfnWZKpRB0e5Fiz6WRkISlicD6r
qXJ3dO4+2/WTxS4CK36z0Qsl6aBkzgoVS9uZWOBcG9+QlNdiS3TlEsphqX1P+upMnfmXY0C22mvc
A7SDqaGNF5g7+Z04urYAJdVrbcuqx4SKxZIM9xDByvLVm6E97gsGESeo2OeHUqIGWseplaVSspAw
Cj6qRsk+GTJ1SAAQFvef55bXdpCbhny/V2dv/c2iqIw3fPCo9Z/P+VlHH6Umb7KxDZ7+Qgzor0J9
VFYUrlSnZ14sNyiykyBqaukQUZua7S6EotZTAAN4sOg2HgUlk2noynyx3B+JWhLOQsWNDP06VH8a
NlTPKFjdWqB5QBr+0ozJtVNnBt7NcWBr1RGr/+QD+P7EgxSl2SczRpH33VxRXeszYKenZYKNyd9y
cDE6riPjtRZTiMAMeEpys3cWu3JRpnqY3Y3+Wi03vdnALR4u9T0nVVfxQ8QcecVLTdardDbY6PvT
Wf60krQ19/cSjfETgjiAbV39sJ/R05G6fdAoiLb0j7OP2EdZmEaVUwUcDPONWLbrHe4mOMp0165+
7o5YE8EERWVXQSOojRp0YfFNLH3LbqcCRaifnn72JH3dSpDJXofu5VfJEQeUxp+DQ172/rwrByRM
1+Xu+7x/Ons2Y8so7eQ61iWaobWMjSoo2SsDZC+k6xpeDD5ZHVY9nPuvK+CiWgHP3/UUbjkV9TOq
IcSbAczM9biDeQK1HjHdhWYPyUBRZoNpdDoE4XkVWxTW6MtbVRpA8S/wfGNQCt3Izyme5qqxVJds
l9a4rUhu820M2RYc64LHX68a4KOsr17vxDyEPA8KEjTgje7PamBgTODF54XLzahZYXfekqnDSgLW
zF0GaIjqOMe3CBXI4sUf0XTBeC/LvnUJxZxIf5Yb7DFobSU6OcJie17+l8A5kzl+RBqQAl8KkHh4
1pAjCVHXYOvwXqT+T+IzYrQF2F+JQekfx8P1MEzcsdonkKg9PEz6qeJUglsTPDchBrcvxjVuSKXK
8T55Z2fliPZHPqxMrhR2h9kuKWACE5/RFJNURgZGcBpSkaRL0pU7ALrKT5mPXozUTAAjfNsuurkE
hokJPpr3NuRDmFxK5rTOyGMSYfDTAcB1pxvS/fLQ0ip/7vjwYRzySS4hEXae4AAP9dE6tE1zV2Q8
y3+qZ3lYb7yjk3P28+6FYlb5EgZlADA2d9T39pS1fiPWFBbgAgRwlNy50DAMuFrVcoV/gqYoGz91
ng3KvEMQKKhhJNX1ZQgyncmjSCNKQYI3c447CzFldlaH4bCVu5NFoID0VMoPFmqiEDBYvYjHJF4w
40C/i/D/4fgdbCWXQ5z91Eqqq7MWSlA7eUXJ5sWQKfntLGAf/EzVLxXt0Ti0xSlBa9k7M+SBhzrx
EzeMmRPM4Z6pdgG4GRBu4R1S0wIPW7c+hPvkM4XjGRMtcYaUDZrCfivdZLp5XIi6o0NfPvzzN4q4
Y1FdEZKpTyEDVbmv3Jdc6K+yJeVe+k651CsZtS+ZO8iEOJ1Gs3R9D8f8wAoxK7YYC+Oxsvjk5AhG
m6qDMppylLu7EqBT1e4DgNkVu0aktv+F+ounoUHcFz8gGpV9kU+Q2FVQeOzP+5yyeeMjQT9lWx3X
WdGbCuQ9An6y6ofcXjPUnn3F4zyIedSaUifFmy93C7qEgdSKgPjbToJITtewCa71xj1xuwGmiDeN
YYhUpxIbAvr1s7zjgBDFYEj0g0p3/rX+mjnnaZz9+DmTjbvXxngpsXibBLOG6L9/HjKJcKCHicVM
xRu8A34SXcTZAR213uqGd8md933kV+vyWdoSwjCIP3z0sN+N0CkDgONn/gIfFIIPIGeQa4FNt/v5
gqE8z5FU3anfZvALOrcw2F+q9uMqVwelHm6NjlBvusg7iH7hAByiwNkTLI5tRY2Zm4+FajMrymMv
DX62zhPvME9vgnAQ0BXXX0aHg6XXTUUk528yEnjyUoWzb64VteMbsWBCtBLT4A8M9mTKUaf2xcN1
BLtsYxgSkX5A8iQRlsfkitIZ72McptvducLaeyibSVm426JDjt80EmVZvfwVWQCkWwbj8MnGboOf
3gZwrvja+KMpr5Q3Z4kA0mwdLCcRAtNkWtgKXfbFq5P7i8PzxzZJf0nsZ2++x9LDfl4PeO5R//EQ
ipK2T+g8Rl3KtNQxWA2uAj7OTw3MowpGKzzzcXq7hF5uhdmMy/q/8ftGJ1W4AiASal65L5uJgErn
KsRPmmoUAnn72AnKnE/muMrrLowuYEKpE9Egt1a657Qcwti8E/rPbUquzuDLBN8LEuwvMBSfciXv
dA9NXw3N+lcqvtGUZhWD4+sWdUezH583EvhLncKMEWyobyzDGK2XDz2KCYH+3e8m/N9h8E79RFed
kfGi63XBLK4gFyIy+DAez3hS1kX3gY7U2VoVokRVWIM+V/r/bOq17azb2qWelsD9+8zU/KvZfHoM
Pdg191r3G6jbcW/exvX3lhJHl4CktaSLA4MZ9k2nAFVN4A17ebOlMp32T00+w644PGOJYhHxrTvP
gKxdl2jKhV1RXrm9OBL9iNSgrWKpHnPFnpCl0DNTeSbJpYj8+2r4N2t8gyxJ5MBzvGa0chszPPea
Uvprm6RRXbP/iaqEyiNIJpjAsaE6oAMQOgpuu16YPBQWzvAECEib8rHMrVr2nJWIZVAUIJGOGIw+
IQ/LE0RWTdABrLsVeAQ/Nq/lRW8dMqyxHWI8gfN9NvZGztyEpy4rmQhrDSDKIJ4WoxmwqsPwnXci
d0I0sgC8mjuWZfaFJepjhIFeFcZTvAehup0bmn6naWTKuVhwD8S/DsQZDo1rvNB3wsq4CyQgW+Di
IZwnKx9fhCfAq2ajgeor5tylzNkWPYeDwZy7UJ00wvRLwczvVp/8J8k32DicfRhmR/bCgxyC08ks
arU1dpGI1G6/Xvh2DM3AGEMWL5/z0WjT5VZx+5lcTqECXixm9/haXB3a4XIR9rZZcat+zGNrg23v
09bwEKf4+q7yU6mj71rTGIsEAIt+ZywLhbW3D2MKbMky1creUN2dYDCW0vaHVT9D2vA4h5D2tQAG
D4o2BQ+qyXXqKwgIJeA9a+L15tfZSxfnOa3wAtX6LmBf4lKC0XQ36c3GPNhRgh3CertUrUoZA/q6
33R7Y3VEwOoNVFglTWOk27lj2BjoGvOoeJUpdn6iaP0TELzAl4LntJbFYsSZbeiKAuajS53MXtpA
qfMJkUcwODrQIJKUa3+pb7IZD+jO50+0iuSActIH+q0NtRD6RgxbfQ8WYa59jM91Y9xOk3dK1qzx
LF4zmPxDiu0f+c7Vm1Fv8kdD0O0Z9d5RaWUXutVdWxzTdQ10kg4xVWs2MvQvThdDPrYraOBY4Jue
5p5U99vE961Pvgyv+2YKDyzk9GvCpnqqxY5ifrrxkYVtoI88WRuIQybXTEhT2eD55AAMMFVeZY+v
iyRydONSvUTq4eI3mQ8OJZUI7EqXABuxt2iJdqjP3Ea0d9UvbYPam1gwaI9s5xT1RmtUJd8aAea/
ks2kBTCax55+m3R3uDqvSDnWC5FOKuZzr/29jw/kAL9s/Pum4aPeTtZhGP21L+4QUnC69S3UzHXl
vjKRMIasKxZFugSWE4eVOdQFOvRRlqgVu2Z1fCe0DPrxc/lbsYv6WF9kKtGHMfB9sAr43ZN7Tj6Q
D26D7rn0w7m4kG8zr71tasYlLDcyn4WDqUBsRoTc2Hl4j6vtEtJbHXBg+oXDCK2u0R5osrtifJjK
F2MRBtt0oQ3IHhpPmmy3LBoNXF+x9IaQGGwJsTb879wxX7AJolySe7oS5MJwFDRZt3oXxsTp7C4n
cpFaDZG3HJQ0lmW7PnBetZYiKVqYjpLa9huKK6fAHIO3g96ByForQjO0LbeoNFFPGPTXgfxolg7g
H58njvUjsQfvZ3ClwuFiHAp7rA6jEzgbICPFNLvQwCfUz5G98TxdU6UvUbXH5xMca5ZFCalXZ0wy
B7SeAxVt2IkZNI+o4CBWyUaRKnFDWe5QSn95GyVNIRXjIsm/mKNE29+Nehul8T790FKFQrmfc4nt
RAxsHp5/BWtypuRgLrQXV5OM719Y16l5cPcTDaTQiA3aibT1rQh2moxhrAenZNQZfvSaRXFPQTs1
XsEV4/N6YYVjgDeWQwf6Vuy1N+DzsmuGLPTKKP6cn+7j4cqOtT5S1SnqjpOpC8uz1ZcVw+aulMPl
12403aQr4L/DlgNjLvq03u1tIDKOXr1CUIRy8Bsu6r7208DfAXnebsTmopjuGcFsS3k9hcp05fLq
VV/cdFMNxnv9Iqv8+tMYRf8IS5xQ3CN6bqSY7WvoLNSo13rasO1026dnUW6jAW3vHDBMlnCiLluZ
bZ52vc2Mgp8ZuVWhuaWjI6ZP2qY831zbobj152bFV3Kp+Z3oZDN1cPc1VVlsPGsa0h4GXEqeSIMO
mtaRl10KS8hllvt346uTpvDphvcAd8mrH9uehD7bOZcUY2TxCmMl4fdXHy0atyF+RqSqPUzWhH5M
Sp4KVCoMB8dQPGBB1rT2QnskLuRUpgl5UzRdfd57mrrfhcxlzaC3q5Oxz4TmpGxMDdDFrycrYlPj
fWkJ4Mc89islIq1CzkGcjG/AYfHE4LBHsAtTrUuBKv2TRuschmyWmFDc3Ka92lMJjQpcAyNWX3t8
jOtwNo53QcCmrnZYK3/0AokA9ZnP6Wp8dI4PVt+uMTEqanjscqEsztlXwbHCZe6i04ofOWmWh/Ed
TRcOxfx+IdcTyQFZTpsN1/ezxiD9WxpYF1Ge0C5qIn2ukQf7+mViaZd2d9SewAm6wXzaC/LJkazo
bqWlIP8L4mmj50UTXBzv0s954FrxYwKogpaxaNBJIvt/kBs9h42HPalNIo5KpMrq4mEyTcFUmnkg
J6CYR6dMRi/Li5RK5oT/LEngF8ysvOt/Ic2RV/HYJQKpDnnLBrDcpt0Cgrqy896+Xd8QBSfLPUK2
zxib/tz5gauwLKlBCQEgunhuFrs10wSW26gA6/nRCejTgyrcgyjyfLPmo3Slf2T0kjHt9uGw8jMJ
gZ9o62qPQ0vda/uvyneAizuEaS5kSRmiapb0NiP8wXdR8pkarSMv6bp2flRbAKf+m19dSWxXMKT8
R2IF2T9BeN1qvyqZ7tKgF9xZ4T1lYq8RD9XCJGjWU4pF19FPFBEGa5RBIhc/lDIO/x1f3wZ8nQZh
5Y0e0vfmWWrCw08bpmXBZDJtBhePjZq47TUrNGzyvSrp45BWNH22oyJXNqPio/lJ/PtEud7z2qvg
jh/MbxY5FAdDSBAFA0eIAimxP9Q+vCupFzGFIcq8IFLY26QBbeTOlxMUDNuulEgp2lT1w4c8mxs3
uZb5uC1QjyRhvMqfv2K6e6/Kamoajc2dco9YI1g2kVn5Dd9EPJyh3boIs8sCJiWU/w6p87JG2hnZ
DLwy17MyhJxP5APg5CIcUNg/TRKjSLye9ammtoz88Tj2321r3bxagXjAtHNZsvfICN54xHsi1xjM
hY2eIR1kzkx7qqu/yNPjQfvyJWMlLv75PDYFvzhiWoABUyVBhWYHewKvOBYkJHJZwuO7XTI9jO5/
63inEPkgzijMKPc/tFQapqZAvUeb/U2gfkO6SWYWfoYCsxFQJxh+rP/FnLdQZn2O8TZBVn/uR+Cw
0O7W5iTUPYbw4agNjhEXbBNXxL7htMT7HfFIC1JnUiIDhFNGizq2ntomE+AQKd6Hoto3zpfaDPcn
v9K6fbJyQrmBvL7oHl1lvJWdVAJCiKdJ75MGY9D/n9QWlG5+HzVX6H8yVGMOTNfnKGu6qHKu1Ia/
tsB0n1TCMCxaUZaeqiXwtDeIXE/jH5LTFMoDUm9uaWqmfjcCon6hYx7WLnnJwLdn/kIz3/YcyhPm
hAYEe2T2XsKQtFwjjKPwT2fdOm7rr5S7Rx0/RA3w8ojgbloiqRhuX+/ZnYnj3tpY9H56jeH7pZt9
iLadaCp6qpNcbOnQaWWiutF6qSYRD8UK5ZFqYSz9DD9FP6FvdQBRVT9bwa1jwlSv2MI9HLCQpK9b
E3wFMu+9OC1eXHgNusQ0RcktG7lxg+uM6ZfyjtQUOakV5Msmsuhj3BVONqlg2n4uQ/boCkJuSNNB
Y6k5vltqtXGtN8/Nm4HumBI4mxc/KOjJictC24IQagTLRBhJQV5idaFD8TNWwzL0rfQwt/nEEPiT
LG7FN6iv1x4N+9wybSIp/Q8QcEaCvXCZ6qx5gfGMvrGTptUpTvrzuFvE8ALBbM2x0i5l96wEcb27
maQlZMK1+GHkyXeLFf9KG+fokhiwRQmK0vBZMNV9FVM27j/N+j3oVXnog9uHeIdlCHCmYZFazpPW
dRV2NTOrk04hlifyca0z848jP0NsJhnzGOHWDXRovMSkp8a7Ttc982IrEKUGl291aFAcBW9C66zq
UbMafIHriaejp8YHxL2Ho/VpWSXr6bFtPtdBlg1ewdkl/PsjGvpAQykY4othXbhgohwhrfgzfMVp
9g5tZ/3axPdsWCfOtX/vxNK8GWAKQJEhFYMj5BuUqfRCuttDvKCRTKYfNKyXdi8P2QirNJzlEE3v
Y+g0NlBhMowDJBdmRKOILPMWOEw/ecBpf9nTy8Ju8QB1elBmgwunp0ycR7yn8edcimB+Qei/uWHp
XZe8O14W/J4B3FiaWYG0jeL8ivq/IPnxdHm5cT1Q41s9zgXojxm4t4YQVltYL32in+h7eYagFreV
wHMmYqzf9kpF0Lf7jbzBcxDuRY7tVY4T3QXvuoGLiisNs/+b2cJecg6nnuaWavLqVIfXITi54Bps
fMz9ftg7b5vvjlB/dGSbNC9G3x8xswvmcCgLAHqfMubglDJ4UurZEnD/TFQWTG/uSQYGQoVJbU3o
W+LwctIAj1i6jtlSK8e+S6MTWHcruz46jpU2IEj+V10U2kZSZPDtyhwi//wL1qXW9/TVxK00SUAu
3NqugbW7Y23Ss+qu14DSWY38asM0g/EI6+PsJ2lKqEVGJwo1vdGoFehE59SfMSZNrfze4/tb6k1m
KhiQKAvjR/6waUd9wU4BHCJto8rFTHZqXWLYlVzlhYY+iWaQl9WOvDz2eRwkdQ956WTVR5TXzuAZ
SDgZeto8CY3oqWV7g0ieDWrLzfIDtsxWy5Su7tza8ohfPqYzDVQglG7bHo1YKD3mIfW7LjETjTh4
H7AuKOWrgCoh37C/YhwcjYg92InnmAQ0tO0qoeYyvLjG3O3z1lunvdgxmmH5WeFIsnSslbBgINSi
sDxR0v9YQbiEkVNiygGLfb6B1vxY7PDPJ1DljPdgh/kB0Z6Rcb+xCwAQ9rg/h8xt+l109hF6L2zl
CvMttPfAdHuQkmzMUnTmtjoS4Ln1Hculqe99zNs9vVkP1div+3kYaOLf53v89WEFepkYCpWGCFV9
Ye3d8bBve4wQobtePHJ4f57PjnfUKYAjj/DmkI1jkdn+KrQpDAzTwImstp6dBvGb4cso7DAEEuVi
XPQzGLS1vdAhp/CrkGwl12QhShuot9mgXRr9D72bHzJBy9XjoklS+hP+N1/Kj+KCNXG8RVQ2khlD
DahosrCcf1dqQWx+vXdUItlXvL/ctU7Somq3Lu4PItJdukZt181AOllY5ELtV0accfOHWjHGYu1m
xzqr4gQdP4XYlQRPYXQCJgXcHLy47tZuoy1Fght0vf5BXYMlCIvO+Ydd+OXNHTZvIfen8jhtFCsJ
GziPp5BiQs1rVd1cdOwVnTByVZSlyvHJgWEXeR5nko91ZKZtLmZtnRBzSl3mvA8Hc1PXmtrvMlKk
HMzRvs6CTUuztt/GiQhbSgkYIv7KUXhYzQhDiaP7a/WBBTk5+zhvxlcEV64RTCqPN4u2z7iWLQMQ
wIIyqhSkolYpDRZOw/WNa+A8udm44gs47kvKKCFplM7557+OY5Zechs3kfBDJF7yXg6TLzHNz173
bJ3U6G08ctIRpEfIRReyHNL/2PJChE2T1gc6REFesKHV6W3x+s+7lZ91QqV4MGeEoQEkakWC2BjL
Wy6/Z9mH3i684nASAAMrBDCJ3ej+SciNNkC2WV0EiS2QFANVqRLwRdGQfD0+pP3Fk9SeABUJQ/t5
pkFVQsu51TegqWLy4JLm/BqJ/vN/3qCTt/Q9/Homh/l/RAKyYYXkZVkPcQitV3Hc4SnwK6bsrKUN
c//r9GMbm/Y+ZL6XQoFes6GqO0egcfh0DvSVPLc2Xk6bzFNwxp2rlCba1vV++ATh2p4yAZeaDtSR
bj+GYmg7UX2nMfChj/bb4k35F6w48Pl3FFZy5w3LHZ9sXsIGURJrKqj4g/v/W5GiMMcvN3gb5RHp
Gvgw+ma+B8LajlOi1hoJ+AYj5Sd81B7erI3DbX+2lHmh91Cpzo2ZEhJK1jlOYUZaTBZsArDZoVSD
vesBVF+nbzkpoZ91lnCPYnt2jDlzMiDaXHtU3H9mt60Xi92ll0Y/CuDcrB3x6fifKowjvbiCe8EU
+9n5kF6V1fWzRO9mlUe3Dk1SOO2/Xu79ETbBqz6aV7DULTIr2ZX8ZYpJhY6ART9vUE2UduKp9c29
P7wtNkIvoxePh53iISJDCiaZIIscMjL1ApVd7jqW2g9VCwvgBFNgEiBj43+DTDrwG7CwJy08sf3/
Yp1EsPkH95VQ5KO9TifulZOo1Cg/PjjDnuEo+iA3AuPt7iwLqtAipsMMIGzV3KmznYPgpwSHTdlL
MzNaV8poKF2vGcPnANLweDT+xnI9E8dmxt12UyftOp/IbP8hN6NyhAC3kXAYrg60v4A/lA2/pflG
eVIx26+f5dAVbvDqESMmQ6X209cQtKie9V3CeG3XRHQpXHa04KnurAmVm7TlEvm39OfGPEL/DUQC
ivAMI/jQcU6/we8PGvbWn7FXEujG01M32gnlWzhu87A0NmG/xBb58XNVXBYSc778kDy5LnKNYkZy
ZFAX2YVKuE2/FLrZUi7goCmo+uEaemyApuARSL0RervyM6wjk146hjfOj/WGnU9UYuilFOwj0l5t
6uwfzNLBtQG/sGJ6tcjQYDlNwLUa2h8nMEoVo7zotFnVZDgANwHx+vlsj8Po616eqCz1TbAR0D7z
FiPBR1J8lLotl7ZlBVo4wxHOr9JgkYTzly4o59WeJ83C4M/ss/GuC+hihmN5TrgANlvpkhTMbvxH
yxsDXGOLLvcR3h4dTbO/aQInNfiYSe8RLFY26V1XOPLk7OhGuy2aoh+ZOkdEI4fSLqXcLGb8eYPE
po/k/4F4jMImxWTvpc00kJMaqGE5lC7vJqe4fu+WYTnvj9VfBvH6m/TlO+wWQtcL6ueGZPKHaAN4
n+r5MdiZ6hwpnavVwzOmT31T2E5CY7Srt1JFZl/GWS0I646sQNQvDX2hHBfsN2+piYTQmLWHESss
Et0DA42SFvK9iYulHsMXL0StwZGrwY+bgT0bV6oLVOwgZBlKUVr/GmR4eYl3e7ECOb/94ousa0zb
FhnOExKO3FUeOSvHRbmmLef529nEF2mcRpJoeAIg6Tkgx+3HzRRV7SZpuqW/LwZPNDCdhVfRQOE+
kHggypGCuWfJ6DfUVjDBMwZCUgBwBjN3cvaKMSQ3ly2ROp0S7fs3bxzyaxohiH1VQpllqIWQdD7O
AAfivCs1ZEU23BH9MTYV4j3YbpqqO4GqnLGbloImbUTtKY8wPjp34eLxf5ew5IFuHL897E1SUDxE
q3eBgr747GZ4PR5Pe1OeMe1MzfswK9ni/QtTpw1UjZlvZWPkCKO2e+IMFo4gURgoSYHPPXrpvw2X
8xEf+35QyfJBxusEa/RMfM8+tklcBPsfNjxtFfPK8s3fCAtrjTRqngPT12/BOyLNzxAcaJ9mtkL1
IioTnWIDbbq9vjY317r9PCiPRqx0Eof1VYTgGicWzf/ZGD3DAVcVh8gC8wblg1zK9ELiF+JJ6md/
9B5zgMIvJw82vQ/j1P91MJBeBCOMHqfpX0M4mutCKTbK3E62VrJHB3S7t2NJ7PIfPkC/6VHm2Xfq
f0NH7NUW4YfsoCQrb20FmZwKwvTLymECSWjxID9WeTPi2/MKtZ4Y204Gb8HDuoTpAvzGt9cUWQS7
gAkHulpTydwngy9sOX7r1RCSNkbQLVYAEvXbdX8D3ZFf3HH6KpKwswimKYK7oTnvHydBup3ek8VJ
adDePLVWNTh62emb6GWTIpLCItsKWfHV75Hb8i9rOAdLD3vdhaju8vJGueWQ8m7tteQE2EsHffV6
wVR9XojTE9ey84oVqoaa6HP3o50JmgAIYNe5PPBkNHsOaflPDWOggo4iA6mB5TR4RNN5h+szMqOO
1RYR80+MOUF4dgvOh+u0EGWFEBbgNpAv3w2QIJborYYpnHUlZC78WjKMZLkKNfz2TXYgLkaxkDgl
0Iam01E+dIspxCo1U0cYFIIVnAXzMVecy2I/NjYnHBXu3W3NuIjJpt3UdQInLxsbtxJ7WRslCoF2
wE1HlBxxy80xpBv490t0airoWn7ADcWqa9K1TEo7j2huenm/85RqaxMjfDfxt5qi2OxdGTIk2vvc
EzV67UdUPl1L4/FH2/EZsYcBvaB+v/KxXZgeTUmsTFwW648BK0wjJABeUX82txiJAm8lbzFrcGu6
S/vtQJiS5iTP/HaXG6Si0lPWJzrT6qQeHdNQZsRfYfLbek+2QC0Dxt9ONqeW2M2L28W+9oWhoRl3
of5/JF8/I81eX6KnpFV7pFqYAIO1A3BFWt1PSGSMzSad3dIFc7XXYykx8FVsJNx2E+9Nv6kxv9fo
yx21xlZNwRHVgvprTvwhsurydtDFDt/ye+tJsrE2KGDns47sZJxxqo7zsY/dwsYftMchfqVMzctc
pQ7sInxk/1G87IWTFy3UK0dOVIradNrnb1kH0a0dHl+XxJnVF2GphuRSzuBUDsgDJIp2g2HtVIuO
3l5BetlsHFcVy9mFHO3CWnHu0aJD54f+pKY32ZzV+slxGGVA5GZfm/PXW7GOLPQjsWUST4qs9UZf
8W0KtzpTA7ieO9rx0mSovIGEZmRlgCZPKAsWhhg1LkhjgDHtN3BDka0U8z2WOssGuFl9jT9Agggd
jrzf2Qsdj3XYHv218B+ytfRirVryZYy1YyPzgCz4if9qvtWmkifeEXytREHv4B0JmNqNmsqU0wJt
WGTWfNGiRJmZMRni8pQ6R9f+XTti5gEEPq7Vik00zvaqbGcxuAx+0scFKhRbwbBy1MC5KcDB/GSL
Ktg0I8smC7wnM0k4fbWSvoYoV7yFTBj0V57rkbfVYz9ZHb5YV1qw8zQv+xfUxo5JZA83DL9yLcdN
/99EvKJLk/+/DEXVBtE8GCC5dLf3h7fr1Mdm7IBz7Y7iOGb9w1yeYhMRxo4Dgx6gfL4Ra3/xA6Fc
tKRvWmtZT9k97Wc/eED04KkbkUwGm2g2NSvVRPvLsJCS35kEqaOxbGRaqBfD87NFGiWkqJ3SXu6U
GWrGZcD5n3hEUoCxhA/ljKavl+PTikURW9G0zGk4T1Kej92KHoRFKNiSiFsafB8dYvzUQ5B2OBkt
aixDlukQt98sX6P8/nNoraFwH8ho1ht/JArxdnejx/K/LdWYDgHZwlMRs1nU4T+GTFOcwwYIsGfC
gyXaOTL6Zfm9vNfoOADpmn0sUJHHa0XKQLzE2kcRXK6Sq9iaRg61TEFbn0pK2S6wKGGo0G8V++lM
fpk/wX8TCOgrh7tDoW8OhD1MJ3TmdWAZyAyg8QWF3L7Gyh6Pa6b+XlN7QDKcHetxGfLbM3ZhPNWW
sdMtiM5Svv3ILHQxtJRdWGs2Hd2y2PbWaVcE0jIr5v+Ma+3Hc4D1bLgXJrv1SFPIXrHSm8DW5w/w
Js19irkmQfO1VikMNZBEN5JlWKCLfceWsMnL6+/DsLCnG6vpD1s5HZrH6kxhk3tkkQghsRAUr98z
PyqShWK2wVj1S8L+wX+pxAzb8N0BZ21XRURsvTEDNRqYrETV9gPIV3om9zfMl2PKIWoD6sM+4/Qq
7UdTsNMAvZ8QZIzLDheNHTX/DIIcpSJjNCF6JNM0PqauIly9HsSoKfXxGKr7O5znHQAGGQDXhXjY
qomwMLYBOK1HGR0eeS/utaXTC8NBh8siJ8fxm+4+iR/VTG0TSWGNqxLuhM8PFAjcDrXaseM4otcS
LImVwQNkkV+IrGGBfLhs7R9BzTmeALopzc17qWPnQtF184rlPAneP90uiDfAdAdQWHuUtQSBdezW
esQWcJgNAJcTS99/Y6JIiKDN6WC0dSPeMiSWI4xAkpJFX2NFb1KHKXpGt9nsCUZjTmKYz5xxWL83
jWxqMufzuQuv82Qr4eh70ozAILPtO5jNT8UypzgC2SctnBx9jqadhaXtZqq/IlfyQspyoJ9/iz09
2bahB8+pGYvWD2qhQUpB2L8gCMbaiFjS+7xzl+WBWP7vSfHy2GZaxE8XhQxS0eck98xX08UmAVZ4
7DiyPDck59uoT5A2nXq81gmfMaG1P+e8+sgRWVlm5c7YjNPS7DpuYP4Bb/5mhVvHjOw6syTLObDj
6hxt3LUAqyJyOQxTHtYNcbGAMfn/DJe27A8EB5Ejjgsjc9oGEIqxM3N2MKZlohJDGP+Co2zfTLTG
YptOlkMjTjS71j021DsAGwGntomiHyDhDZmJ+lLEMxPvJTMCP9oTjHwmhHDCAFcnL232CMxbsA6O
ppsSJFkuTdBid/hDNFS3cy2IKCRUw+ZblzjVgx+Jv/gXjjO9/RlPCfNJ5/pN6hZLom4xI4RHJRt5
A2+uyQc6jwIDfkhDn85A63RGxRsyJMqtTcpTZK6IGqeb0JBnZgEyJgswKUzdktdyseH1SWOHIG8j
ykg8wZrAA+DGqe8Sqn8BGqN9E2rNF36fqve40EhGQSDVZ92+LGIYornKg+plfvWP5HSXQ10TZxzE
ZiZQBjYdxf6Onb/eI7bq2y7pk+YFjdbqElmd4Cz2IEf88rXsm8TsE2gHWEGvSQCqCwy81xS8pEwe
OjRYp2rbqpbH6KBiIwgubjshUQ4ZBKrYsLJzDBOjHCN3wMlnsTE4kx4/4n5k8vKOVWY2P1RKIHHN
yGWd+yCZxH/GHoVkJM3ZQv/qMw9vdYV6KbR3f+5RWrRIa3n4IdPd+ZsbBzjkxrdqqcrVpwjXyslf
Cb7Do/jXzADVfB6+P9JjM9BFNcDsrVuwZD52VJp4BQIeq59kMTxqqETXepf2/f2+t7mYGEmCf8DA
kwhn7NqwN9/i6ANgeuFqx5BDeW6tpjyJMcyoZ6JzAxIyHNn2/6u4Awz/n5r1BaYkJFplSbSNzm+i
JtaRmWJqRsFRcC6QcOWito1+lqFDz9iSu13qEYYONKpxNn2rbMF2ZCil6FWwDbBYIibu+gizJLKH
SWH/JfjL5u/cyU1gRmqVFhd5CWzqtX9oQndAPGGtunSwB+aojPQcnrxVvl4dR23+NgMAbL1uews8
7wHfdG2uGWsletXTp9uOK42AgdjkqAz/1U57t3LaWNp4lrRggRE7od5fRzeczLpnOBFDbOr2k1wK
DSiRtvdeha9JQUeSlIb2knfShnTNgOhgQFV2Hk4VjKyCdlreL8PG17unYK7489KA7DHnfyZ2+63V
cmS5XAaUwRFU66QCwcNfzw5gkpBUi4Yfzy4hLmCi8QzVDVOTC6wrAah1dIW8snGWrp3DFBb/JMAz
RHuUO1/90b44Cx828M3VQgaJD8lZ7dnqV7v4S5KqRmG9GyL0J369V8dRNVri1OQsBFGgMgdbD+kM
3js9cELKcLHq1jkINBSESUg1/dHeCbIOEybPBxJ+6bl8zJVH3mc/dS51IPdZpK15gtAoo43VfZNq
+YeZ18X7Zc5fyZlDiCW2LvjSV2xb8qXMSVnm/eW8gK7vCtY4PWVNAJQM7veJYvbrC9l4ZoUTl4X5
QaDf5Hz+cDXhJ+/mUH+2H0HHcHurU+4l9yB9ME8tUhzffovwNQPGp4anx5rn/BNhVEURcbNl5aEC
cUZYgGS529MC/fjlo2khqg0/RaKqecW8YPOqodqjcBFSaC0g2PFe3ySAR/Om02gjm2vuC3QEsqUL
HjsGc/80DHz1zdo2pVYh8RlOvqdZA3wyZqLNOuIGi7+HfJNEDeFBy0xNJGsh9D2KV6LZYHdCBE/5
Dc2gb74bQ9wzF27KG+yprmy/z2V2dKPNY0m6UxLL+PyFDWHu29JgvANJSs63WnP3d1j9yoSrTGEl
rI4b0W4nhzVzFlsbBoFY04TG1foOszcUhEU5zB18NJbkJpmjnXrnu97qrqiERFW9gnPSmQHZBvu+
D0JQEwWmFGO+pv0SNLabcgNuE2LYRfkFXWmErXoC6DDHeNiVCybSLkd7DUhiQWYKYkfubhnJU3CQ
oPKVKvgO/AgmTtsiNwFeFnI4bfQvLjSvTO2ANFqWEkpqV2oRW0NSVrbQZ+DeB8xrKz6TOtXwD7BR
CotqCOI3ii4nIO6tsDUDoVk7lavid4CGZ+Cj6YTpGI6pKIZLTXaJ+gLYPTmxm+cKx5+d/yQ+Wj2f
RV2WD0gP5nc61exwbHV7Rj2F+J6zyKZGeSPyf+MAXo/KTgm5WXyjwNZWhhEYuNCPK8u7w+MsOkbl
JBiIGDAddex/dWXiIzSDTkvBT4cWDRWop4XJkf4Q/sJqK7QgiDYQGjxLePW/snRq4mgfxe2RRdHj
+zRTn6ZGCLB7RLNkJqrHKjMMVUuuB8GmbXbw7vQEvD7O67yG5k/+juPfNfswRG28jcPPCshcpXts
G4pqjVFMaCbltcuj3vRMDCkkAkp2d5kOurBCLUD5yzYBXxCqBmeCKmClvIQKZTDs9dcpIiBt2dPC
GuVK+NYC8v/6R61Bwd1P992VgVvETwPx6+dSxmXw5EHv3XlqIvdf3+1QExZww9UopII9ZEHcKJy1
bCHO86HUeAZ5e6QkFxl/ROF0n+sa4OfwlQXIqYuA+DzhiSJLK6/H2QUdqIUyW/1p5jE0ZCniu77J
KxnITNlpD8RBxZw1WjkUeAyuIALSlywWNkPDxse/H6tikoV4VOJU8EiotQtdGe6BuGmfCJNMnq0Z
V5r5eLrKXENmhjHnmyMxEdNK7zsBGEbiVPc+tqQAkBkAS1z8/L81db3RQzq4gfxcUUGaxtU2vojT
9yVyVPXuf6lgt8+pWST7QtzyOTYcAWmIOA8fIChnqkl4plbJIpY871TvE1KQvEXZbnOvJpOVnsPK
tcsJDPEiOlssSsJXRGXuBDSKzTh8wPm5esiq2zxcC0pi2gNCo08Pfg5TCuFvOdLXAL5QtSapwtt0
w/ylkPSnZISJ//ivBkew9k3zYWJ11IhQZykVouY6dsVRW75vTgVrWheYNLvzNxx62SjzJQZAwPHE
Sc9QcLtkIqh7FXQl4oG9JPVnHcZMZ6xhnXIH04KGWdeRt3xtkD3q40O+ju0P6yLeMbZPl6Ewztsy
4wM6W0Ii+MXnH6Myj3KIheenfICmO0VIqQXRXfRWE3RWfM/eTIiLzHfSHkDnaynhsQVkmctX+hk2
RTHLpLVQUb8TZ5TULQDX3LrgmMc0O3fYNcYxplGmXk8mNwxkQLslVpHufUbWRmQ2DRNJ7ZXabtxl
1Yj+8NC7YONkg7Qz/2NqTX0ABNFij+ZXnnNZn5unfOKTqNehOp29s2iEJErIMfwOvvzjo7SkHFWm
g9ZXdGe3EYKfRiLkKTLzTkASSnE//UcNAG1iOI2AmdS+FwrVo9d1lKhIyxozbw023/AmfQifQuG2
PySLp2ZjSc+DnGzxsHaF/VDPhphgs+FksXQ94ZIW4/1Z6bGrgQzR1z6aYsmPo5+ZX04q18idFk7r
8Hum7KnirPgSAsmQ3V2qBj4txIx6sFrT/VKDAHIMc38ebjYKzPch3rEHHENd1fzreq4IjNxrteRQ
vUnPjmUJbEHpNq1FYixE3z3fIuyNPdVdT0WYgSTjoLQYHny+6nynewrIx6u5eJ7NwuAtszcXuDI9
AZuFbAi9o3Uoxpnmawi+Lkp7gBqPqkjhpl6oiyLzB1p4mMSUdv6+WAyvPz9G+NZE8hGS3T7dhWjU
VhD6ZvfLpOLhoGQaBScE05HFUWsSn8qZeBf78HHr7GJQNmBx1FOde2CgreDljOtS3MMgTfn0kcO7
zcVjqKiiYuIXrMxoNZHKf3vMHfmI3kLCdc7mKMMfLM03cyr9RAJ/wLpvd4eWSsGu9IK9e6R8OGr3
PVEKC6+x5cKpRbanjscNIc2YPyJCy0ct++M52Ap/AC2uq11rD/H9ZFZtBrZCR8qpSm3bUdeXTnFm
vXa5sebWl7/72LTCwXrqUyEkAFXjRt7m+u8V8okAlQl0mjQFbnBwkZCO+NYgpLSFrTb503Cra/6o
HEXiYqnC7q6jxg+FI64pgVpqzkE3kKLff9K/0EfrX0eZyHb+8ISxE7p6bGBhb0vd3bXuBZ30qtYP
+Byi26PSh45EcABAiG4TZvuEJvW6N7liB4HgyaE2Y63KD882qDSBvdE64QDh4WO7sqQUkC8GeqGm
9VMPyqtS/vkjxipPIhBlMecAQNFfhEMfgFnpseHfMzFBAUpVtXvN4xKIybOp2rrots6/+HpgoBmc
+A49A9kQJKGBjEB8Vjx/ccRucAxMvvujzWd4VhGKdx3MAMkLP+xkKuCy2/BkzJluM86g5Z6X+5R6
E6Q35MGfW0mYvVwLWSYI7mmDJbh57cwMk2aPyaI0oxQU2VSgLfBJwmY/pqyU5MVYM8QiUbzouoBE
wWLyQL/IELWXbVPxN26fCfV8GqHscY9fROMyaIJP8jmexWM1bWhyJhGI1YQPN535zXqaaSCI/HEB
bi+MfjJDVuzEl6r4mH8vCqzw3YDhJDIMRmrbp4vK1LLMU/iM/aokalronLKtzOt3pXBYyGhG/3W8
u1ufkCkoFg5zFaUA8JJHKjtv0SQPG+GalLOfSScpNblwaPIiZ1g/YSPHaZlzFQoRcQe/9rPuALgo
Nvhq6tIPKEXJMHJttT3Dy285OSX5kHowBqogkLr6hA1eZMUS38H11G47RDGW1s3WWW+B9eAKqgS5
gqQkFYon/8YadlHDOKECiPLg8O8s7YJ6FT1lST1fbDYSjExIv0s3zz0kiRJfVoUmqpKPadiIY6IJ
wpNMaxAc/1vkBanJiOc324fK3Wp71MtWb/OTjpY0zv+vpcYH3fjb0MWdNAvMtYUkTILcMlgihbIT
kcrUC9lpRHsS8umN3ciSFpCzDjesnVw8Lw2QLnlDyfeR47NDCdX9AmmnV+HevAaNCkDhrc7tCK2j
xjWncwMelR46eaBq5wpLlyD40st8PfVyeCAydYCZ+6JKPD3JVObNGlqOTW8gesVDX8HxpRnxg6au
bUmCrTdtgipzQB9P82HATWKTrqVzaPODPVRw2V51/SaUeSO1SFZQkFOq04bmZCCMCwaqaR1YIJWs
ixswNl6/MDuFZSyPmL5X+NcEsdV64YiH9kVEDP10wwmHtNMbw7g+FlGe9dYd48UzHpTbV9Q4W5Ne
fgR/VZ75M2xYvMj8ho/glTddB+3OoXaieclgQOrF4CFaPke0mv9mMqkWuriL2EE2uzPj6MPbHGHO
2Y7lIz2i0gcGhugdgtZ61CF0QJhacREKJf93huUabfpdbFSzUpgoRM26BPwf0BrJDps8zwHgd1Zc
buxhYT1+zQWpskW5t+O9CVWel6xWBtxN+IeGjaSMf/vpj/CocmG80jDDyy5YlyEM5rEKw3tqalL1
HwuhMU2cVXq2wfnnceif0bbqbksAYNyNDrHMLxAC0tneyqEvHYwp4iEDYq/3uYQVe0BkVuI9GmKW
6wzQnYVSTjX1180tLIUSfJmPDZFPft6FH4c0UO1dZ8sFTyS8rSqJMEl5KDl5sXAGM04GtY0ouEhg
zrlWDPX+nzr0FE9cPrKBq1tOy223Hm/vKRHlWiLKPl7oOtcmqub96tm8R3jy41dodKB8UiZ7mI/x
RPmefNBcSjr5xC8w/cfM7N7nmePF1ygIFeUh/YEOseX+dwSm2n1zUNb+GAKxHf68Ornd1XecSNDI
MSj2Dv6LWbPfzK5XgfnINm1BqVUu7ntch6e3E9zIIXaENq7E6EcT+7ivylojNPRRRTGMLJMz58VG
0ukrBnD2GO5+xjZWSSJZm1ACmuj+Wsd9IqHGXrQRC/BM8MWVWpn1d0IGhC7aT84wmTJqiNd7cwhO
4RQV4+tW8zSk1R8/619NXdxAbul5jnogrS35vPesXLqdpjeudRJzknoNWb5v/De8Cmr7upVz6DB6
qZ7n+6yCV6Dazavv1045bQtTdX8t9oH9+gXELizIADHMO59HsKAgRq4Y53Dzyn6+2eaIsbHC8Ime
AX/Bt5JcXAWsBwVSjm/pTB14sUx/8uSe1jtPNsK9xSAv2cTAH+kOsXl8Vq7zHjt9rqjlF16SUf53
n8pATYllPFzfeu0qzOOfMGtG5OnD2zqefoU7fYHrXGv6aUrz5o2uinun8JQ2W+nO4NWcH5efxC19
GkzDX62ZxoP/jjqNm3u9EQyGC4PbTdGcHFjx1TTT62CnHS5uqjsp5IhQ8ACE5Re2wE3rhUwT0a1E
TrXutqcTb2FDy8Vi7dEwIdcOZHQ2JD74nLYAE77lUWTxDgJRN/EV77eWKeW9+NnPHwGr4kXCKl0b
BbThX9O27+rX4pLh4ZFEkkY44/NCAuzLhznE/6Ia1Ani6U3ZSN5Gwobsa5yi2QDNDGxiNmGetpjQ
r7QxbWINBCgumH67F0Puy9bjPAPIamZB+BaL74tJCfZVxEuXz+m67VBsoR7oLqJLGspRcrLzFvq5
nIso0TzjUNPvuBB3vVCp2YsERT1/Doj4Qh4Bzuk4x+/bBOH7dNqCsQWlzdlpetY0GPox/XinfN8/
LRIPQFLN91rA4xfldXXDxth1PsGxiQWVz5ilxQvnH7yQ0h4hSbzNlEVB+UryjmRIRqXSf9aMphvS
6fC4drXPpDuGo23oxir18aY1xekNJ0FGS7+D/MGcWxYZPRHonws+SCyQI56zzv7RoJgiYH9UPsK8
Oc9e53A23oDnw5BguwfjRQcdrhXv0x5x3+YieTes3gtHw253YLLgXoEyB2r2xrAH4SEVBKqqMssZ
9vB0G/qPASab1wBzvhSbc2Sp7+pwLlx33pr+AE/jplfxPFS9IQ69og9VyEjtBx2gmu5CZ7Fm26Iw
90M+NmPBLvGFJhQPw9CFsB/Qbsj9drGc9rWN2jv6RaVh425YHWM4t/q/t5zIG8jt+STc3j3ps7aM
ntAIt59MzqjBEe5EdcNFFf/wdkwvTDMmlE1u12XN3/NqULmfCu4VV+gCDn2cKUWwguCf4Ve3Lr90
BFeCbn7OKw9WUFUS8jlKBFwbpyaMmOwXdFVbTkn5IgJhtkoja/4QAN+odZcQ6xB06wDuyYzN3ACO
PWR/m4+gLyn5Sxk1UpBV16ZPLTwVfM0ypyGmlRS3sRzjoi/EgI7KBLdSyRWGEaHoxU+D3/ZU9Ub9
UqmQxHQvV7JrChu1GRAC4WjC8krI30hGuQMRQ4jI4U8Ttf67WfXUBsHaZzHILTaLiaf5/vl2Pz5c
uKTBmluh/1kif1jdfbrayzdmumGIip9GIVaezhaLHlU2jInpmJhqgZgzHEXP01AYBsfuKbettKS6
jQHNuDdhtwQgnluN5iV6Oe6Wbh8LNx1to5PsRG1hGIFs9HCFT9UMTjEBl9Kq+9VZyezLpFXp985o
l2zqhkuuCcnh1+HQbe7WWM03bPXADEvPIyMs8fhhuZGBOfCqlrwSeS6hLiX4Tw6YuyHtE9lVsFAa
iXB+FbD0TZDoQgqAhTdYK/D5e3hEoFB7ioRoDE2uR1S2ymeaB+X/T/x+rhV9rucpf5TtpCGZbTsR
y1CigZRFN+ntjRSoE1Y6ntJgSvkz3gRVYIfJ5jQCLknQZX8XR5+DQ8XfVP4w5gRQXtLUvQh2t+Ux
Mv6p0tbM0iB/zpkDZTqPAboSmYnxOwu6361kuMEWedc8nEZvboHtU1TZI0cn8g3YM+p6hxXrm7j1
KhTQ66vLezNbmD0FRXQrNA0JxcTUkkxGx8PJ8nzjqRKb6PnpfCmP+S/8D8uGWe1WwkFLFc/wNnvA
KwFR7+hmgTHz883jDryTYCrm5FAX3JuO6ZNcQwb9X8GtzYr3U5i5102694yyQSmYYAQ1cN+IoKb5
+HGGeSUN0FcuDzGxJYYS5LK9J/Ukh1ojDAMP4lNdg1Sc9GIIv50U0GViyA77UXWX+omg8W+gA2Ij
oawvnSNiVJ8FWnYZgPSgAhJZsvMc9NELFedsEAQk4ZU4ZOapWiv1EenMWfr+KwJy/1jBFvWYlKDT
G5I3DVH2Cwm3e4YHn6T+sFh7Mxv5qQ0u3X2riWk9Iue0ZN+b9VsZ72uu+RN0GeT4jl7i6/jnHwT6
YAb5ietTwleE4nS2Vdw9c0xux2WuwqHNY8cWqba/BnYd9jhpMUF9X74PYftwfxaMFFoUF/nICbl9
XcSf0UPnQYtWr5I82cNFf/85DfG9aXzlJyyxPqalIz+8JJOx5sF+gjjgMFX2u6XnBHJ98DJBVNIU
tok5gDOOJJFEuQq/4JvtTcwKOFUu0bddBH+YwAAv/dMP0aHsaYWQ2428AT/XcHJDX1fkyplHnWIT
wPixX56O+UOFjAOPoaAni59SyB4iuOVr7aDhXx/2WsvtXq4kMibnCMtpWOXp7qbkfaIGQfNaGgVq
UhPNOrZh2lMxHjAUOQhR61JeKBnrNZr97aukeOexqVo+/gEXAmPBR0toPb6bqY4LneabxUDskeKo
CeDzeHfdeq2wteGkpjZ8FR35nJuVI3NCEKZCss/UQOAGz+IfRFYUhgnqFW3yTiSksHviqdDo7wDR
a25Zx6+VyuY2LHIjH3kq/AxRGRa9x1FrjGplAmQ+P7p48OyfCWW6nMt3F8wUrFs7lK5emvcy8YSz
c02uXfbQ31OmSZERrpoT03MJFGhgwxJP1oRwRBClg7tyuZKU8Az3XQuGOeNSRSyQn9AGVkPU+Jqg
oQCFqEo+UrwheUqx8WhZHJeKfaRia+bGt6lTdNFl9AGXN0bnm3sr1xYx+arp+9iiVmmiuFZgjZu3
/6YBkaPCfolMRyPhwmMVeZKql1+FkxnCyahoWtwTBSBInDQFh1sbrGX8YYtjNGlRtMKuoMbK1obH
1mTKUcmNUd6+8BGb/bFzKF98ISxUi0SAskUrpLSa6PIPuHM9cdG7WTvtpb0ZGBtvllbv/SdekOTg
CxGWvgRR1GAWMVjnx9FufR/cZaDrvrtPqX4fYjq0DqsetxU3TiwNZrE0ysaLoLQNhFiDnqlfnAFE
QxRsTwNNF9bsTG5U3mPylvySD4mT4EzcPdMgwxKudgg6f82230UojCctrP1In30WFplCcn3ypG4g
5h3a21jECBb9C1NbXwzM1+/Qy1wstCoTaplAI/PjUnCs0aOx22nwNsQMZ4STHxqQrUh78m2lOALh
xLSvokOfz9GMZ2bjKmAwC+ueBe7yqbWCqH3zFTR/TOHPxxVUCrM3yPIaTLxiUWJ2gBGiUbltWLIp
MEyvTQNd2Smme9y7JBvjFRdjO5YKs06U2qIb7pSyU7AA0blFX1xNh0vlPFz2x4SkesU/NZtx5l0U
GfexfUcnB0uOCEvlkha5hXtEXP6KLdR62G3JXKmBx0GTjRAd1oV1wRgK5FClOFnlx+ax1sSTSVNg
Zl4yqVOwWPQ9TlbLhw76EK3ScAAczhIteg7WVcha/rSPDDGIJxB/f3pswn0c7tPJwTq9z32jOelV
mdyriBY4zoFE+NatArY3ebR/tazO7ei1F3L0PDHl6huKRK7F8oNUlgh0QanWjosPiYoJKAPUnGZY
tkWNgMGFZDLsJ/KUvR6/SUljC6cOYHsiD1RtneMryOuRuACLPLhXugX0GPOhX3yV0XvZD2d1qYuQ
KqcqzpgFF6EQdmCr2JiAf9Ow5Uwyu6N2nvgsAtgGFIE3wovXky11MypzHCM+OyhzSPJqR/STWhWr
nxGeYnbow2LxR4BjFtQk7sNNpmFBh33R9+WE6fqVPYs2Gq22+cbSSjcXD7fpCK3aAPHzX5YM1xoD
49kOhCQfz23Lmax145tm9/8OmA8XDiuy+4valbOpI+gcBrdGXwXjZjcShV8211F+wG0b9BkdXizO
+aeDvIjgLWUFMzfYLBX9xezYhfPUvrkW87wlyqcaYrKnqTDV9a9cYVKQSyvk6OKZg2pk/qBx7Ivp
5Hc3KUCXdsw5icXjdWBcudBSVvf9bpvFqS3gQ591ClmOdM2mg2gNfnjytU8J3TBnaVi/qQPpJ2F1
+E1uQRvCiDCnW8lm3yOdBNFF4aLUDp8eqlJMAHILQ47ih1I+Wbe1ErSmjDwWKk9RguxM+h/onttG
b78sYg4XGuQvlPsCy8XP3Wj5kjFj/EsG1pnVGRocuZ6IwmRyMX4500GtJ8bBa+b82o4mLjvW0UG8
G45/yOE7h5Qv1ffiJTkd0/Bn0R6kdgKW61rCw/uiLA4O7jLbJD3BIG+r6tTg2Zdk+sTzHDxoZ/Yc
DE8WWlgKml+DyHIJgqv2EljdPBD40evN41pidf3XA+Gy1yyHNBvWD+yXRGH8rg+f/PArRXeYMaPB
KSs095MlIRmTKt9HQjORG66/MvMk2UITTQPFnvgxAHlEQ0hg61FAP/Q7fs/LE6iLPXmP9G3grIUv
imHHHKHyJIGCwKZB+FCcSsxpXlPCmypxwGfHWHFel7TdC3tW5gIwDqZTrHGA+DSp9FG13kucMArZ
TQLQWdvudpyLehJi5LDg3nE1EHR9XfSyidaLVjtaWyb08u2JvbjUe5Qzg1xBHfmRRp7hRHZRdIHR
It+d9EJRSwhhPV6fTl77OOqGCtVC5WcD26DwOL+OInuBGYr2MPhj76PatqzNh9tN1To5h3Jreywo
SDWujOdnkBtk+JnmHUCKA/xUqZNfSDDbqGv2r7TRC5+sg7cGrwVE16wccPoUfzTqkhpqiUt4iLFn
zAvISB//xLH7YSNKMCDQzmw02YX1GM9dic0ZZCXkQEjaGVx5STbz4M4LoMaPpdEBN3xpJ5M9NVbH
wQEUKSjPi+Sl7WXaa28tXHVycVWy3wFUIbEU3i06PZ7i6llFQECQ28CaDO0VpIhDaPzmBYGpiUNj
cwCpumcEBVcCTUitpeTNjn9/U6dLN5k1tG8U5SCTTB6CW+OcLiho154P++9beOp0XVw1e7kkfmZy
ILjDFQyBvXVLsXo+xe54ig/Sa58MH6BpTFdkXITBTPaqt2UatgEB8Sb+34XK5LuwCp0ImOTZwokY
lOc9odfmtMUn5noLJU51zpuIKmvzzfeIy41SzKnqR+qGXK05eSL6qMjn58zs8Y2aTxI00YOD3prz
N6NIFo/VyPDoXeyK7z26NM+AU7vohFX3PHYkEIiqJQD08fGXjVobSTLSWRZvZ4WulUgpk/RD8do7
pZIaElv7fJN//VzmuP6F4csXGT/25m8W2ybOHNlQdeOffKBZjak4G7RQdG1RI+DOnps4ZRk0srWc
RuZ0MGGAu/GIwtZdmhJnDXbV2YQtj5VBEliGTXMOM40Ljq0dvqlXLGvHQ9SB6I3vqxmWOjbTXXmc
hhVK8RCaRsLcrsngQjChA4WsX3vmj+iBOxhNZRm+EZYJR8p+HFFUEnvAnu8jT8Fy2VROVN1R/sVI
T5cDowHwch/3mAog7+NdZGJ3J1FGXMFmXDkyPY2cIhAiTUAS6B9DMvyRmHPGUpROkvhguJMt+J5j
W7uMjvQSjMQNVvz9kdiL3D8qSYpSAHHHYka/QvfaNBqo1Mg0nVXyCQ46kB0jHLDaEbdU9i55tv+n
PDGC/PzW3EtRgvYlnuPIEs4SB9TXGVFB5qRQUXXSmZZ+4og45TZInAoLgnsZvg/8sj/L2g2yuCBz
+RGwsw1uDYmiufaIzFf3aSC6PFvts1rRW6ZUoGnBDcQTOQAEw9EH1TJNoGNBGpXFhIrOAGKtJmX+
tQ0NsFxha7j0O5PYD0i+xYw3B6UMzJEOkn4SpawQAh5eLCbDDYSCH6WgWkeAxek8ffacGTU6VzuK
N5UQqHhbhUqFLddWrAJ6YQ3F3ZPj00m3SwfAa5vjOQpupIfwhTroHouaopmdhq5MMMzVgNzjsPFm
xCmlvX5uu6BmR2D0uQHhhqTMV5tTzlR5EtiORXTNFABNsBTuI37XUP12cJPVCK/rXbZcXCEIuqPK
uRSsh8jyIgda0y107Ks4I9MmJqciMhhiSoUxcW39d89prZzv2Yru7D7+SNBDnfVJiLYlDPOfVpSf
5n33XcZoyJOUOFI0eKP5tuA1hd5jwKfaROFlq1JHB9Ea79wfSoIqgE9yIMbpaT38VcRatgPhE3Vo
IALRnBgKwNn7fF/B97qPXEZOgepqrssDv80dN7QfVSLIMM2acgjRYyiMuKmiSnZO1aenwpnTYTwF
0o5uLvjObbXiEm0WFJfWpzEAkvSC89xCMgsvnXPZ10UK94Y3n00i4ajsdtFGjDVdzyaPUX3NHIvr
CzwGM5EX9EjDDVZRnQbIMLCowjvTgD9Fpc9R0vde4Fg/EwrKiGD260gBZR8RY9JrJwbpKRULQrcf
IQQ+qUs/zMiXcT4/CFLGNQeNnoM8ebW15KmyTg6mz8+aj0/LY/xcjRY1quGiDseiMxgZutQkKkv1
zufgefcvGRovr5vAJn34jgWFqBKxccARV0WMswhzxhizLFc7+IncfwA92WOh+6nczd8eCf0kW7ge
inCDVK7NjjBG3OWZqsfQjIuFEpq/+l6UBT+sIGkNfUBagOHfZM5dWSrvSlGzqBuGiWQJq7H7xejO
n5b/Z1rbz3pbsRUpKMJIgwbaMjPl6XMhJmrPoN+bo+zAOFcJb685UrEhAuI43DB38q+nJjovZ6Vv
JXUlUkItATSU1dEH+GXGd9BLBN5/gBaOVMhzDr/icXM084gG7zLbUZeCUCFt6q4uzxIeRtwS0wEG
jt7Pe76mJ18XIBsMToxtlqnfznzY8HmY5n4wpoyls8+6oHMrUfJYLTk4rWKjnKhknbNxCH17kyGH
WyXg4k9RrKbcJEaXjBZFYL8YYY+YSQYfg18hQhBe6OQqOsi49qWSvFAdE3L7pUVfjWb1p4MZZc5i
tjoecvLwnqyHxxG0LdSjEwHcXVWRs2cFMMXudsio+mIV/CiAN/8a/hD0IXbYRIymImoAEhRhRMjP
Rn4OiOCF6EV773ZybGJK11qyAW5NqNBbYiFsPzcQwvns4rpx/AQ4A88Tw6DiC+0cvSU0lXyL4N2v
B7QOYSzAFZnmlnFVhS+1DK5ZDkuaIySSispcjiGTZNKdd6mt++7f21ZCvbhmqT0ifTWoSchqSX2g
ajmdkABZosi8nrsA9t5DBkHXkY0iWgID6AFoH/7IacymH0F4Ac7TmgBZ1+iwllhgF3T/v7bti36N
ZqFYFFa0lne3RF7wnwZeV9pJ0Sr5RnyyZEO6qud5DcSnDBFya3tHpm481PRdhbWf5t51mR4W2cu3
/JH62d2lugdujcoY+CZL8UC5SB9fZVcPYLmWEFsOX3a1TkJIvvKdLPaKiFXLh2DaslOj5BF1ECFJ
mnvwoEUcRGOHLXZMIsEGvyqeWuCquoCKAYZQ3B7jsoGBo2PKg9FBC+pHsNcelz+9zZMEdWAMzPlY
oUYAIqu5AR+iqgqmAkWz1YyoZzfMYzNfOvM9WE3kzCzcsDyRGZuPGeub1+42sbPSEf+UdTBjzE7m
1pwxmmfu75Z7ehndWT0C1TfDY51keDGrXDKQH4M1Bdrl/8/sy/2QyQOF7lGgtahufxeqC0UEW4H0
sqlPtTffFjMiAend0W4v3fVaPB6id9Rt0Ppe9kMp1dde0Wb3OKmpVsXQARG4hicr+IKBRXNa2969
XOD5vypZ8hMyatBmU5cq1pmla6k6e088x+2JfeRqGfEWRFF6znc2yrWz6Ra3V0wYfIwf0z5abS0Q
dgHQ2Ftak7VgBY/Yk1u8JEDrymfJnqqltDBmRJJ17bnSfkUzIvVBXh+2CM4cldRZCQlLK+j8J36d
L+MzK3/vskcPUNLAOQn2ZE8nb94UYo1mPi5QqRgmaop0HuEYAGhEDnDQEtg9t1WGGr7IjHZTEwgL
1NqQtHEmA2MtGeWGndjXEvRz1X8Cmcp0+QJlJu3XLRGAHb4u1+/MhUK26C821Jkd0P1UAcce4pFT
3XA3wcCeQ5+T/SpHrWxGiEJq34enfmqCLdDY5kkixUXEDa8kiNbQf2ghV660OY3GgmeS+o3Q8T7Z
2m0e2IFW8nKyOHlkDDf4ded/H40tBOJC1EGpCcAmzskHFkWUI29CczhlWX6Mf0eKpOK1KI8ksmvW
7j2zZyx8pSJk4zq8eAhNKWaFqxsyg6L9avl/tWkqrnjk1S4uv9FHuFGA8jVFcUPaUA9F2WaLY4WO
ZGuiy/YO9FrvOnPRnBqhY52uWsBgRAsjg8u6cgkz1SblrzAldOCD6wPhaKd3ixEYHnkvp4dtNPzc
4HB4HcIooO8ntsHEwbh06FFz3B0zF7O7NRgWiJg9wd3/y3UP10QPnzoOoRhg4FAoZs4rgD/gvLdS
mz4q21j55oI6/4ulg8h6Dy6O4Dps8XUeBILrhbZzmOF1WEiMWuG0fRfbQN4Fsd/w9r68OIko1iwn
v5OZl2E0bnrxwbHB2X0zhUEX7LdsXftyqevhf3JOMNBf+/lsMfXA9vKHZuNihM+KmeCtfPQAXjw6
BeCj2EpSEpvxonLOHfTbATcfOkSsN6qBKS2Tz6qD9SrbX7zs7eMdAC8mdWQ/byWSMczuwZBGWBcB
Vf+c6U85OGQCV4Zmdc9Ao+S5E9ha1z3sXQNXh8RfWtW/+o1wDfo1VwVPvcQpE3CyNCVsRni67+KM
BD1KiEyBGBB7oP2PGyE1obiMczPf3IHFq4J52fhq3q/3UcaJWfWGSNfR3SkKsjhLPfXrwuFMf3Rq
IXezdPwa8Coelbgs4N/0Fatf/QInqEXQc0ESkuCH7CGpTPvcu7SIkNVtz5T1N1xx+CVxCM2jqB6z
ldUvnIHdPLy2avggL3CbGEXIL7ZH2F1dVmHhIn+t0nyxLRZLSbK753psTuNiVJzvP6R9UnBLNpMx
6DLK7e4PTEXxRMQaI8VGxei0I7hOIFt0XbjU/zbmmr+l6AdW3UMi6Rgml7n/0CfGcgKkUGYbetH5
/EGwdfel3Vnns5UxuafkNkQHCw5Odn5+CQ+MYf3T4BHURFz4EjZaySVpS6n/dxx+4RIl6DuFxgMW
tnGQSuyahoSLSpND2w4FvoER4uStlujf7Oq/PzlSjUKK8o3RX1WFlhVL4t9zhs6VCS+cyuD6QdKn
9sWDU8TOLt3mHfRs8OeAsR3946AkDsxibMOqiGPKSArSUePJ1v0XUO8U5Mhobw6bQ2Uf/qXezUOS
T2E7oy5ZgKlPI0myX93weXdV+TdDQ3O16Dm24/AEdGBMAF/RFTAwiFyavMhP2EFjscxRywIAX3Mg
v7l0ZBn/GJOtpLFlJjhJkfkGOdEytnnydiVNFGpcbx+yjjEKukyEKomIkzmeA54fiiuITU3T3UNs
ODKEUbr3ZW3M7hHotUADfgezALvfEA5L8FM9o1B3ASAxF6Pllt9cgkxwJ8fldHlFWUFk9e/Ii6Zg
/eCFHlFZUbjn7zxFRqa/b2QYNqwcxOD5M0U/zLhmENeJtjX63k7vBgKjG01oGAfDiH4wb4iV5xdK
+cCGzI0nzMBpES97pQn4azmvY0h8a/3ndGmGGHwbDAUDBbHhndbUMsBkUm9zqvCPN+snIk8mbm1f
YynY5KsMk2BMcyQ1Ds8h69N4pc0/xdmHq1MmjebXYvXnnZ8BVW9W5LbuMsKAq2slIkFkS2g7wZdp
xoRG+bkDHtLMRLZcOn+DbVemlBT2DdrIMAPT0YdG/x3xChtVwAfR781VzpGYDZ7WNZdrQvn4yYR1
u3683iW+iSSTTR5owP2qDnPQrifVHwznqv1DMxzbgdCyGpgV/QwGFtncAMDJGanISsI0BluulnCI
Q6/kYX4E8letwv+DJeJcfV8qowhMK/CpYYLT8xL1WuKqDHP/ToNzcYsrXmEVvoPD50TRANTpDrk4
IBBoj2GFdCspeKks2GJhg/vqydGinJzeVK9GzS9xDSyGoVSSFeaLY3dcZVwgE0MS1N6nFwCIp4lx
F5KHFjQWam7g99TOQAefvWE9DAINHgv3Yh8B1kI5nwtBHELvcSdHpxxjsFovltlQ1l/0RlxTocEe
YX+P4R7/1P/F6Sf2qUQVKscgyDCvet8jb3FdYJTOYuRQQwSxWtBfvdg8/Bi4Rmyy8Nq8z6APQ0pt
Tl/fMIyU6Zyv3o808yFOZ0dLmqhCUiVQ3KAG0cEm4S9/FGrp58qZSneNJ7RC1N9ljdXCbiBOt5YV
466u2NfwhW9tosNfevXnB2iPKrPlh0tlSDtuzGoBFTkwsROcB2hYN4ovkSRDol/EWHVolYxo4lEn
iKTsX32zOCl2xGSOAOxpHtRKfMWirvM9yeFg/APh4aGcLW2dzY8eeVgLAUaz9x8anz4YK+otKOLN
oybYp4G+RnRcEiiZ4CpEDwf9cv5L5oOFgisSERB15Ay9+GVIV8jr0ZYcDFbfxHqb0Iu8uO8NeBa9
Ao+ItSe/rzAMXyXG3H1c1Fqw/4zZjp49ulQOhLmgHWH57pwXdOIjFsOrY5S4DHww7kfCC09ZCvWA
fcij+8UvxydMT74qBuMRGaZ1cY1NsMjEaJrvUwJWmxMMM3oZvBpfwS+ZbTqH4Z4HAbQgIZnPbt+w
Y6OiTxy/ShLbyKXXm4RmfRsbv4gpWx0t69h8AK9FSfhN47AkEu1Bhu44/3bSRlPdFxnsktFIjSuo
EGCEYUwjXPpOBufzEbWntE0a6Tb0ZxxHanlFKvBCsmYnF/qs956BqUNBFyjNP+5XQA2xkvKuxr0h
0yQZEGgBf1uzNFMovBJRJOa9r/ISt5TuTOQguiFi08nDMHHTYG898HcxgbGnWCWwPWDx7TOaIA4m
jnGuya6CRUafh5GLHJhz3IlmVlS2bjaOhS5NU16IIJKk6T4EPq8KLyXO7d97YNNGj2/njQ6qZifS
yI7SBEdW+kBxIH2kfxljjpobHXBeVxsgd0TVkvVx/6IjKkOWFemb4Ww4p0nf2lqfH6C6zWx5fu/y
Lu7tRcGVNVKzEQr24weGGVWbq/pQBe5UtrWZyNsA7M+KLTpxriNNzszMUhr5s7d9vIfIrklxGqFu
ZMUl5pY82KtoZHBKm6o7DlhFZFwSRtMqu0le6XXCZlB16mPTcnNQ2OvJXbz+w61Bc7hgYFN+byez
YBKu7NttkznM9jlwAUSnJ8zwor2pzelQZIOBWT7Yc1NJeES3CShaYK3JGV33z9evXPgjov5sWyDH
4iRp6n+ihpJ9ObZ16sq/PlgRjvP73L3mCp5QWnNDxLgSyRWkVbQmUTE4+xsnw4AAeVf/WhyUgGCx
zE9u9LZYzRDOPQdp/LIy9/zRuwUtYFghAf37RGI8B+APIe9nsCpSr61uBP7QMcQAt8VVNiclbDYJ
hx/+LG8MOD3m5ihJLY+85dDPpQtC7Czw5/mGrnE26RuoQNIaRJ/k5MDs3OOKjhU2SYizhfk9lAPF
OcJczf6wrHia81MgW7UaufNXzqoxOHR1RW522YI1/HHjC2TYfzXpAp6SqHJy27/uYm5SxZKIGdmW
8/etT354SCJuZUmXfAEtjOPoo3CVefy1LpA4XslZ3gqcjdUh3KC3Ke94xcPObqnG4jP0c2rBD6VK
ptMKGjzVyQkquPNsTTc3V6E5vo+rFhZF1CIRZLXrIHiwG0cL6W6moCVkhj6bx5/bjl2nOEhhx/nN
5RauBxZkfCqk1e4TmCQ9jfMFpo0k2yTexvvYlV0IYBW6maktcViZ5shzBDTIXvAwsGBrPPg2ROtP
CIscF29/gWTOEsjYpWfgm19aOlyW4OMmbd+dGeUwv6Gp3VFcuHYOd5kEJC53kKbooRrTb6Zgrmma
n188IIvKorBQedke9Z1x5WuBdzG+BLxDFkJFTvQ879zlYOVnE1Jg+AYF/kdi5ioobRrDwVgCAWg8
hqkcH2Tma5mbAuyybnZpaWPpH9Mb86YU1K2nI4cvClyIsEwBFC5RxVVT2OKinFA9gTnTltQUP8+X
qnbbNp5GrK6eaRzLhQrPBpqKl8+rAv3epfrmqeYh1Os2LHGJIMYOY12ZdqAQMEEb+Pvey2UTv1bG
YNBcp12wuOMEGTl7ueGYXOQIzo4kqc25BOpgun0qExffqBUM/qZeDG0zNVhIt8Mh3di/dsAesMxU
qYFL/J394Ga+SKpulXeJbvNQoOCAiurNd8VdlARLI7yh69PhCxs17Jluu1O3mlWUmf78spYUz4f3
I3YX+AcGsHUJhOrNkwsMkN2TKPbZPyCSvGKdjTzD4ItnT6YwHe3ckNB0RTIZWBc/Wg0QeTKs0kVh
nSQACVrktGA/9tP4qJq772DZMOu266WNwgHnGRLLa8Tckab8XcysQXZTa3a3dO+zhGQLxz9YpXAR
VWge0j7tjlgzm+shCSiColBUu/s5qgQ8nwxKkRzJAugSuQWcC0NRe895SgyH7vgE+koraRvhIVQm
IpaI3ygjegKo5jvbDj+msTjSIreeE+Lau5cEyqieQBM9iin3+NJ4uIeGvUkCvdj5bMDG3noo2pUm
gKbAvuOB2TF8qtHOwwYNhcJxIfkZZy3EbzpiItWhuxuTb6w06Wte5snmI5sGVHqk4hwyS9MF70eF
sc2C3gHXfe4AO6pZRKskNxKXpbmxMRojrOV9ukaqwUX4WoztMXgZEzgqC/6jTn4f3IMggaxkdbVA
fM0X3/Y5jSi6J+6VrwYN/Co/Kucv4oYcEsPMYMKyUVe6OktnlBq2xILlwB8xNd9JtqvG3gWJHKbs
Bk3Ox3v7LrZUd+ZBzxH1GfF0/ehCwidCjFHoDQjla1WR9g40zqfKmZSkR1jCs7lNUOTwewG+H9eT
Q3zWXjiq/LgPxxQnM31N91xkLZ9MDKDDmaJQw4EoO/WiSRY2NR1iQSFxmCnQaVLGVg/6SVvJyd94
8qTlQU0LU985Vn/MiOTm7FRKF1Z+wFCco72FG6HZ+UBbzNKFJNEmci7d7r+Qb2LnmrgKhcwWblot
0aVwAy53/NIe3lU6O++RnB4qZ6wLUS7UMphRAs2ZHskWdFSPHtQJDjwgDVc1j5e9NgHaILT1Rlr9
B13scQkUlf2Ov998GQqShuhytvl1Zh5LzzLUp3y/3r62M3L7M+88ornzNh4qse3a4vIaY7lJkA9n
taZTAXjgMvNFIVTZt1zCYR4LmGoyDP7V7XneK5f1N/AB4jV8Tya35L5XHMWpv5Z35vG8P2j660TR
hha+pvS21ahwqntpobq7R48I3XQU+nv3XvGhnRc9noBQaPGNM2Y/YikL8xcvPIRYLnyEjnINjoYe
9ZCaYo4MGxWQllW9KSUVZ0IcFuOv3JdNAvLFfnVNYxBtnqqymHnzoH50HhV3R9aJdn6ENAkqVqKf
zIu+RWH65x/zXmzlD+mrGxPdj/PbBjQguclqh4DkR0J9r7cnrskVjQkK+pX2XEGnMTXrefkJx2uZ
bQW3txlHXGrLSvQlFY35M4Ko73Ta9Ob8WhU/S0x6Gs4Iaixkd00VpuXohmPTqfLKxYY50tJKspIp
AfT1Z1n3yRq3nYtZBVZB0Axa9cHAkTwXIwUuh0PfuVsId8jc/xnSLvyAWgn40paCHuQLkqW0de/C
uIZ7OwbqEe6DPyjJundA4kQ+RZ/ZWB+RGg2558Kjz9fHUM+kQVR5CSocryZoBD6Xpzt2HwMrJksE
PKjsa/YLil+i2oBYd0wn/Smeka1XbKqDUK06pOzDEWcuZ4lgmb9R7mCpV0ynJPwZdRb1sPQQjs2G
QA6AB68gHVJZqGP0x1xkS2EDY9GTTHo/IKvcRZv6rCFcOC8tcX2SdMiOyP4G+V+RhEEE8odILwIQ
p/B4ZQd5X7JntYV9IUXB5XMeIEgVUyL0X7XXIFEiiLDMk/sWDzyTC9b9DWc4xW/EHd7y8cTgyPoC
czeLRMRw994FMEA7HhBOVXboaaXsFj554HyK8sX5aRh5VoWOKRcTwbQuuj1i2GH1t5mNvm73psQP
lN1G7eEnjCG21LpvDv7PKvMaJrI3BEIQoP0UEraIRfLMMt9HoSvphfaAw2MxZM167/AKovlE6sVM
wYEn2VZ6JAbvR06m8ErirTcT5v0PchkxwV/2jyIx7T0cEg5F0WjylRxMda4refj2VJXCqrq4//eh
fnA7s8MIRyoNFY+GZ7pZepm8hTdyx6uifASu2ppz82t65Q/Mjxs/8xOoOHJN7b4BgZN9BrL9wNN1
IOhe6GXBx2xUujIq6me+hGzjsKNK1BPkx8X5oB7zWVKEF/qgM/3gqui3JckIkDEbQG4V0WoQu2/o
p/Vz23ZwXGGW+pfhUESrWMKtdPO7mTAwAXParLDOUM4QQtqzTe1TkhibDLaUBpUjsBMzvMvKc+Np
SPyD8Y/DhpC/acV4ZyUCY0kjPkAD26n1MtN8IWHjI4mr7r/fxwAM3Qx8jZ4wOks83IuQncEV5Gd0
4bazRdQ+IJCcUxfzRBW1tbAbBiSSnErcXtxKl/jTmWusU44LDfuDDdRaRkyMur5DMy11PmiSOyAc
jly4EomR/xzomfYID/L0y6pn2PKWXN/3ZkY329KrAeI/je/gqvhUkn9SYEjuKu1OBqgAPZyJR0Hw
i8cVvnPLo7FUdtg1JR1DYyTMwCJ3R21+Obi6QaSdVMEkohc/ACh8fuvcjrPZwFLGq7n/WNldsgv7
8NqbmqIGgjP/ZRIroCc1zxpyw6zv8ahPIuiaNUNcRQyFukXq+lWfMu4/4zSEdSl+9a7JbLnKDHoY
kZp7UzTLzhenE/0OQEeBWWkI6iOX+T/LQgXQ/vRpFw+JVYJYyqDVSasxaXlvTKl98WF6rpYLYy2+
7ocpthi3YFk5HZ7DCnUf4ci5rq3aa6AT3WCX2t+MzC17AodavZ6+GI5GCSLi4gD7BScrKQxBqdXa
jAY4OwSOBIWcewAeBlNqpWLx99rfMOg7XfwR30/SMl3XcPLL8h4Zdivzte3oB6fs0QxE7njPVSg2
+vVQB0KN+4XBKfBo2Pf6qmXDP7mob5h+fLLNAt+89Jyl8ecOu95J8Fv6C552LWzVdqTPhAgOS9WQ
8zBjNFMfTMe5t79DsGYTgnTm0C57gInixFKpjKLqNkhqo85ZSsKeBUJ5q9rJbtau5ipLKok7BHkA
glIG0HB2b5fcbjI3gyf4DjLW/srybzhwlUc6cRYismN665GimnGzU8niJbeGvYKaWcuY7OWMTzF9
oBKghGzhd6u1IRgUvQIgbu7ltMUiBGfnbDKoKNFLSi+rZokt8MRYI2RvdLWtFpkL8yew+3DBJOr3
8PYZxR/ZPknHOEZBzf1ZiP11Ivn/lAxR462IswHQRd0HWsDYw8hSECaE4KNq119FDs6dEgG1Rkqi
306M0jqrDdTXPq8U+QgjscQhGyhZVVnlZsgxBJzfX9/IpB/NHwumZINlEFzVTDq8hbwb+SOQF4qm
rJzEBKhhiWGx4bsnRr1gpiYtuQ4NBjyN1VVLgnu1GGIkje1qehxKNtq73jCiyy6c/ry5/L7rd3BZ
KhpT2MGiafpSs4l/RU6Xzw81Pj/3g/YBU8+si6DOMPHrC5VqmsblUaLZY4PWVQtZw6MlAGzYRWm3
Lwllkdg2zWnYnvElqYyK3LlQjThS1mtQQjtFlUSmvulJYzSciHxF+O4vyJhTVmHnImn470V48bTm
dyLd14NmKW5HO26Ow8+eQ/1EHxs/kVJq+deWWiCYAU173xS4zsl9GZJlewLQl8PuUAcVPfxW2xa1
IqU3u1t1t7d5x6JfO4r8WVw2ZCJKnT6w7cqVa0x4F3f4SdPMeyFSPp9hFD6iPtl5sJh7A0Pre7fJ
Tc+fL2IoOh8/X0r2m1Nyc1V0gj+JLyjJk8LqSBE2xE1TssjMm74FfPKF16FOe9Ir83iaLzVJRC8N
7y2vbtwkKUa2G7nyXAJ5e4LZR57TJ7SO6iROR8Bs0Whr05qi1xTwUTyvQHHktlPGJzkIjIDvXnzd
TtKm8kc0k4Juf3lLwxS5cDmC1CpRNkk7wMJP4B9sYA87KKq3+45w3disNHD7HgYy/fqf3jNXFWrL
wa8DHVGwhxCtb2Po2TlJTafnPzDSwYRUJOLagNw0+MCwNAb7wvLvk2FrVmNI+QtTamw0QQrEOnnT
2seDs1aFPq7oGx/9nJhnI+7a47elA8bGg187YA4Sxtz4kILPG0GY09eL3HwWh1kttDB5aPbrTZy4
kjASDj9WzPt2V06ctUg24bBFIsgpnzYa7FOSQT5jRcYMWZaHheLmHS4vsn8M3/HWDgvPczHM/WUo
0VxmbFGRpYqyAqZtHUcLxzQ9u4TIj6QbQIoGGz9qvzZo6c2w+XWaRgFUd+vCUAPw1SZNkqwpdDD2
JXKzAllTQ4ckB+80awL6WOgP/lQTyobLMkKoYPtuK0fIFEVMVwunJxspLSWUGMpu1MopVkkjbtaB
UUSCKzbQaLpuw5nsc9uAWp4G9KAwGRA4TFk9IcU1H1Pj197JkRnPDwDXlRiE5/SzXndLhT+PQus4
hWL6M5S8CFfClQmL3vb0uAbx5K5alxdgTU2i/NxechUDY+hUE7gkvw2OPo2yK8RrQlZIxOmPRF8s
Rux4xrlyKTYPDTBF520p4tdw/gsWIk1oqQih41dL9RNCim7XQEmqkdFQMfTvFVRc7LZLVaxqLZkj
MiLRNyEOoFvI0D0e8X1J9AQ0WFSt0BzDC4xw1A1cP9LpnL7KPtlvrfWpWIPWCG08cInpUDANHoro
cH1/+L2DWCe2RpqqrVtiyJcs/4wI9b86ArAQwSMFPerOS4pSaGEBrNS7/qF9Y+mIyjVLBzhlAT8F
sp9iVTmCXLF4IoltTCwoUf0vDOw8lEa7bIbHtojJdzHywIqI86B58LbSQ8KwtHoe/uPxTihEERx9
zQGGY0HIrUQKkepMngyCEW+zpupeWb99xlhYFzWcSEwC4oy8NJfQCQeAYuUVhhwNCsM8UkrgsbHM
/e78Z6ThGzz/NCy/2gQqd+NyVfkExpesBi1zbHOCdUnnkXE7BuBCVdbDM7ya+PHh+xmfoGJBABQJ
UfLwREpD1UVGLG2ZEPKa22BG1JbpDKX+ngNFXVjdtcIiWUemuY65mLQRrYTQk54lo5zEDw/wBDsa
ZiTElQgRGAZXkOL/76FMxtxyUhpz7VEKTho1m77DVmBRsXC7l6tXZuyoKiM578NhM8VEazKqseZ2
rigjv0UPUGukC1BHOT6C6U80e+D/3iTAYKdYMdlkB6wQkaSe9WioTjGfJfg5UMgJSxWKXLKLHMAx
vpUC9hy3oyfvMdYdZeHwpf051OL5zst6CJyb1DFcd0FeE+9LxMCtTHCA3o2ENoPlTHXFFzp6Dsvc
mjGC6L/EnnSNEm1ccXq6eTtWDfHZyjgNF2BZnn9jEyzmwEyXuv2LEXugclTIh4lD0GXFaACIYK+h
/0RJFRVL0bbB8QkQIRZ8wh6pdhKvfwq+PFD+N1iDeYdhkB4Z3no7tvcnWfmLfJy0G2HEMR9WTOBA
QxYx4zxAu9WEKM21bgGIsbOVLEE+vJB6KyXcWxM6bUAJUwjAWUzwqdFT6MeIAEyNc+xQxugKQOq1
UR2RNhBLUShDrp1UWc74oM5yhaJFKkQjboTtDvpVSAPcDiTcsqDMqnqhaknMDj6rLEwqeCTfaMSF
MCdWGQaOYCnWTd2BAKB9qEoI+6UhdM6ilBW7R9t914mnKnUHAbzACKArAcQvZuvyT7F+UMUZm5bv
yKWfcQZJpMNEVkNcKvun0e/YBaQZ7u3Vt1o2bVg9lAvhtuD1fl129gInlhP+OfrTVHZECdynIsoU
6r883TTOycu/FZXZdjAb36CSdzVQQ6K3b99RKIV7nI3vwcrAfe2zqMAkLjFJO6NlOgt3+UdpCaSk
vgG2iSlqKhr0v3y1l1ZXxiZnl/iYog0qoelSZnMH2PH5ZNfuVBxdSElSPvZxFSsZQ4nvRd9zhiQ5
ryh5A+V/H8W5dkWa5xFonbU9RjId/0p8FnnhIcYQuIhIL4A8SFPfG3QcyobssAz3NcOcvAJdHqMo
Nvm1UaPZc9vhn12kJj18UpT9pzlJ4ADtybzwD5GPgDjpvWi9gfEAGs8uXH/25ZZxpp3YBQSYhUso
fW561Eu9ADU3WPyaTrrAED2WcA6mIIdMBZ6KVvgiZ+wayvd2iFH3VTJ2i20V80MSeYEQxmTmxYdC
vpF64GyyJgTeYYSy4khA1/lXpC/OnO9vuVWfXtqCOFmHaajioItC+B9F8YT5H037+BDo+GI+L5Bt
WxJz9M4mgNz0YAylc+8vVgdFxWCSUD0EJ90zGF/4uxiZlIN9QsUCfiXjUjQsn4gFXD82g83nCLBa
eXGqA9QlAWF1ljQYVmejnivPaMmY7Y95S3gF3WLlzeTxHx73L16Mjm//rQ2oqEmC2I0XHs5zpnqj
Geqxtz2WritlFkRXYiBd/9tFFHwTij49hSTjZfAQoA7VkeAHEbiLjm/x66paHArJxkTIJ3uBIOi1
RXKdhJl50FuRS9Q1CgZJkfB57fELxZSvVfT0hT66zbh3nfZoPn3W3i4ecrhUxAXg88KIhn9bnigu
uvpN0gIhIvrNkctWhfuV2tErNt37uIR8Aet5A8o9sDLUreDaki0d49Up/J/COStR/1bCwi0n/XWU
9OYEsm52/KAuSPytcth2jDgHaS3AH287yK96G4W+SkFYREYnRkrNg4AvoxJU8TkNVN67/Ebc2wJL
PZUDw0/LLaBHqF88i3sX3+fYqHaMmunMZ0ZFjQqaGVmJuFsoexwnHBs3XFJB0DnwMH1yOna1fwsY
NJ5gyaAdNSn3p2KkrdGtAvEg72CM/Lzn3lHdVQiqCrEPLIUF0BJLCk8W7mtYOCTqb/jsXaDA5j56
cNyCmLgOZzVrIgDJzQx+OmpgTdkuGWFClu/JOEZnnZqz/wV3qjdnsZLZI3sEswR9VjhY+5K5uO9c
ndLc+JbxX6pQ7fJRnCJR/j+y7Lxl8fes2ZPkIjuWf7bs31vlNd7Qj8dXTQ3IDN0/oMcNfzoF2y9g
SAF3iwehsJbyA/gH/XktLbiHKW3eCQCkB6NsKk+pwf3OZbfDaIrok8vLcK+oDv3biQNx2afmnDED
/+vY2Gs11LhX3CmzaNBb6yqeDr6gLg/iQjV7c6sWBdAqcgAGy2UDPDOKPtVooe/dZy0LnZZ9s5Kx
CvW4Oyd+R85UtH7mDwzNbnrYwMTmR7LDEV9y97shy2GYnzCFiQalVga27dSNkEEGeOV/kFM2jv2f
cin6pma6WKRk3bsz3WARI2y//ARUEXXx92vvbJvqpY3wDiVeNWuYyQWUk/FVq3yT2VZ9FoWlxfks
62CugbBVEL+gw889cHIR+PGJAcdXZHiLkF2XhN7KLUqWdRDQdsSfy0CeXTBKEzVXXwVIG8DfA5qU
rSa92pwmezCH0iOBlBJAp7cQMqeSpcx6bIIWmHW3JN1GNx74bUqPI2S7tRGS9T/nia2xswKA2RPu
LC+h+1hBRWy56DbkwNzRLC/zu+AT/da6Vv3bGLZ15Bv+vpxyC1tUHSTaILHXsAkT5Xv0Y7ILja30
7zY88KeGBs020t+svFu6mMNXYEO4XZMgwGpfzOytNN7QhPi2CcMAX+XTuZGHgSMJthtCq4UgUam7
fJt0lujeznE2bZfZE0qWWLJcsS3QdIIKG683cNwzkKIrmkzlNAhRutGR06LCoZEdJH0HUQYaPnMj
ZRl3we2W7vLnI7PXYXU9nXjnPqhz6GwtkHzfk+7csEzh42JgkOOGmSdDePfsqZqcdB56zptwqQwm
5GB6BF6NTg8gTpmwtmqmy/5pvej9VKHrHxVwb6nqd8sCH0TbHgyXnMiFvuvOfvhzCewI/8mL56d3
MCXjdFoq5+ecT8Ylpc31ZEMWfD+YFrAYDCFBmJw1gyeDmwTCkIR6tyUoddf0XVhDPN6hfqpAWAHK
Ck6SMoTEBBzhoVniSw/LrVXWIs0mb9ysjALzrZLbpbpQryVP9AuyT4vQ6U5dWKiT7TjqMGKXc+Vm
HtMnTfhetqXoBeQLJ+OVuufX7x9AlgDraOZZhQmUvVDTQ2kFasaViplO041JovrwyBxGWAQ71/MJ
hAzzG780vOBlphFGnNipq7cpsIYjVUkx1VlYwfoKV0uCbDrm69jDhykS+QKlWqAxCMX7bSGtyReh
rH6pCgbZbZKyy7PFUq1FbkPVg5wwuvfFgeMobIgfQvxXmDCRmZaQMOhSWO5gYxY+NVyb4igVTdy8
2Ssrzd1JpP6E5zsPp6Er16a15ipoZPszYqzTuD5OP3+c5uLYUf9D8p4ZznpjQIGr6PK3/WGnytU+
cK39NSOl8lJwF8HOo6o/GLWd2RaPG/u63aaQhKxfK1Y2+wPl+wTpz71sOgpSrxkeMTZgNP7gYGIt
LppRkikUS+79pkfILtkIOpHrs1uDaTMT485f6XqgbOBk+ZZCxe18DhLVf3e5Q44u1WC4oYwU2Yya
Cf1BKyIl9qjFFbZRa5ADx3ZtmeSS51pyP7rf/S0Ou0DyhsZH9O6nL/P8nihZ4pPDCPmRvn9dOwJy
p52SyIqZ4IzEZMvbmav8fYUc/ncrKRckubeafOiymWlz2trEoQhyX9CeYAtapyt9DtO1wkS3vrPC
eQSBAEHNeBxj/Ot8/EUYqim9gj/YgD5D2ZPcG4iprEntq+mSTANvg2wUAdcg1tdKIArWuqQgPabf
bnVQm9lg15LXcB+FtIfcLdDERwmmERuPj75ZK0cdRiRUKlINlUEU49fIpQBWJZ2szk+myynCyxIQ
k0ccknv3Omj3bMnUDAr4YDegVG/vZ4VuuUg5U2oQaJO0I90Xv6KOOPcKSztl2ruii7APR+aAF08x
G8hJDa0zWPSeYPA0qxidURuCigIvjVu5eTL++CMLXARRSLIqygVqcZSmayusFK0pILndgrU2Ik9L
POzoLbXAGoFjs7CeOiiZhCuTAOIvCO4ZEMCmLjVSzrl2NKTJGxFDyxlFaQZc1PwRMpqCgddVdNr0
SGgalJ04xzx/ZkWOxGuDLG5lMVMlwT05NnEjllAd0zSxLDQiMkbXKLM2vDSghT0hEDahChNJUjO4
MPTP2D4Cb3O0Y/hsMnqIeHZ5zvrsPL5KNPPxGdTGo3NLCn8No9rQRpjGwmB2tyfSGimF/tp625g2
+UJaQkN9NIyuwmlFecBl/VEyZ5GODfD9dU61JDnIkUuQvpVkWfPgJR4fmCiD0wYpCRNgi0c7yeGr
i3ZclH4E+9wtCfHwtqJvFOohJ8c/jkDomElA3RzF09N0U0vkwyvR6YrUT05dbyKu1FIDH4bf/yKZ
PuofpYYWE6DEXQ48M02O+7aH0wFIqoF7TjEU6uLDtuxQxzvq4eAVtfDmRTXgKTkbmMstP4ym15gb
84F3tpyXjqLM6YgcMcy2/ntgACouhmErZAnVXbJaNX9fKL56PW6keiTVL0gS8iolaa+s0Lf/1bS2
82Mr+8G32H5Vv5h0K7GwO7bz1bpgJZjpfa9v/GfRUhbApydnRGGvziJ5sFPe2Bysmm0JLImTpyq1
WtwzCslDpiomtbsTC0+QV183OW7WhI/c1GcbMSIdhto6u+R8yvKpSRfOAOyQV+arZwMxatlLCxxG
TIeMESW3royAq595JVDE1Xdd3dZXdhRnwBglB0O9KaXPXZxRZ94GZLQQioJORCQniPNpSqr/ZvCn
gakTazIDrWM0BXfWfkY2Sk1tPiTIi2utZCAsji667SxHnRnjSfnm3DtZJnQtNuGWPjTp0DiySo+F
xKmVRdARJw1vIveeSopfAQIxj1OC31tutm8g5O8+hkz1rNV9m68deqt463QiDj7FaReBRc2gM2LF
8f9nnO7tSmr8uIAkeJ2ufODFm6tWmH2mRIgmRJW7ntqYFbNQ4dYqTxDVWcN/KyOkqXsm0PiKb1eG
CVRuEArXUF6X026boJ/5eHD3SAI111IGjk7DhsJrhxQNRei5EekGIft1E9VRhRk2vsteaVRHYNFO
Jz5IHax/JICHHU/D7jnClzlKzsETWWjw8bEIgAcAjYxtbWOKkNvstt0euMv5q87UcGx/v8vJpkVh
nAPZKEEG5GKRQIkaQZ4yl9gjdpUrS5rfng8OfSXhU9cVJKB51/BdNF3W/xX5SgADN4D64Ci41PW7
S0FP9LDmXmcOyTc9cSr3ajoUguG047kp0bGHT6wjO7nkscG0rtwFNwt7mCfwmpsUILodT/brtwnq
7wpXLzQ6/3SLfle+vO5LHj1KF/zNp/RoLgVNzWiuIQnZQPpEprs22Y2DmqrOaZeYpuHYNTKrO1La
gI6t28GiK9zUbXyjPV6I2bCP4WUkh0pXTmnVMj7iD67scLNLBbNVf3tAorwnKs8Ppw75dKhuK8o9
uoDT+3XkpUo+kRCeYGf9dBcnhDumzAcdAAWR+Q1w2ZtraPi5E8q0LPvSEjLBRAPeqngZNe1GJrw5
HzCqkucJ90AIzxHT4l1VZT0qKS8y+hcsy0/EjEuZcYv4TdYgR6s+nIRVw77dWzd6UPznvDGee98w
vPslylKTuHqSI4/tBCEqP3mpoqEapC9C5gyapE2RHGkS1sMTq6xylPBU26FwTCekWk2L0griUlI7
LpveiGjg6WPw4q2cJCkWWFL89ogdDDdcZFIrjgZLiLdJ7iEUJQekn66zLHB12gZp0BkVLVlMQqvn
F+Afrza4ppzYSsIKH4u0zDs5zIpceXZpbgCNyFqWqWC5dGNR49JoqycOwa8JTSbDzaAy/322MAJD
9VWKCRC178aJFOO4r0r8FER2NOXN5i5yIZLyTPK0POsZaeht6q7AEa3SSOxld6ZmNH9C2pUy2ux2
uRDjkPeLd5OGcr2WJkzoZKdVsjh6sNsyJ7ZhLkK7iYArHc6aGig7eN9I5B4RztL8rXUXFz0IYRrl
1+oEcFcnsTj6SYJDAWrn4KWRjvURBQwRbD1qZIlhg7tXhhDsNYiWGgs+0zef0bpgcFp9X8qjChuc
ZBp/K/06evJ8vD65KGyxDkb5xvX4D/6dGcqlMrliYBMJHWjS4uKYHBJ76eGpQt81Zcv40o7+NX0+
k67OOP/2OI9HP8UaFKg3dY0ECSnnVsilBi2vRj88WSZQmQOsqGdbgdjrI/Hc8gm9h2aXlz2/zc7E
puQ6+FuORxnwxSnI6X+PeMrTx7ZIVq0zWg6D3HKBzobKPoD21cyf7xSFCdjZinAptzF0ahvU3P0x
6036zuyJMGXc/3ihZcH1hwjj1DnucH22oUTDhb4ck8Z/1R8VLj8jmRZod4/l75NLeBjj2zm8y6Fr
zA75Rg/C7733uC55RWRS2fBYBD417azyCXJfa7P8CtOCdywSn/PlFIIrXvKgF6WkG68piPAen45N
V6y/zQrhu27eSaDapyvAX/IAOp/Ca/l/Xz80pC67watjhTbQvcA/D41SpVYcJCQI1xPPgH26zZHu
METBB1MPwVve2kN8RJciKV+CRwiKUDQfX+PhMG+eaCvAvjX2ixUFnUyW+dEDUZkWs38JG3TCo34Y
UBiPmP3DJcPONzvA6pVxz4PyIAMPfDpGUWk7FzlGZ6fPKBbbMPI3f57I3Tz4hI6ov9X8vZdRW0Z5
JalfJfS9pe7koCjkK6IdM6/AYqEpYksfCWswhrXDztYs9XX7lF9UwB1L2iOwGTipdLOo3im/R6Ql
9+KlFEwYuXFkVe1KFgnDkW2lX5+CTQoVo8HarLyWLgme+vcwrhbYFVobhzLihyCpVC+RxRvUpkNR
Wgk6/xjKIs2GWFcON6r5pBjSggGsy2cGh5CGnqC1gdhGCkghPWOLs24Lv/FcIVzmpi9dBTziwAY5
GaTspkzxTxFVPpWlhhgNAUEf+akgkrDv+RxXkgGzX/mSZBegeFbsuo+Vl31wxOrlp08Mf+iOzzGe
pyDQBji33M4lY6yjUmYGRdNHKAuXwY0zRsEd4ShB6HEr6W9be0sIJjm1MSN4kRW73PKd4BvH+T7x
ie/6NynbGVMEPAIC6cf6Wb2a2igSAHU4Cr0P/gUH/B7p39L5fm3dv4qDHbN8HVdF4kXqQa4CksI0
eGZ2B24QP/AhaZA0xbdIop5UKOwtQEkav+KhXKD0t2k02fDQoMOV5lGOMTDJ3Ch5pK842/uByTSW
7rlpaFtTMuwQZaeSQGNXKijV0r4oM/p0faFqzhv7lmfpt+uWEJKFdAz/wc0FnXGHIGXhJlRZQTRv
nH5jv9umdAVE4abdNK2RdXMTwwEebnLR9hKpnR5QlyAN+izsOnAV6pANdAFXAx9AJc05AM3xtHsZ
gKOZsLtqKPsuQSW5QHABtrvrECwFUeOA9/I2y5fnpvg3I5xENAmR3DlXtvnPhada9qybAMspiAGX
fjHEZRYwggLXoSCYIRRrOwyi3mRAumUnbaTQFrPo3Zh/84z0w1j+NzU0czdYwAjkespGNJdw4HXH
vg5iSC3Njd8rVcvDqW5DBpH2sZajJjXTuy3nOL1EF/O3P6xDsTfGjesNCC4fg6aYgs2IFv28AH51
LXo29Ye4Ttnxn6In0lJOYXGK72o1w8WsYJ72U234KSq6oCC273LQYqlNI8WdacIUM7QnucbNJ3nJ
gFHeULuBwLxpbcwWxqDfES7BrTGtLzh5fvcV+oYlq4Oh2KAP/YolPzPAe/cebVfJvtSeLXWRzAva
elEJzs0GBIBIK/SPB60EpBAGgEj2zIfLItPElDpR5oUrrfbL6MBQhu2lwf4hMWO8AE6qcfs5XWOR
adDJF8Rs5Y2kS2T7T6o6p6Asow3qDuKGlNN9OzTyNxy6mp2v8XpeAE2lJc8u0yTlDk/+ky4PlIeP
Wh12whd5LaimuulHS4SkX5T2OvJm3MMSUb/GfF934Rao0esfXU9UJ24gieKrVp78bLPkQvKm12Ud
hX/+oPldN5+NTiYfIOaTu+9lXL8SHJMYOuBFqlxojJylX/dqkgYcihLMBNJruxUz+62UWAdRCFWe
25oJ0Mbopr4965jwd31LmpaKboxItmANrEkQIOSuyA4MXf5uT9EXr92J9HMiTZlROXYx6RyRUy/6
d5Y8g23bnMWWf6xPeGFVC0bBne5QHL3N3OXiiBUUbLp6a2HbzwxQWhoQ4VJ0tMyhXkDfscbld2zP
iKLMTabJ+1bz5/RH3pDqxknVIPWzI1xxom+wYZsAF2ut28am2bRxeXWXVBXnMyaCALPL1xZPDobE
yLdRWygN4OMMOh0y5gTkKFbK0kZ9s31MGkFYH9HA+91jCLhNNEh/YZlqgvqBrs9jfBqAVqS4vhPh
o9GDmbZCZ/JrMWpZt4HJ6e51Ml3frVAqJhH0yNvIFMPcLm0L/RW33UkLBWfqxlRQQTDvvHZ2+foQ
i7je8p05JCovMeHDboBkLBZ98RABB/sTb0iU5D0Kwj5pMS9wKNUx66tFGxeRtVpavx1m+r0n1dcS
ms+DgAK235NL2L/moonygG6cnAadRCXJ6o5Ehzbm4MJHAyvKHj6WwXEhVioM7Cog2dszgYochXSS
LiJtVapUP0EKNauC/HQ15knqUgnav0bn07sVnySIGsbwoNQvVQKxkJJg0+w1+0Rkgovc0RQHW3Zm
OkzSADquowpFbhN/4DlVEA85X7RMl66uUJoO195eXhvP3lfVmg8mRN0ts8CLKExWgylMq9lbrbVN
NHu3x2bacOruBdY6sRc6WJ0kdhPWHH2f+Zud1iBPCFUC0krU3WARp7tJfNNBQuWP1a5z960BAoEk
KFJnbm5mCQ0q/uo8pDnOKWeWh+rJxEeO3S9u5GwMJxkIsmsotxlOVE7rXOiXM0kQGQvyKq+CTtq9
MQ6h4NsV0sm1C8juot3tKf8m+7+Q+/YzG6Bt1D/DUpZ+jLV4PMXWej2VmrrOsDqXGrWH4b5U/Rh9
kmEmVn8Q8edt/mn0gvV0Q/xqj0ntooEtdLrR9uFMGHLeImBYlwfd7kDMHQsy5c4/mM3d9k795C3j
gP5WDeFwxc9iyOEAKUuo4baPVrNcCBPUfspcB/EzBme2Y9jYNr6eRA74M2r3v3lLlCxvVO4JVCVo
M1CXdPqubtDCWRnJ3OwYFZSVwQRweQ/NjYmpueFRUlVVre8hwqJv0yfC3TD2Sq3im1oj+G7hq3iD
utfDaXtTjjERUFVrBdP2hT9xepaJQDLYnGTEI8ApjvemPyq5kPfenQAi4AtD7SN/biPn0m7Ub7Io
3nHitOJ77uWOkC/oDs6W6MYONRdxuAsc01klCNjxQABaPGBM1eeEib+hPZb9wgAhyBRWnpK/WBpP
SHf8FV+w8pMQFj8U5jht6IcSkJczpbaFb3H2NvtLKkbLh9mLIQ2i1zlZKCnNTRsBQaGor0JXfLYg
BN3nWESiZnQYIySy2vL+eHo8bIguec6rmtnj4CfqH+wCztMzPGir5YnKUisBCRo7aOXMyYtfBRbC
g/hXNOD1S5HutOVEb3zfGLn/tbLY7DX2W6AJsaakEPxHTqY+o65iWqbdYbGpClxuFhFDhoPW7vLQ
/zNr+EH3e//bTSsBzs8IVPRcmjam4f9+ncMoCuA/QbBPUhLkT51ufvZ4lfUxtymMNYo7XWqHjKvY
YewpRDDFVKij9ZyoGFYcTvX2rHyO6Txath4Ac4Coam072XRm6xh6TdJlxJb3Fyfhvm9QtrP1W/rO
QhcsX2p0/YS9RjaBEK+omYrCC4kNVQAOp2BAZ+THCS34lWMcMgS4oOBwxreLzx9yktZbP5w31ZWx
NNE1NC0UslL4cAbhG5yZriYP/Lzq+vhB7vJCKQ/iaOKfBulLQmvyUpdO9rXjC3FigaZbXml0rnRk
UYrtCD4x+DiH9Q8bt2cuNmLz5jL3OQbPAbEwRA4j1mUGmvok8SikQ94/n+sA4sG8homzKF0QSAzH
cZA/+34V1suXLoF0aG2VmY7cJU6avhcW5fnN0iGtjRlN7ysgpAo/0BsVIymvYDLJEJRO+gmGvw7+
U19WBlS2L4UGB6mCjyccCf5amrEk1ROWLYOZOWnJ+hlpFmfW8D9IgLXNZlO90ryC9NV+U1/vMVeT
APUk1m0e9kkbZwge++/2LXXJpGQQRF3ZuIgO83RAEjHbG/+0yWRVPLyCAKqYX9KpvbMxCa6rwOVK
Lnkly92OIMH/ztFxjUhy5CmNnnKj0hEZFXVCEgbzyZdRVWEoeRz5TNL88yva69HbDXdI9OCoPld6
VjmE45jGEKwYlaLVb7Hr+JF201X9mgVWN1fmv3gqsIo/XoJpPuHQunPaPyOY2a2ZdhL9Q7hVTEPR
UZk7OkSJ1RlO+dDE3JLZMMVxk9srO4vGxIlOSfKmvu787sIku1JXXOYW5bjTa8I4uVjrOsGl6uLo
fhbOcpwrgFV4/Myx7ufF/17EBlcGljceVKxVd1ipZjPnu0qd1Z3avm2irK4+ATwf2lTVniQXgAjD
OSlc5c9KcjEZZ5SDROkjgBPszXbaLy3XX/iY19ePgu9RswgMUNhSFmdoi6qWtSEfhQDHEohLP4j5
O+nDmgu/kFc/rdIHTezQYlidgi09kSxRXQ5xqOYw/iIdifev9Xhv+bl8wsSNB9hrkzFJUddR9miA
h+AgEgF+pZqnIcfaddR9kMgHellIXh+IfE8ejPyZkbQmAZ/F/WZOvTwr4VFv4v9O7d7Zn0xXG46O
UM9MVfmFFsW6mk23pkEiHMoodqaSARboGXJroUBsAROLpsUc1HPFUM30Sx2DKPOAiCV4Pq4eTNgj
LoWAlOD6c+C8+alnrTreL/xsTkjBw/iOelaSq3VO71M0vWqqT84LzlcHmSSFtdTji15hG/ISIXJo
weHfV8X1CqbLbgJZbHSN2Z2poA4hN/r3LD4DEXtEjvOK9l4EhUFFdaOP4r/+foRTZm2K/XZjGG61
+KvZerTgroo7lB8+3X9F60KcebBkNUBSLHhEJSi7AC1LNYMzmVa4UAfXlCoMqaTOlGfUvcIN3tvi
ne3WFHU0MD1ShwLCJt2TuhXkuv+3sV229z9QcPRrn9bx2aVazA0f7lHxjSg0IQH1Gb8EPI8Oq1dW
Xl+3isvMAJFshLfpxL9ciaT+l7BoBtfcpu4eHlB69vCpbv+jjk6H+huh12txLcSJTbAx1E9YWRw+
qCwcjKdabIOlUFdrEA2nlBQ42mH+MmZH3MKkhmI7RLw3MjR/pwvBYZAv4udLmf+2C/0SHgtgMAhm
rE3NUaoPWGvu1L0GUxyDQsVyTqtqRFoH/Twvo2Ti3SHeQhy3tATCkKk2LTitSgcKQ+JaYK3M9I7D
LW+4PkONvG4BP5MxFKiCZkV05gCJaqhz2MLRdFnAR05zR568Tgq/z8w/LJnbIqdM7J+t7ee2pz3v
ZpKFW+C9YAyCZypr8ykQDWljDUb2nwJhTVtjfl45KEAW+P3r9fyKF7v0tYmB85vD+EvcahMcBC+w
7rs8rFSz+POp/bbyiSO6EBPgPYraIEjBx1N/+yaf7juwbbwVsEzH3aw6C90j6gJH7HEFwCAPF4O8
8tySQfkTMxPbgIyvTriBFN1+rKoccZuTCExIi9zbOZFzkccjPspAOc029xv/YkVoGZpBKNz66qSM
9tRBYpf4ambnzyV9V/CFA+YyAntPyxhXuRhYWLeaMQ6zZ4kSe7hqtXnXhRfAQJe3wQVCjeSdJggl
Hf3QEVz4O7FTK9M9KNsDsDA8xWfP//r6nvE6DypIumhUUxRLDK9xn8mMm6ft44fn34GLbi8FGuVR
9hOIczKfkcVCk1VjEBQ2y1LEun10y3Efsa6NP99q34bp246R1N2lGqPnK66Ag5fKFnbw9amyTp8K
D1R8mQv2APFELAgqGBPpqwK/0HO/MyOBD8iq1ND3X1V1+JMsr9YgLqEXAMQpVY5XVenRxGyXhVAU
2qhGoEaISCQJI/Y3aS5ANlzcV4d5UwlHJho4GeYPVPQEaYB89BsWc3jM0jsKPX69xLswjDtG/0R/
NF0a6o4UYiorDHV/C22xQITPZeDxQoVIsuLlsIRYlG8EKMTHLmbswIl3jK7lVkw8uP2Vr+mCT4Mc
A4zHuCR89U2ZfXDQ3xCS3EM5vagXd6D+1fsVJIhLGeRAW/uGbnNK3GSn9VwMufuFLcgkQ9N9lDN5
ABazQkXMiOJZfFPwuS+eXxGohpLKYAfg2OZhiTG4Of3tocNpH0yQXEPh1Xa1bWdm7g6w1bw/FHWS
nklOian60EZh9VcCT8jYV0SoQkPyh3MRPNpqaUV46o7JO+0+M6E6EyMfIepUW112nzgUgEeUMJfg
TdZ4+2UccELOYLXIyLzUEXBglNILcYW26aWcvKfvEpkbyprSpphXkSvksrim9l7qXio14Q6GA5uX
4dBKCbH30eveTmc/dQsfZ/b9magYiixZbql9g9M/RMKw5yhgM5iTOHB7Z1gZHlHF+nSnS3+C1Gni
Wr9n79pKmXjHnOzLR5abnbC9r1Bnhubj6ZGYY0tvkS1rIltEsvVWaAFndDfK0pevdUOcV3iU98vH
0jO4/Ritnc06VmDUEiU2NAAAHRpG9dT6+uRXGWLtaKApaYOxPbcjBw3g7ICcd8tSH5YcrCXGEHcS
WzmXpvoLweba7goX6IfE6wjVZ4Lx6V9ZP043F+fqxUHbdm0sMX5x8QI4Xv53Yob8V8ner1a30FVE
cOWm2ICcFGoyHF6CkjKJ1GlCx21Eqt/x5INNVjFTcfwn45yhSCcAiMskXkDZHBoKU9hbhi4EsHGZ
vDuOJAOEkg+P9pooCBe5sXwdkkukmPamvS5oTGmUiGXk7Jr1RPr6Xc1YSLE8ZTyqW9zp1+bzos0P
ru2O2bVGZpmL4/xgdXlaSfe23tghH8q58GnSGWj/37DeUjWlLw3ih9emnzwWcjVYWcdo7tRAwuff
hkzzmdEC4MI2Q17VRFAJ2ukQvGOVBwY0+Shg4yQRBCtML755Mbyx7sOH1mf1q6pkSu4iXxi5qTi2
TuEvZEfa0nAgyE2apcWiehGTBlILm38K8kaw19f3j2sPpAhxRiOb08xUmQlriW5Le+VUA9UaYvt0
qFfd+3GriRMwXjlv4VokwNlR/mzMaxYWrtBPqiSMn+iK3t5Lkk/HFGrN+7I76Hx2/3RmsnILExtE
Kt4MDv0ebU/n3mNFH2ccT7ov5/2fu/JcihC3Vtx59qvClmDE3LS9j0x4hscubJqSXFBLxsrdo/8T
MGQWiK4EIFCYuMsppuPyd+fgeaUhKX2cph7WH4BIvcChr29e/dQrnOwwyzOgwpRHdFXdaetq+d+K
gjeMtzOIyBFa0AUhT3ZXh76/CzOgpWu1FrR+srgeiaN1u9Jt73KgSP/IjrevRJHciSncB+N66jDA
inyWgKouqPZ+D0DUDK6DCsoaLWJzYrz3d10h9swlWpVM5WkwDqObHuRrezes6ybh+wn6eNw6rxr4
lsKqKhU5x2qiyVvvJnKUBIlTDzruEiHJjyBANIlEJeR5QQCPvLkIXADa8cXuJCZiY3opPn+HK2IW
UQAxmNBCOHJ3FKijblYbMpPRqXGzla1MwRDK6NC+j7nF6Az/10ez7xwm8/T46okvC6IZAffPQf3o
heIoOV9Gk6E/jYbG6vBn9XBLbO1Slefc8St2Z/6uZCyRjccOoVo5ioC5TdVqjSpUTlHdQm4BmN5q
80w2G5Fm8enmrVz4E9nF37EjupvnhkgGn2TCzDR9hAw8NQAOrjISGWkJcUUXUF7cpQp1rD97Ma1t
xg2LsLDXY8qfxeo9t6nhSYE/iyqPL6LcmwyJMZAEWEY+q1NeMgQavwuIf7ObgLOO8FyeD+A3Uj2X
pbYFOsJq756GsShsAqUqp1z4cBI3xmfH7OaHRkeFuqg3oqYsu4rMBTJ3As9gHKidlVFTdUugggqv
0ApvwiBi1vUbtv19/xQWiQvDGdADxr4xaZgKw7pRSR47l+H+gG09Nrl2dDjq98FNjF2dJjLDsbbO
M9CK4ZhhyIyxwV85g2CvDKa/5H7JVxfMfxvK9LdSsAM5ejFIe7rG3iVolDDo3HgP5/ONiDxtpQmG
x2agK9IUCmGwF2yGlSPWy3br5Vf5phoxzdxcFHq//VLaKQsFloggK1yQAySZM6cQg2MF9kkCjG10
2lyudkLIvHq7fjvwyAeWNr5J+I0ZbRiMwgOtm54y6bdzCR6Hq4JrjB9vtgrWzmSG4NBJI7Ey6q8H
X+WSQq8mDhl9jicKjsJm/x0EC6i6z4TsvHVzR3ZyZIvdSVnJSdk4PBn3+RGKtb/Bl/TRXxV7houX
x4X2X0/gTHYWrtEiToFupE9xeYheBJOTHgGnD+skGLgq35bdoF6Zp6A7xF3JYULNhPrblFRv/cNU
QcmPoCQm1JswP8g8KT/bA9XfFxPb0fa4R/FedjSf4E9yLCTm1hFGwcfIl4WnfRUhxc7UgdpWFMEt
LLK2wmKa1BQzeNC5Cp17BpjwgTOjzJyfSBOfNQ6QE9anE7cdTp+ql0cT+wM3SGqhkIxOhJEo7RCe
XN26xiYaTUfCq/WarHdUm7wlV88WeJU+Fl5j4F6sZJPIMZAFdrILMMFnA3gaCfthaxTRsNEJaZuc
NRb+UTY999Qw2Ixw8BiCb43hJW52/OsWoKj6LiUyzZxiE4hxF3PdQtFRU8rc866Gt3+4iC3if3Ll
4QuOEh3NxOcC6PhcslPZdJcD8h4giKWFzqsh2KkUC8is7oMqzVxrzPrRjr5nRvbe+6g5N7XMjX1/
CEa6r7jDqsv+HqCadmEZ/Vjz2mWgOruxpOAtLJF8CyKjWEfXzttXRr2jXlBpQaeyQmriKu+SEguy
9fiQsHhNsCrzODDCPlKwiSi0HUMsF5ULyT3ZupWj/bD+xculYAwLsJ98sQSYRfgETEZkVs1sGtqf
rHQ65k6FupJqHpwSnLAuZFVpdlW5cVVHV9jCIsTGin9Qvnyu26He5gHhCH//GUr5tfr4Qs0D5sHr
O69ozlULtB47OmPuQnPK+4HqsxGm0O0DAdb0kzOQ9zCzUdNscrfnwqk3+vsfHIzNwp75nFBLxiAn
HLOM+9v4ZyXXVUVM8kzf1T1W7ISw3eBHeUqJt00scJVbDLYlNZDJ9Win0EhGatohXD07QKp12t2l
4B+6YFyhwGCTR1YInQGkjCwoRSBsDudCf08Hcqn75A3d2oCrqbbE07DAkS6qdVHV0c6KHNayxOJO
tQ4UMvdssmWaCOOXD3Pb38rkfdfm6dDBQdDOfXK+ac0EeHr8HhDcezHOLKUqq9DodonLKX9pwge6
QZSuj85HK/iPCAEUTMBtSRp27uyPBa/0RZ/nYTcgKhBL97loQ04eajX51XBQMt2SpK1w2wFO8ggR
PNWin9u/sadVc7CfE21lzBlBQLaVz749qBcUDQIphd96LkbzmJcrik+htBrWjquIF0aUIffGw70q
duOge09M8fEagPiuW0wSCL+e6L00yBpi6/bvibwklE9OyPHBIozV+jJFuyC0jLTQD1LYr3oINFC3
SrX5XnvLSnZfrM0Y5IL9jqMHj3KT7BtP1eiDctXDLItQpuM3woGT1SbD+sNnEJ6PVlnzgxPh00Xj
UzbnPKcG2IUjyD/vElQTJp5Nvyn/9W/fBFn3AbpUIGTBAvNqynth0VtMgkubfjXLd4iLmiYA36a9
K4BoWaOw/M2d96O3PJarbh4l/1CIfSb5dGRYZxX/a945i7+efVJT5/l+bN2qde0lrvKRT/lqJvt3
xP3gjPEDyI1HJtsi4zPz+EMcELlpV9gqknTXW9Vzq/UWPLELcBIplKaOwGNZgS5yg3MR/cM6rQgn
/1xMFBlyrkIhtmKg5Gvl8+LHnhiQMPsEoT/7Gm8IoDeI1a77XYR4VDxxBpALQSr8XdRBBLS/+XxJ
J64EPOqMiKskvemrrFvzmm03wnrieCE2kpv86Umx1LqWRvCZhp2YWsRBFB5VuJRThzIQHCbR6tsn
okKOUiI4oZy1R++0b69hSRH2AzO+iOmQkf6sEb6yMlw9FBgPANo+IQM9b5MbYwtNeaDQ3rYgU4Ud
3i7G+q7Gqk+FZP9Ag0PRoIYNSLFKI2NEEVzci7cR9v7b+aT/KQ6sd6Z+T+Gem4j1BQ76LHEQwewQ
oVZdKe07Qr1YS6zhRMANiLeECeSnrEj28y4es60zTuaJBlNc7/5aLUrsOPVxBbkZqvO3e7OHdB+R
6cUtpDypje10k8S0uFBHgRJDDiwpkhMpSeWGFjPDuFccFVJ6DJauf4F6xl4K5o8w7iENGo05p6Jm
VfcDmH1Xg7ZMprsZlVGlS+1X1qqMjiTziMT3m+8ubaw0x6KnSwHBPQN3qcSHTYRJeLZaqsdqS/WM
7e1h+mzhUa2Nd35/ggeo3Du3bj/JKX3TPgXZCzSh2OEVOyY1tO0OaJPkMNOLFKK1yUyiW8F0b3JT
qZ0Nf/j0Sgt75DnWbXkwJB/wjjUXZN4BNuaGy4VnI0PGycyYNhOGO08oqlGrh0bwmeLu/t5QDby/
wW4GOdrtykyq9Fjzv44sRk1THzVnuPL50mzs+R/uZNCK/sJGltALTJ0+sij0HIhuB1dfWOt5WnC+
T8cMeRKqpnaSy0lPUdlmJ9DhmV1KN1Q2HzOIqdsSXnjqpP7j+l59w7oR7xFRMJV4QyA4WgNe9BqJ
eJQEKF1YQuRj+5OWtpOMcR9eDzvlk40OV5WbTh1BC0sSI/SPDrewUor+4FMrfJbEA0d6rIsH6K9a
d1rIE6zOLt0wUaJUQ8S/bM18xfLAQaVRRAYMMzlpXNlWoiVOTInM+2N2dgMzbhB8KDTLuwpbxt9I
uUpTIoNrd9HubnxEwLOIK4baS8+lI9IF0Tl7A6LjznGEUrWiF7K4tJcRqkR7F9+eUdIQeigIGTWq
vY0i1cWtoWdfj8FLUM808erJq47w3M90b4liNH5msGI/B09dB7IaRpJpU84qVArcAKWMjHxL7m1p
h2gOPIeXekBU2YhMwnHSLkB0c0C0W9zoiCk2e0dvomUbV8bX9upP+T6f+vcCOzB3uAq/LExBflML
0Mp/pEP8tN2VEVpq+xeX0ooLDm23jX4gc822L9XoaVsD/pYGSlG5I8wi13pOLOiibftbSbWD5HcX
NHpdrEE7IOk1B5WvACSm88L0JxAWAyPLtIqhprVZp6wXOvAsJiCr44FsG9BugD6MBdZpIbuHX478
36Qm485oPr/qja386R+kXHdWiIr/TUpOYik+qQuOgR9wxIR0uEnCkWycDj1Jm5e1JxU9b+471VxY
PdDDNeC0TP5zeErcMohmr5wziKlYBBgwXv5SfCFCdrYwjfGlkIHgpT2TeKQJ7WfZaKFKMIPUj/g6
Qim7/STg5fYG2iJ6Pf8F4bvUd5RkOGrUb273Iy6dYXsTrqVUcEhOGB+NIcB8Ppeist81Ja/EwiWe
SVgs1s9JN6GTKLGSx0bfvM5ChQpOmtX0FwmgU5bpHV0jD6JKuI4UdZXLTxPDn7KL7j4f7+ugj9wI
axHMcWAvY5SbIP2p1/YEZ9jqwsj/XARSThrrg2GSgG/VA/Au3eUxOnQxZGURmxJ4vOmN3ZYwl+a1
kEespafTwG6BEnGzA3+A2Y5i1PH4jAYtwkt5AuZhhVYIr7VAOvFwgOou85AHpUtL1IqhNO48y1uX
E1flJ8zZjRtRzX11PlaWxEb1ytlqKD+h90b+mIABQ2tJ5yGQrtYzhCzd0YD/wfzktiH3nGX+cV7F
6bj9lY8+XZ+288Ll4QE+OgEKHUh7UYNIUblWqSktRAthFsrQJFG6sy/pOmv5xsUBRQSFHKrumFtE
N9vZfhAYdTo4tNIjCUxK15O1xeS9nwJiQkg14Be9y0YUdt5E7QFuUBHrqBN0WrW4m5ykXdTvRVBy
wpZ4cszVbJ6IPSiFC3DbIc3s/L5Y1vNnweKdz5vhZbLy6+q7bRpLzKqvo8pgY0KH4Bv/adT0n7nQ
KY8Fs1PHqM3B6YEC0lww3x39VuwLXURFQpeXk/w2mrLBjTh04u3jK4l3HmUJ/343LC4Yo4J6ZMfU
eejg6jFThgOWNm6WqypoJWuBrkQv5RO/+maFBmUgcEBTT5Qh8AZBxQm2O2P98aaDnYhSPLcHA4m0
a6CMMkplMsmZk+B6MNO6yC4mPrYb/R4YbVb/rTSQLu36WqKan4WQwN8gcU+xL6dYCd2rRyk4mPpz
8+IEqcw1yfrciv8WWP0e5g22ux63kQw6Iib0ugq0cSzFEaAnZaUiSNLnquDWOGt5fIx/r9oRppCW
NPt5lN6X8kM6Lfmw5Lp721bL/lNrUNAFLoqMRTot+rRDBQ+TJocInhYqSZZRFN10qd/tYuDBxL1x
S8muTgLPI4po9OpsbwN/w2LZ8DMcKJUcFtIrcC3bCsdsbxHTst50tM1ruQDig6Psvhy0dFD6uRP3
Kxv+o9Jhts1red/T2zIAFzNDB0FWDvx5ohKpFYft9CQKzq51HrPO07pI91b9EWsOyJT82B6odByV
A8eKr+K0qMZr70WmOkb1UEO2mIe8ocmr1hloUfjcEsLfRTBwX2mo1uUNg+HPNqrWrmy1lfS8184T
z6462WRqAc9gJ+fNy6zj+1g4aG6l6a/GwkEM42hHP6Qb4BaXvLmtL7sHryvZvn5li0VFKppIXyAJ
Q3i75xH9Z5f1loE3PSLtQxA3L/ppkCQBBqMs32VbWDW4k5m6A0ZU2e6u06XBJiuohgVs7HWXKsvj
hjDK090XyNh9lAEMKSIsY9Zed3zGw2Fj6YkeOlWUxM9zLmhWw0nw33p1xAqnPt3e+yX7bNDRBY4F
pD7vfjN2SdAz3AB9V7NBI2qB65KySa250IHUDGuIZQRCgv82uHWo2o0/5kwndAsOqIrXu0B432Mw
nvFNfkv2zyTJmFu3bxtHUc5dbiuSURg/TIuwlVP5Ny5MkPtNWBgT6FEbz9RHdJUQt9ls5gC/71XC
qqT3vxeD8rSl+m4y05hVVotPoE3babZAkrzFBQbwTEnU6T9rkLZQJn4iCm+fLdcqPEMl/P62sBxY
2WPgcYPrGgb2Ua9IZwSuFVKyzpDktwBwk9rU5TDuwGIYB/3Wlrjoyyrcy1QfJCUjN88pl2g6368p
cmIksl2Mk9j2M4OeT2nzT5hPnqXob3J7qQRydanq4nTH2L6LCkyrA/llc2NjeWxhNyuJP4oIxVkx
qYhoEvC/FMFN30tJCoTKGQm3SXSbkOTbk78mjhQDBH6Rg92aLxv9th957G5nG0gJ7qS14AW3VsTG
4+o1AAqTynfBpdTbVRkVcAY00wyBaiHPYa/PmKgitGAl622zXt83BWtVxdfEDqJgWCiio1KcmBBQ
OmUOIuK9tnQkSZNNxblsivWMTCcfz3BMZgjaVNjTQWyehYfAXB7ei++aCIhj9e6/aX2Ns32u9Txu
iWgufvlx/QcaU9Kah3Q8KZvvJ5qBUum+UMc17C1X8FWJ5XX2E5Z9QqIqZ5GBYdSiwa+nqSlnZPXr
rnrTmUS5YWMbF7VoUfdhRikaGIcIaNvQ/bNTXk8j8LQoSzkN1s299/DU+ACPqpW5mwcTy38Zr6h/
sGEPacnvObDBJVERJUUyZy8YPeVk6Qvo3iU8SRUbc1jpwWUmFMTN3GxDNA0ESbkJHmeBprna9TWS
vJ6Y+1qsX9rQ0ZTMV3rRR2pRL9Jyk5qg3RZUHynUN/12k6ONqLiJQMGc+7kklPXSyl0V6GoMPsRj
l6uKs6tZ6y46gU+3R88X6sqVgwLXilBwXJrnrMVFvvCwacT3paEp4aFV7uBDbvOZdzMIKXBs/bur
66wryEJe1lN1KKcSjEq/jvdoWdmOEBHoN/3AmOQ8fHatuDXt71RL2WXU2ZkdmGaXDYJ/jiA3sBUI
y7fF1aBLCDyJv7UYJPtLouuaRmrAvf9AezTOpuvgvNlVdBdFC1JtihvhhhdtWHcYhzt+SFwnV9gm
mZOx8rol4z0teIZ+3MC0BLRRRGaqkNYPG0YA4Fv29JSzoa3QJL+N0xlo1I6qGS+zJd8LIqKMZe/O
YHX4LAIrkvZsmd4vjKPR5q/Q3HcVXWs3cvyCJD9CHfQmgFifuI/xTOBqSndsTNDgcZVxCm8d4eP9
PzRJ5OCUY53Fiz4t7jFsdI5It0ahLrK6EHDEOhUKIU8NMTG7rsnEKkEKtxVJebzDsloVsRVuY3Xt
r9MYh04cFTvQVmEYuTK2KZBuPYsI0F+tw0lA6tqSa1UssLfVLZyz5QCd+AT18yP8pqTLx4lwUmIr
Io57NwkifXezY9O9kdUg+C5rCERosZnev++6QO11GIrwHWOYaFzcWSD//LiJGVbiV4W8yYsGLSM6
oEixY9YRuIsDKOkX9jNGClEc2rOMQESuO4mHnfjDwgHhtqvXX+GymcTLpMAWW6ViDbuTyZ5uOD09
Dzp67IubXUwbiOSMqsKX6yer7x+tSIy16Fg4FPELpXQhwSax+qq0MMxTEXYPkPSGw3ZII3UBVZIP
8wE9iMoh3nKvA7mnVh/o48p+mOidXVPdyeYB0bSUHBHYwYJWuTS7CFmdBYNhlZAkN1ni7Ur0k3+C
8Xtb6jqVhaoSIg4JMyYHsgsKKNDm51wcKuD3L4Hh7WfSX6i0DZpx31m61LlmTdunN+Pz5rpXI53B
0ljatJdqyHEDTA8YKGmJupr5RwfDtISkASh5br+NHB+1UgD6jcJEYP4P0tahlYPWOjgGxMXOEdMi
bJD9bxEERr00YeYhzH1FrA6vCs1b9On9c4WlbKDyjSqcdv+bcIOZCI0Bk7tssXbIozoS3mI0hssV
Gu2DixCCwHpNHtkVLWDJ3uPnpQbmCYcUT47QCOcuLtFsyE4eXZsWdVnkQJ33+t3N23JOkEKDt8ah
U22aZ38KgaveOO7EsZRTiJp+3Dtm8xcc67C9sflTPLjn8GP9qZKVWYPLzv3QrtcmcB0j8v2XjyvB
+XxXrKB7laNEkEQ+h7smDSIxPhHAGBA/dHlBs0e9qKcImHBUt0V+aLlvIM0vj0rT7vQ02xaOrqsM
aPCou4QIYPy/xwbPJSrFosviBDVL/73JhcPxemWk4fxfRA0CmDsnUFy3MCFJOlGbLG60NSJ5ZikC
ikupH+nI17+lyBbuKmlS+nkK0T2Q0a8mm5iHbDYU6z21GGeOQWEV4ERGjzU4yJt1fmvmZWgZ2L1L
X7pFe+/Fqt0UqS8YXq+hTPKXGLWU4Z8ggXNw+Pe2e2q96FG5Zr4VMqoPlFMDqcqk5qTH9anZaykj
/mI+y7OzOSZa5CJLGqZy+s0BX+v/IOgW4sJviuLeiCR0o+o9738qFE9rB+xdPT41sGNET9nPkzSQ
5QEGV+FiFTFEYFjj5/D1W/JmY4w8bjQOSmNa/cO2qM/B4CMaPL9akHp/nFqfmuqlLnoPLBNlStYa
loqSAV5hDvxSOElXRKakpC590Tv1R6b28rXqjc4x3aa1VFn4P260ETjtBXUUjCs4RdSh6wkOrWHi
GQABeE+we51ppTHzkxN5aJb068+1DtPx2OM2EQkPqUAlzqp+lTuJkc2sOIgANCAjKX0NkClFsBcI
IgVKABaS84BiDDJ/jY8HnWTIQQcK/At+8m6GmGjEQ7wGzcMyTNf7LEAzLVNs7xjnYdSYPUc8hyW2
6hVXHBAF38sCuvBqX10oQnuPEqaKHvCLFRPsRGYno/T3xiBWTDNdoRyHVj+06WlXc3pHafSi2R9D
DQlxR6SlGM4eF/ra9DXiwKLprK4cWlahA2czALps+KtnVTmH/rvppxgENTQq3t9TuHHzYks67LB7
daZXKdW/atgF1xKi2YW/sqyv6yAodkWhvtTxW6sjTFbO0HXtaKoqok/VWqIT/xmKvJncgy1brcSm
QWhTYe6Q81y62J1u0BKP8Lzh6OKScVQ2l6tROxueBerELn04fTFQh/W3yCGRKny+hfIkmYTa6XkR
+dG7kNvpDMN8m5pc0N48k6twEAGHwVfOklg/StbZ91wAubXbYpuNhrs+V7CjpDQYxdThASF9kLpK
or+OX9Ien82AWAwFZh2SHZc0EzDafk7ftS0r9cU7/gnn56fpwQBpdUb2GikDoFAICpbPa/KZ3Tec
us+nCXT2SwbcdbJSRmmgMgHjf2Oz9SiGluHaPYqbJDulXuPd2RldSvyygqOEskfcEa3WiquwiqUp
9teObdC+jdZxQbUNybx+u25OuLr2BTi9DRtzyzv5JkIbT+3egIe7SKSTy5bVdqtJB1cJ3pcn95D1
CfW3eL9cCx6+awVnXWMGkr09xq56gSkadqQdSyq5yYeGqPfQFUxZ2TAhQDlj5A4xZFpKiWdI0zPE
k6lRPqjmmmFaH8j2DAWkL8xvip25EzGLtcm/jIkaWzfHI3JIEg+3gozRO1JWIQygJ0lywSWHxemE
3xnSeN3+4n3Wma8rc7rh+spUerm9T1OxgdDNyBBBqFmNbe5jZW8OyCKYf84s+l1gj5qWiFuHp/tI
UK6y5dCI8DYzcbfHOBcamYRIjoXu7xL5IhbqcnQnXYT4Qgca62wU4swNV8nUrQzwl5hBHeqgcawi
o9FFWkUcZTrjY1A1XcTGW2VU2S9bC1AskkWidnIFC4kvWDJLcCnaNCIh67ecOZH/w4EsXKWMpUa/
kFjteY1g2Wk9KPTa84LglGcHO66GGcbp5M+l44AcpCAHrFm3mcYWD9rkIvFxPRaEzGdn0ry6okeX
n+Jarw+vJK7psJmQe148O0YIOshYLoHznUiak4ibX+XM8wJwLkAE6hC6JQTPQk38k/2RINnvU1UI
NQVew1Nr0kifBfUnV/uMkKIDhNzUkgu6jkVrKyu7JP4HuVTPD2wRBpA2eOD9+YM04pDdvVJIlbl4
6mfNYiMKtoOliRN6bkhqcP97grRDK0fNr00GH1ciTos/btUtxocKHUs2BLohRF1eO68jR/dY1FKU
Lpu9dt7GlTR09F3R+pxYGLJfeB2E2VG71oFwGz/Y+RRWgShOr9f0muP8OoDqPyi1ZK3N9tAEd1BZ
FlbsH6M4DjvW2sJc8ayE8h9Wp7RMzhz/Z0pFIAzk1i77Ju1mZSJTUu9RxLRpAto0uaSsfHlAQG6q
NL0ehl8bY/xoCkU9x99MMLkXR4pSzwPL0j0XK6VJDm8rmV/BBRfyB1qvDGy7l62bINtjFrz67Lmw
troeDL+GYrWznyN+daeVVVvVesPtsyE6Wl52h8ZQ856r7kcjQyzPTsMSg06IJlQQ6DwFnXzJUapy
kswFti46OB0lhXRTOB1BUxX3CjTIkl/8aDPLXWUKs3+Bjw70K56uE9rhRhmPhkfVhhlr2QlPHyUk
jHE2wVFJv/RVmsVwfn06YF87PjDzrbXIhlaRtH9OEolmr2e3GxTZI1WVkVK5MExQtPQu/kfxyYX/
H3w4OgLIv0M04LYBW9RP/xoV5q5RVW14QVgg06r0CvmLRZfm5LeDBeb+N1KVg3KCI0YVlOM5NMtE
pNVBJvVwhcnU50xpP1titVvMw4eeQwpyiZ/uBulpGeXXOKJiVki31hXFuhcBFHMTG9VWt/emAb0D
7Ch2cuOyZObWjIZeI7S0j/vhrlHSuMMrZ9WJGT5sHSypO7+M/U1BpU4bumxxDcQHbA9NmJZEF/JB
z/IRFOKw9khxpyNbiHVU6wDSSeCC/lCjiZqf/QcrHMx+ltNQC4Cek+tFLt+dn6RZUHNrcZTiPGRY
ReyrEBYYixyvfNHfq9CD02HyDBZt06TawDiRDPvJDCddcajKyfOfZaVmZQ7RDcJOm/wYG/PlxklC
ahzi5slF2ZZrRobJzO2RcWWbbEWsHZONt9auM3e3FoyyP9vlPJsFxU/H5L0A8iMrEJ7YVPVX+RPe
tr8DcgXqnbpcSg0+s1o7JyWaw0EnRtbMJSRrj9SM4JwW8MavZKAWY6fK/xLzSTVLXd+Wx459QLV1
gOqaJHCIKQanxrbNW1bjXap1YLEn8cHGPMLTolqLKnRvusrDEsh+vqJ3aFJh36WlB1qvmGUNmH+J
PaXHveIo4yYMLNRLrWWou2w1ypn0EHjeX3WWiLt9dQevsuk92Z+HCqPeMy6uVf8JdxFGH7wRtVq7
Emu2swG6IOupF/TmrlAe6xV8m8u4D+q2ek173YdrSq3VA90mXic9uZRCrlanT9z898HwHtxv2bW2
WTrMHsW3EhZmJ0dcR8uxfFKs5k57sDDFSkbcOrSp4yVrzosoptRPQ4F/RIu4A5/nT1bfQX5EFfrD
XmPj/YQf89rabwaNE7ZG9D7/sNIj8OYuhLrKIY/S7aezHpXMIKaVftPlEY5Y73eOvaBcNdN7Y951
niRaNw+Mk3U8x1mrpK1MGXoffZdMxQLzw/NEDm9FmFibXwgPtdo+msc9cN9NPLJJCT38batHk2Sx
Xbe9Thmft4jHnaIDoZkjJnyb3258n1eJ7lviaMhUfdN9oMu3cJ9V8SjOz7QHo6qWOeA1pWKMLjSw
BG8dOpPN6djOx6mDOfSYRuILwJH7danbYiZnYDe86fm+9UC8k9VNNqvF/PQH3ItHYnZx5hxX9tWi
MT2B4Pau8bchoztBIHGw8kdYil2iMRwoH6iLUifnTXtyJrou40730Kc4GE11PBnBCL1VK+skGlvM
xJhF1m0d7KkoTxKLBJ/oKuSjgLKFUMVYhqXEtBsPNk9lu5pAIsMVWU3FTghxcK+ElnEFZWnvZBeQ
KVu4K4m6eatKHZgF0C15QfQv7kYUz9qEVQaC1WahQaSXv0J7vf0qceGY8go5HbAe/ND3eiEF63ok
6CWw4X6D1B58/YUWyStLr+Ph2d9Tt0BHsZmiOhQtWuNYx46cEKyCZWSM1X/rR59cOGEKJ1S6Djl9
lw7Jt0rTXeRL1fg2p9+2aGphFqxJ0gzhw0dMCsEurmi0D/MM2l2teAnBREg1LIz12E+dhuREy8Qy
wX2WsEG23yBfcMdEKMKVOBnExX4JcKRpU/9T/0JWWU4xilWQCWFXvW24ha74rGes/q//xKOjY2hs
C0s9e5gc1d9k1F+wMbFjM9HNmNxall3k4s/XYIz2irKWvONIL1Gv8MkYJcjGqQmLZlxj9kOlkcmk
jv1a55f9gwZQIDUvx9Eyc73dokgkzsCNV9i0qhdpiXdM7E+CO1ETR+l5KaUGsSnhbPC5k+uQTXb5
Zb7GZAaYrLVBOcW4Euign2p5tMOehYBTIDEyT/kQeqQFvrgiQuiLZzUle3Y69JRBHgOZ/uD3ayj+
tTpnbjPOkGN+y2QOkuJtx7fFdMcz1A0mavU2FxKpaX/LrtXbFT7+aG0WnywZRzH2Gp1QN3Sa9BNv
ELUmzZ4rnsHStZ+1a+jyVZgEokcFayDAXSplp3Z9gKP03xK7V9++9bsyLedCwH5LX1s8Si48OVTB
gFEM9+XQ9DEO68nhcoaiQmACfzhwdMgGmMK9mRI/lCmA3H8sY3ment7DxR14/qsTX6fVHwwYCQRB
OhOT1lY4cX+0tGmRXMJHJ2PTbMjsIWdvr0gOgsJLsC44bwBE3ic6XyBugTGq3I6ek/PyTpSAOrTE
r3EXKday6UW1ANFolMX3d9COCMkKRL5D4Zc6fPKf2AfMEI1cYdH8JHCKiuSeztSROopiKnZHZFld
sMxC452cBrQ6d/jVImCWI+sCKYzp7inO2OHS3fySnWqRVSHkQvYo1ARwjELDetp/oOsldB2JaThl
Jivl3j7eB334hB/x2y98Pj6eZD2MSkkIleY60/J2FuyIkL7lqY4K1UZZNhgLJ6yPMX1G9pITNOwC
ysGkAsxtUka9N5DdzonxTdiQ+6dLkBYl1DWBSdnOuPukRbTQs6EU3wqd4G0hGVFOzh4tg64B+xut
s/yP7kvEzgmb+FPfeFOLo+YGQGKy6hiObpB/PZebOJLk53/pXXwqQKa5ZQM0HJbnaGAz6Caan/+j
XTRtVovVjmx9Hvg7kED8LaVKcCHwSwyqsDrIjSKMdKTagnGVRTAmmCv3CELGZl91OKLmFcH/aRJY
lsK+DID7MFBmjT78E7Ss0cB4Vnv2hsNbq5yDhZkVkN7lrbnFx8F/5Iw7EogzYpyTzvexF+vKSn4b
0xtUjPJn+/duV9ThfiaeU/hWZTjOZRwhJbEWMVcBYl9M0jNUNzygWvrzqutLsuIwdJZv0GPD5QeS
aq8W1NhrwNAVq3aH5PHqPGauNd6AQ7qt6w/4fbtrnzBYGqJ8DGV+3G4nCxMU52RKWDbo91xObmTU
J+HCslRE2fTak2FEMl2TgXeHMJvmR2zn5u7Jy+hyyfEVjDknq8i7MARwpPJJHVyN/k50KuzOOcgO
gT0lAKMIcl76wSQRPg5fcfOU02ZGcD9q40aSWwdkQtJHTJ0cJYS6LbpjAqL08pxeR6dZ9z7iz6Yg
fMo/8DtHUPGKmBtLsaW6pB3SZQigzH2bgAFZLgQvm1Ra887T5lGJc8+cPhql6AoYLv88U823w9ON
8807Q4MdlTon3TBOWYj9vMVsWLbTAPadibdWAXg5GWJoWDWpgdDmlaKzZDX/si2EltxbwmMMQ+A9
dAp7MDNNzhiGh9FNGpcYNKT7OiBWJLrmhSTJw7aIKALOfO/S/N7QSHd1ojqWqDe/IbNWnXAJpov8
UoyMWVx9kYapASaxI9/U6Vezg9YTxRkPp/KlI2Fys4K/GGxX9la0MsjkkQXnjAXoKJ4TvxGu3kRI
juuoOEVZ7FbXir0izM2s3Ej3vac77b12k9rBzw1cGZItdKrfaweuvig98HKNfhAD76jyWv0GGNEU
7rV5UAieCnnihkVehg1r4tuTMwA5exN96JAgw2f/JZCCIRR0cwssX/yf2MTyZYROnL1MO8r7/eEG
k5dN+uMCr86XHf+kPUMPMv5CN5DXLumHnG761AtCEf8XrE6FbYvKWY92l5gK+SmG/GvXxxb9PETb
OyH3tVjCWhfZ6ZfRRPXpL11i0cNtfQ1K7CXksBx23lwvU6nlby13moyFUf+2wKIyf6hhlrPv349u
ry7gX6yfF9F7UtzgjLC5tcdH07lKTckB+v3VOWsT8jsjnr7AweOOdzi+JV1Kh6LSKGtqkNym0SS6
JU2ojIbn+QjdlIWbuV4MYb2fVskrdR6cZWNoMyF4IKwTSUn7U89bYreAjcPBtDjSTrDRjy8wC1O1
ZKmLNDr+qdSkj/zYEaYEroYic3CgJdIxO8GBrHNjRdSdMOLYw/heBUz3QhkLY96mIKOKt/Lt+vbC
t0yDkZc23wLMeblHoL0pE2pBRR3rC0SHtJIwkzAqmA8r0QfvRlpsISR2fh7YOn2XTQ5vceqFmLFd
EdL26PJIRi1SYBlGUhwWPM3TaESoOxwRRdP4PPRHgw7hYMfom7AF/RNWDpO2ZDrfyri0lxSzp4U7
1sO8PJwCtNrbLixXJWzJUCJEfTeJA7/M1f0Z1vuCaR9g5L6r8xsvCFrzRdtVp0iF6XwHLwrDHKgJ
S+RMCChibk63lXADy0XaFzEgWo3cXu2wgidKVxCSpGeuEuCKHrg07S3J6I9Oe1LZvv52d54vC8iv
RSgvRTVMNQ2LAe04DyVLa9/6hIyJsQKL0iViRg0i0Sp+Tq7JcuKyLczi6y7LCD19wDPQCoBbonfn
PWCMWUHJ6g6a7oa/Fl3idPD9eLyenfunIaFDHJNBZ77hLJltO+I1DP6597f4F0DvVSypNw6c4pfv
4vBZIFJxTFAi4kgaO/zfTrbe1z4E+mvLIj0sTNUFVb8nplIyVMZmjD7Xj/SZBQBaKcmD1fCHRQ2d
FXwb7XRNVBcPN/IDcNNDbG2VcO2V/LLD/OLDmc3QKqvARbSeRGsZJNJK/l1nTvGZnggOIU3V6zAj
CSX2PnoCsvMw2kptgjPee8gNbEG0mRSTsSq8gccq/eEd/L3N4zTnieXi8Opr0vXFUlwLWlsnNWkm
bzltNnM1X/dnqhhvRu9Xef9oOLslNgXVaEcFQQ4P+cnXlr3DZ1gVtrbSJqnP06WtGt86rRvJP9nJ
6Hj96gSX/zSGLDEhQTWSi9G1fr/crBou5QzmWmzy6TPvnhQFKImEWAiflpyY4TRE/BDq4XsObkUf
yjUeIxkJ32DiIeKNHP78MfwkaCYBblX7X4e4DfIPoqa5gZAbQUXRPky2kDwMWxLOGOUQ8NTpE4tC
s3uXEoLMOKDxv2maJANTLskiPoghvnG3V6kU9krhYbw21Du7MUYRv/s75OB7Soi6oI9cywqa0/IL
x0A7ZdH+sRc2ht4fjLn62qTWOGIHjrIizwgkrhxB4TWl9L7i70Tbd8WrzqLWtxAX45FbHkXWCDwc
5MEUXii+IYxVPUPOaxYFp07w/N1PWgTv2a/sp/cozNjueMQAFTNJUaJlQto1raw5XcsN/VaujsNO
RQUs7W+oe4nNLFeo7q0V140rKYGZ5IZW5NAOHFE8WAKzHtVf9ffKlBOtstixBc+Qax6X2SlPC1nB
BYAQ8Fz9VK5wzx9f27A0RBHhpUGKxmhwkHovRBERilEo7Q1iOOJvBPZhRZ4NyXijl0Zr+04cMOXy
4un79BhgSsXetmy8NiVtI0PyhSZhyCIIGUcj2tUClcHU5DewDWWD7bZpW6+SJsW4KafWFirTRhPU
t1+cCFN+Po710pSWjTb9gIKqfDbMy2Z/DD2aoHaWRiUJznXNJsx3Sdy9ImKoEdIdmIzS0jgCbdcx
dCMhmzAHSSEWMHy3JcMPOwICUa8b4kpqCfkcjeOnzzfrvOSn+D1adAOYjL5VTm5Mc+d8njDgZ9OG
Q9yB5o48sF+6WHyWsQKgW7TT1Z9WIJdwTa0zXQ8ZqgYs/PXkqB6YjHTholGJxX0M1cQNabQdvDgm
MjNu7d1gtzyT3dL26wy3qDs+VE3/8hTOCi5IKxXbkY9hrlg3ktPsYx+sttfG48qYltUD0M/11h7I
Vpy9ls9SHCojugVDPYAUBxUfSjfo/UivXhwHeH3AFyrgRVveY7PWujoXumSspKHEPaC0XiwZIHWj
s5f/YyvnrDgTlWTGEOoXnIq1Q7Tg7KWUybTRS6ryF8aqnQWRKjQVvuxhJtm+Vcu3j186L0wDXMhY
u9QXcro+iQfWWBD0+t1bhemhfIJHgdghX10PjnQRnxq64ucCaj1P+rgn1f+18Mt+eDNltaQSfp4k
bqBWB7iOchHFAh+p9jNTO412K+s04x2mk6ohSK06ARx6kXRQ2lBkc1rQ7C8UiuXA5/+mx6gg9K06
mrkRTf90cCJU0h+gHYjRvuiHm45bOEpj/b3ALR2mCI1Z+I8AojB1o+wJHZDC4dr/u+/JQB/fNwhN
aPsGzcC3jkJrjmjJ9xLZNdq7a5j420+D9bZmxuvI3nYypu61SUYHs6A8pMl06gYZNDxdjNCurWIG
tFK7mgV2npierTivr0lEtEQPle0junab6y6ikGSUeNNSRAdSEKjmlrO9Ovdksa5Qijw4tOM2qJho
WeC5Kl3tf8kXyUXZ0CUmmJkmTwqzMs3eR7w9pedaS8S1eaf/9GLmlnnKnLL6CpbScHxnlZTuibcL
GMPRAlfGJdPxUps2zxR9QgNGRB9q7x56r5UuTdTtO365X2yPL4GBswF1n4f92RZh6HXH2QDOrsEk
BjzyQhiKVMkvS8BAJBpxOcHatNXPJS7i38GPsXenchrXAn/ZKdv7pYP15IGZDs7ZOjMcj7f3u3AQ
NCIK45/4LxciXOWjrEeh1yFL9Xngey4OvLT9+RFR5a4+k61cr4qGMj35hb0s5snGhCYdoToC9hg6
9KHiq5GBb8kPUm/flqA+Poajqk30+88O9m6LkqDQl6On32FhRqj/uegw7eEUPdj42sXT4TE6x2l8
kHRSpervLjhwV1All/WkZdq7VeImnYCrdhi22AfqVin4J7Cy8Ja51hCP+vhu1aFLuQqNuSZv/RC7
6GBFvX9o7I1btpp0tnlSEuBB4RG2iSSiELSvDvYwpjYIsR7Wfuxb6t+eUMHc8LcYxirsIESydhAs
hJWZxFZDOC5JUMZFXMgCLWt7UuQ/LlnuqvYLDwYGIVa8sG5O3i5BA2TcvJNO3r3n80UgTLE8box0
oOHaRl06zwzyNmqy7tGTkGO+FOYdgh/hj/MOUHV5A8bQSx7Dx4yKlwqAlzEdzA2/JG+NFU4QR4cY
lWc3rSwdUecmvtiNwqYhADKavLnYFhhjrv8xsMtOEtEjvGnvby8U+8wwCd7vMYLb1qKJDdls3knb
k+6tr40EwHpEpF/EhWSOe8pGgUpe+JV5ZDNhx2lQVqfObMaOcfTt4cciO5jKpXSzbGLXo5fH1C9R
+l/p/oGTirrM1jImI+MAqTO9RBkt2zRbV28JfP98BvpPGfWEHUIgNwatvlY+z3UXTd6HfI5zDmxW
HWu0o3h1khLffq5jk3f+R7NARN26bObwwnO3h2C6pFaMrGVFCVj8N9fMrp47Gr2JsTCssKNdS3hM
0HoJnzUono4ZbktFRY3Qud3dxOv0+7BIF9zgpN3KniqLgGKXYoMV05xd9tehe5gg60fQHO0Gwumg
l5ykXmQCD7Nzc5TY+HJxPoG1oavXzXZbbmbkdS6CFBCd6vT/ByEp404F/nRa17KZjw5z4jl0X0Jf
mcEO2/3BPCe/E+MRaXCQtarXyx8esfbQT8tfoMbHxAM5LacdcknyVrQAmX6338Voq52ZURlu4uEM
aznyxB08rhSe8zNVlLXVcaCSPCbGOiEdiRuVAlJDnVx3Cr/EqHS5iprHAM6IKE+rkJa+WHtLUaH7
oH7THceRu+5EIgGYnA+HJoE4s8exxyJa0cSuz41tEmlBodVt4K1YdkaghjGdmHbesoqdad1pQAcW
9FBZp158Gse8BmLORRYmdNa/EGbOCH/5KUiF5EW7wLSkOWCVbSXOwpKQ/wXlx2ycA7xNIvkXcT+I
9zsDzgUUYTXfBTisNcTFD0ifKa4aTa+8xzgEB/Guwutv9+0zdLtqWCUwLj1eiZktFSLkotEHjyO0
fwEZ5VF00aS36zld3ghQgk3pByt7jW7ZqVRQ7cfWh+j8GIaQypkMP1fk1I0ATs8dLd91vUibffG2
rxlZ0Pro5ND2pN9k92cV3OzjMdXKAbS5r500729tDOWP2g8YThoiwhwTMuVgyYrrsAFynMrRiCqB
CfbUOZ5E6XIt5WjfR1asvUOvGiEp53n5N+qEavzKi3sKBJflo9OvHMNsI7QjSIYxnwLbCm/Jh2aM
iKFvd6vEwAFKCcWXAs4YchP68sQusXro17a2MbaZXDSdDizV2hdqZd1ULOhKfhaquGKlEVST0Qhr
+lk0nCsJFM09DBzGhW5Yk8wox9a1DuBOOVWm7ggVkfCzVfu6Z/qGXS1bj3IDkPYWMfRp0cz9hR28
iVn9Ux4s5qz9vhhWH6IiplSsSV6+3w1hlfoPs0PGvz4CO+U6ra0UH9PXt9bfKu+hyX6x7Ykv+0z0
wXSxeEVOMpmZI3/M4D0vYTm0rMMfeV8+FwkgoHmDkwROvBlgaXPuLXZHMlucVoN9UxgQm5T5gQ+N
o5kuINGf1lsPprkVefzVn/G3m2unhC2RXd5n1GFiosECcS9JDr6B6BVhdoh9g30KZM3u0XOPXE6R
F9prKOKrrnuSd4ldLAvWUAM0uoNu3TxqK/KsLAyqth7/jdS2z1qaEsnsLiWzrXa237gqJ8TvLh9a
iT38EBHtC25daYy+AxzywsZi0w8i64UqhZjn3d52vua/sqbkAYc/t1aqtwro8aDDsdqK0QP+ZO3H
YHJ7IBNmtEUn0CVum0Wf9ci6damLqlPw1osCQvAdg1mDm1A57bckRHsVuv+Xsi3hWUwX8X7WMU4l
nSw4gphEtrtybJX9GGUNgYT7aIbLjJn+BZ7jWISAEvGScA1ebuAf1vT1tzz2BGlCE1PraBLMl8K0
pYWazF9zMNZuJJL0N7zWLUzumAWwHtqPeOunKSYG+QYydbPkrLYG1IrqLBAH4qq0yoqQFfKevsFd
FD2K4y0uueQ+Bx/jfzFx4K3oD10uLqppy9RazrMuvvSfDoOfU2jDjYoGacL2/V6By43pOOqCgQcH
9AGTDr3W1FzEgg3eoeFJ76takodlzit0cyPIJ688sE59I0Rll8Y87kxiQu7s8EpqyOE1Zop4s3Bc
xHze0W6VbM0h4cqGaAreKoQRZF/i6uvHOQFemn2h95zycMbXJkc1TW6vvV8cmWMrOUxXyEwrdOoe
7mlHrMuSujbAcm4cIBzIist+QOJQpQdzq6Hx469KQ5KTyazSGYPgmp8R3wxfEpGZO69LkTnIShDo
FYyBMx5Pb9kj7x+dIDISQHN+lCOMzFjsd/ud1iVTRGqFj+sZGTNDHK2It1xgXiCnSurRew369Th0
juEMbEbAU/+Pf/mdl4WEgMyooikIye/kkhfyseMU7COisq5broq5n0Y36zmdjGqC0ZSgztV8SCNs
gbGrm7U7qPo2NfEaqf4fatBW92iuJXRLMOXt7zMFmTYspyvoINSxRq5F6bKn7Pz/rR4j+sX0vWuc
nBZ73r9Difxd9DsMQU4/G9XxZ2hqID39aSOKQbJ0qQyonoXK5XWDid41FP0cImiRhnO13p8/bp5u
qwA9vuxp9uNj7TPyhmECxLhWz/Z7h8dWfnTXpVrzTxCrbUCjoOiqOySZW6TcT+DsKQV4c4bnD9Ib
bo2ZXcMd2jAM5b1LNYoD/EDMarIlIYP1iG8NxqGGfvLvip4u4Z9fFp0jIJv2Wth9GxxvoP/Sia5Q
H0XyJPRrlj8m+haXIBfK7daq43agLkyutbTbTDWEKIcW3IjkPPd0NSoHdOAhdiodXvtBsna7FQ2F
kX0BFj44gnzOCl9bdq5O68vVAYd4FhWMIMtgzRKkfHxFjU3hLSaQcLRUcWOs83Hnnl4GGTTJ0FJB
orzvhlvVMtiQldpf0tRCg3HcA9qzyaAOUOuavlzGsUaOGOJ11O6VuajG5Kps+/qSWq0VbsT0IZjm
3AkJt9U9IsT3F1YcTMr3z/e2bcz6ygoPCNt7Ei3xKBVmvlHlcae2spm/snsosOu8/GYdd7g+rItg
25vr1m6ViLtQSROJq2osp2BAIzEn7Hsb/lh5+FC2CDdwvexHPy3BenyT6Mbq9P6B+UMD9RAGkBSn
vm/MECDQPV4GzTLZaVIUrm/FeldejC09BPndhmE/EUxjg196ys6NAmZ/CRWpVeK1CFwKMWB/A8pA
8J+eLGI8lkB6u/k+v4PKKpEl2CJfNbuZNhj1PUw/ycTZLDCWNAu5/YoIKVM5uoXJlEyC2mh4Y8ln
0THKLJBS6DLvFSCVU0Wgua2LnSjRGE+jEmpOx/+L323z2/IT23lc4S7OaovbJostFex9fZ431aeT
aLGdxlJb7XMO12jMv2pK1GGAlwAt35XKyziYhtcsLat1WgmazfV34QEC5pDZQBNweHovLrDB2dNy
lc3Yg6mEzi/sRfq3fjdi/Bh5RN2PJ/Dh4S3j2l4m3i1pp7AV6XQSEXezcSQJwqI9odR4tIV1HlIk
x2231/xmGdZRBmzYkNN0LEsSbsbIqzE8+/i2HUnTlKgzt99oUWsFTbZ0Z3docz4fXnaNHYDPUDMe
W2KMbz9wM+oYFQ2EoSHoDgTqf363tBkKbj9vOIGjjSPwOcCMtTIowglv600yOVqgnqT2vKghQ6B+
AJ3q/T4X2/TnCLhPySMo/fGGFQkS//i7dtJymQNif9/ws8liTCX1Rhu2wrOSXQA+B5/mHPVSu8yR
L3dRMH0CmKmZd1EtoZYwpmYupm65qAu34HRZfYNlvU50J7u3GF1JR9R6JpIheCFpcc4uz8BbrzPZ
ymHFsaVtJL2bsTcL4Ccsi0IGz87MhVEsTadVBXtnTfE/LQfVpmOGfvNf71plfQUCFj6CIma9eCLF
0tHsfXu/KCA4PhdTcIA43F8IElvv4SNwvN4FgG+zff0XQvzB1XL0zdoCxAUYoRiWvqp4m2wFtQ0u
my3AIEhrhxQDZi5S3bui++uMzLGta0v6Vb75E4mSzWlzVEKaUHA8W9cut8ebYRK692wK0ZNBblDV
LH9cxQp1LizbzQY50RLIpzk0fNuDIe6jO6ODX9i+fmumNapj9umSB+oSYaFlTMYRgMI9m8S3Vnnm
4jpD1Q4odIE6emE7uL5JMlEggYQ9sjpyWaE1N+jkyW+QCivGvqgpRrROQG+ke/l+v/UN6KENnNIK
nngFVO1D01bH0SijSvfdXrtX6lO5fl3JFvtXTWAl8+L8R2QK0X5qGhCoNW0mSTJLSiBl3so4f9DU
Xp1HGZfEQKkxkSECqP0etccLw+ucJm155T8y2XQwoR6fsH8CD/FKnX3FrKja+IEZb7QL8DgHPJhZ
VyvJCIo2NjzTT9a8TfHFLm0gOw6rAz+zALqiwNhq2nYr5Q/7yVnOvJPUsA92x4dCmxlT8SXVc37Q
v/naSDPy5Be1KwYiskYaskHDL+6JZIQmuPFLP98qXqzSu/keO5/6JLZ5Bai1yNQDNGwIdp1zSl6w
HBoushR3d0fwM4u7CO48FaYRkt1ITUmDxgvDdHg8rjUXQkxHFPmVkS7aYAbq9lcrqWV2xYwUQiej
6xN70tmg3j/D5kLhVS7BXHW0zPdjQhzpzhAvZisFRjtpM60Qmenh6iKSpqOpOAyz/DTk04vQC2Jq
momKGMJ2q/Pi8B1MYxJfbJNGuF7vQwPRtdHcN/yi6tJ+NBaNU7WgzOGf0hW9JW1fncUOt+eUkxD1
sI7D4BLrLZ21fBoWltP2LVz8HJbMVLXMb7dEyqQQtrBxlrxFBtfu8CVgbXPxTw/kip+Q97BJN9NK
0d59N1qxH9u0VmtRRvkdCZCg0TZdPKTt8kPPxloETZwVWcK+ZKJr1o+g+cMBYnoB8s+ipQYyDo6n
yEs1yw/r8s20vmwhZIR8c/xtbDyLo/AVMxUAciuhPVdNC7ebnV54MASYXwxKXKglRqzK3Ow7A3Va
0fEQ14uR158YCUWF7gNLRFy7MtYxbRmXXsY33B0DAwvGYaDLRtET3eEXCl3DG+yDTZqZsHEj+FNJ
MhkQWtOgsTnP1I8GhtMbzbQwkCBhk3Fdec7Lb8l5w9w1DjK3zYhpurZkzX99iwRiFg6mdPMtYCB4
YpZCbiB6vlJ7DTXMVEbpjU8jdNLrJrsrVfYWzTs5D6lxGUhmrXtn+ijvtK2OecssiGcZDskxJ2hM
/e4i80LxttztSeHswfjP7KTIbii/ikEgvZhQbGM/S09tGRm6aLbN0N5IVKxcuKhhfG5p9x8tTaq4
vapxR/YxU/MjipneuZ/EKMKCdYPuqcY3+avy/PfgINnH8c311dFF87KHn1ugEoILHpnjRvn4DK2F
1Py06KlszSffhsIpveAHH3n1Ntwa6u2maKnsyhBllhbfHdl8jwKREgEG0M1DguPgRF2O4r9npgXI
UhjgTk6itGcG3e1Qlfq9Xg9Vw4WZnz31eC81FJhofB0o4fbKB5X5ate5SNGK8cnIsRMt5HpfnAMv
FOXUW6SBTj41j51nmYNV9cpCvXwiW/DyhzeniCQ9gCShFP23X290vk4KYqdocvSDf/D5/nX6dv43
5sFXEQxVZmq31hLNawiDxCq136RQ2LWkCThpGUfHYAT+Jo07BqLTL5iQlV9LKyoP+KPXeADGL4qQ
ic7ugxrKirKuezPnL0hHmBYOacSqtk6caqayORG4mZtJh7FNw5qRPKYmlhzS8tWH8Kkzk66i2JzN
HgazcNCyNYPR02B7WykCmf0ENMh81ij/O/aNNXR9lXXUFr1Xd0AiP1xfIzCCrvaJet7xl81zpsO/
hjOv8sKubuL8Y5muOePdx+21Nvo1DyQEddi3UTiqJEh51eXheecSdZ8942UKz4lX9BCQdxOODDzx
AUL9CXY1gesiZymuhsvRB8ABKldlgwX3JyzlXTjPuEyZu319LYFjnW1eJLaV8XjhOAOknje3y5Mw
i3PW6OsYnYzs6K4XpywE6trHHLRgSeSPeAKt+/RbY8qaY6QIyzHhSp4Lelncca3IAjpyCJcdF0A1
3/YqSlcxjZmTOaE13EL2KpNThNjGmHuuk1ugjhBZzJnnMarqnMzpm6Tfo8GkkDLBKPr5A7cJQxN7
9swtXAN/gkD3gMOlASCVMDytUafeDm9LD3ecVtN/bP8cUegxrOPLFnAZExekR0PN2+bQz33dcVhM
mioF5BH8RymVBtWTWLlyUI5+bEnyyuTC0AIZRvfnrOJVxdrZUKeFVS3qPyGs+Es7ByPOjCdGklkI
lz6oy4AALCv/b1wGmISf0hqnOhfHr8i83LiaPHCTGaDtBzDXZyYSC6fsdtNP74F+G/5Vkm8E7WuU
fj4KuBMUer17m7mWO22kQuqlP4rj3N1Wqha6RPkusyeihYikI5W7GqMiKglZBIjlmvvNsH4TRele
9Urn3iCo0T5z07g8LgGR9onIkYKsq2++usCQcPQQ0WayH0eHmYuMhWCMGPcc7cUInQS3dk5BGfHd
7VI5Ic6Y9Wk2ZqCskwoqbHuFQs0kzuXO4fX4OOAcMqmeOavhpiTaNpJzuyqITqj+NMCnN6t1WpZv
UnK6DahQRNYrlcG3sX86upS7CVbrscnVOMqcnYNkccLuvR/cs7KkXvWHMVs92pWRHLCT7vxqIcLP
rXCdR1Vw8NVylt/J8BeE/RsZb2NTWyBTz/pcAhWRqRUlelMJKK80TotU0g9K+/VKr2exQQQT74yx
PYxSkYbtaEEVsKNQDTkCGRLTFLBO9Uqr/wVK0u0b1YYCgpqkJF78D3xT+z96KU0SGylGlNAIa67V
0X6JuVqKpHcnpPS+ed+J8K0jKMmp0htuk76dLI46yj/C02/xxud228Xd2keHWA7NfiS0MbGlZot5
m4oBQqfP4XwCQ6ouWgnM0UKLKGpn4VPBdg0cy/nJn3n8mmcODj08cVft/lbvIHfnzmSZfC1caSHA
y2LjEjNmjKAIQ82Eq7xv4Ki91e8RWL0yOIdI1yloEJ1R6M3O9RsvuHqmUWyuDqqjvQcQv6z1wHDt
wTwA2Q7GlqtRK3BwnNiFzYj+72TeXERUY+FADAL4htNHqPaMn5kng4jgFa7YqfFohDubS7SeZVzz
EKSohreqt3U8jbtA/V2JsdtoGDcM7nI+qT2Rnq5HWZAUN6QO7v+0JcLE5lweVhSI4+cbjsBKSGdn
2jg8oBAjrnFqowbwauxCTG49pA9eqpKk0045yLfHeeuGb1hUTHHJARwdbpZuXJjmDXA/rjOnqrU1
Hf8FdCGAMfILZ6jCQFv6zPO5Ef5Qexh4kUgUwkPEN42z7zHrNsPmTeSQaZKsyVAv3NPchmErVxbg
i0l5dTcwxeyp3nghitT/7E17h6oM1/KKSISawtNMxoDEHBnxUDQJu4jIhV0Uj7tH9/C/sF/iqc3D
m9TWl5TLuimP+4Y+x5H7yJd7vx8ZjkqL0qxgFK3LoO9W55pN8bHbsu54ABIsTKofjmggkWIiR4zs
LuXfOU0c2w0erMIw9mSTzWu/OYMhtFgbDtacUfVBsJU/X+d4q4+dmUvhK2Ik+0eg8oJsBYuYiBb6
F5SnewLAGje4spD77ZzLDd7giy/Rl+DRo3LkgIXtup0L9k6FApI3ehflTRRdoImNv+HmbKUdT555
C29rOE5fpJP2ckP1e/ZCuNNiXuax0dR02RwDYvZJshuIzngnjNYCwfmwPGKIgfFV4f4NUjOwCafj
E/Wuzt7zWhQRDja0kN8Tqfkj6yd4cfyyRnLXXX2l2xiveVdLIME4b1weBN1f9LTUdW/Jib/TpT+l
Z3CshVRyY92nDmBBAXmL/7G8zz3J3XMkKWtWnCN44DhRq+89Sbj9IMOn68B+P13zoyXlnp9k8gzy
DpW0psRaWxK7cZDena7vp20tPyau0I6diqoQZUZM75QwxZZ6u6VEMiD5rDBJFxGcg+ebyKXfzN2K
vslFaG3WXNxg1gK/EgaZxVtZ/z1Znf4X+7nEYsRM1bW4RhT5tM4QehuK1fu8D0zfzm50zrFOMtH/
0e3vRwm6A8auRkkSnBK6aEtGo5ALHC4+kA38XAuXsfj6abAQYEDRWTPByQxjqJvw+GtjvA5EHEd4
wy9URKSJ4TWcDmUw2ISCi2DyMzemqWn9vHl109fHh0YlmVQxlQKiXY3gMHz9QtKjb6dOOL94Oyma
d4z+GkkOFHn+LCBunG0C88N7BGxlfc9gTk4ZjXmW8mAI0E4l0ILoL6+Xxd551xRDG+4l9ZEKl3hm
TAjw8MFhiKDcizW7MJMtzNy8tAv4De2uzZEnVjdIgIuev7ymd3WUpj9t4IpqWkhvkYPU5NBdgO9W
b9cg4iIylEOuhuY0P4GQs+rr04hFHPtzGr/VOCLpfKUBU683oK25k5XwFCOjZfdC8o/cFlYziCMd
q/+GT3lIqvZELegO9b5S5UppcowmeVDY896SULWp3Ui6zpGn68BowYulR7v1ZeBrE5I6j95b5tqM
aQrSVMVb7prSpDiIK4bAmcrJwXFDtVm1h+fNFaVMV1Cp30V2tFExRYhVwvho606U9BDf46djF6JS
gbSU+jjioFwbM8eN19Lqh3PZyntgWDArYCNe77L9huWBYgxOEhHt/4JLjdnGMAkOV37/TVwi2ksf
eKA24NuL/9jLAGAzADF/QM7Pc8dRCqupWuTKKHGhT/7lE4ZU/43XolVGdmmw6hyxWlNIcnrKEozh
7NiiF2mjRg0fjVbTkDudjntArJmNgQ5F9zsogGyWOGPIbu3mIbL6JDhFDpQPMHIWawvI9Qg2F92w
CSYElpKaxaHrOaOclglGuLL2r5PzUcZWMOrIr3KpxX6pfR3SAQKtWfX8UQOqK3tuDw5sUZ9x1QMI
OTHguiLOdtmSk2Z/KyZ/2lcb3ygxInv0Pk5fA1K79xE8BbdOWskSJmx2hjej094mRI9vzAWh7bP5
KXwXWVbzC5WGMUvToE8jA+jDqHAexYouY5C4RTCtSFQcYGzSwxqLkA8MBeuKbkQCZ586b9EmMhng
ZGcRK37uGOaAaTRPccKu1ufkQHh5MZwrxyiN+nHX6FKMSzSi0hmiN6/Jy0Br8bjWFwmBdRHstpe0
N370PLI6ZdV2GIsatczp6zEAFsKVUwRstL/uMIpoxaHI9SBb0P4/qgrG4J6CPtEDfQzPOyvm72bH
I3YeKG5+pgI30YyuR6fdzhQMfIZn+z3xftJvV6/LcQa6V4i4v2q8dGc37jhP/157TvSQQpTxS/Ex
0psbfR059SpGyWm97FkG9b8MKbmMmzvKpB4CKfGRa5ZnrwfItL1EufgaYb2cdgNfOuDmTN3Y3TQC
IXZHhEfaeGENvu+3YwirSwjl45kuUCdjAedpv3XlzIOtmxtemHFMPp6L75lHRRL3IUfPQ3jEmfCJ
ktiAX98SqAWfY8j/fkk0eee4LAYkSUS1ThTi6V67ABRQWc8PFzuAqozW3dpemZlIukq2U77aAwF9
zdEOUZV9eUYyP52X19f3FLIHWo18EcoyzZx5J2uYxYwL/mcQcnrXTcY6A8J2OqKh+JbYMkSAQlic
LEPVusrtE/YGUBeIGD1J+7aGmMA8G+8mlHxeeHYB+p4v1ROXOPk4Td7B8tXnhV4GnSfjqCSlE0EZ
+aUd9uwOvKrVlOng12Y4exIsJehPxo/c3oZLqUf161pRw/Vni63MUnUncDLsACxoeH8nr03+HFux
wL0KPTkosJjJQsP9zZrHYNztc5XYvwtchnh4+GVhivjJJ9eeWNHC1/buJbpLhLPyItpS2PdBJEzw
YK1Yd5dszKtvKybN3Bk6yI64+5ZgPv2zSkzkFgEFdZZ/1joqRP9yBVn/9EDWfRRkccM4oA3Gp9PD
6PfKkNcmPNw1uRBFQFDwDMiFYmzqXDO54zxXcP/r0M9T4XcfOCMkPu3vW09HtAzwNQG603tlJBTS
CkGMbkDpgBlDlmc7A0OWmK/5vweuK5cww65hGm4qyW0QYM2PHzzhkZPpElRjMvggeWku7Nq3QNQn
EaStEow+T65KHci547BDCjNEGTCkESAPNkO+aOFXXEik2DTNX9q5Y08Qz4aJOZNpdFeEt0rtX/su
F30RZAfGBL5+Z77qujpClOESpWv7NKyfv/hK3by3xdwT2gXp6GIPAi7clIqZ0fI1Fz2v9WFTwR8H
Ce7bUReW0IqDNwoqu9yEisTtQE8DNCeFVpG2D5XM9HKBoo+ulM+C2TIYtmTzXENW5JkJCSdBP7N+
v8aki9q9I8yaVrnntOKjNz1LtyPGfgVEVRhphaXKD7qoGCbHS4DbK0AtkyF6EWe6oOUdOZv11lyK
cX8MZmYALLkhAtyWA7DLoQixzoOh0TPla3hHgoHWZWGMjMCo3GmT37dMvXeeOc2Uqyl29kWpTc4n
O1EPNO8bzsZ+1PjToE3x6EbiAj7k0YmEKbSTIhW5S53BMNCGijOs3QOla064EMkIR2OMOVaL9h0b
xngbwXq1Lpx1PiyG7AjI38kvWx9ho/rwG8DOWfoA35AJEZYkIzXWdZFAwB3CalJAuuG4unWDIz+M
3VWiy0GoUb72yd3EEwEKxOj+1Bm3TzMM9jPlYvKha7RGY6Fdj0k2pkZDO2UT5L23tWejQtxAG8HA
yeRwiLElaiaBYL0YqvDscplV9zpiQQQaOP8iMyjpMPjxBHcX+TCWJdfGtPL/Ajj2Vlkgclftu/z8
GxM0/XJHBlMnJ6ZS1ElphG3G6JaWwK1UGk4twjgmMCDJ/7Aqs8eSbRZZt+PTh1/vlgodNZ/T+8KJ
+jzLIwxiFMQyiOSfFR8hVFZNmwDjnA7OKOk2ln2jUy7JZMHJe33dAyvQ1Qnwb+0r71GNZvEMHoJF
Z2GPydAfKiFlmjwKWb1TCG0KOZxL7c4+Q+tOGH6ngYJk4+nvlTzOPmIAVmoAUSAYKIJDwn8jVc+a
FTZ/t/IDNbgn60DI7/bWFjfqtAs49GOgMeGdGYSCzhsDAqaieBOVHYEeRz2YVyZQtvsI2K4lxv+d
yLoHs1F1gBSvsXfa+qMugiU0dRDe4tavHorBypb0PBlPKSWwhgafD1ukdOOuhH2YdjVJrcX1mrKL
8aV24U83ZP6UwHxsusZFcQfm749YJyv2O7kWi5bkYYVsGx64i5k8TMYJnHfvlQiAearvxwSDVuq+
wIPJFuqpwp6fSB4swewK20ZvfHoMc8UgN63hurBjyS9QXcz28c/nqq/AvZbZ0kAs3VW3YCK1xPIb
31pp6fo46cxQiFtVgwWEU0yuNtJrDRmYnMKCntuxN2baB8k4cq/YGxfAMmxPXvR8HIdk6NnRYxXa
MshA911q9gsO1zWHFyR57+HjCw8ehuHZlhmqRnCMUaQJjWuTC9uuRCE2y5pzCHwLSZlyabwilqUV
axnSaeyB7zlsMGAbQQE4R3r0prI5F5eMa91rA8kpZR2/amrXD0YU1T9+s7GcTv3V7r/31GEbajoA
eN4lGombQER8nK6u7bPz+LsohhbpFyuXyi4nSS6YB2eaUs8WOFM/YazomWo2BI7l4S2ujxpi4IL4
S5Dz190uBhSiqRQDg8mcoWJZuMU4YgYlAJ4gfQPlnSxhOOgzZvHhog+N4qevoy2bzmpYDCctx2vy
fsHzBOHzCMzJfPjJMvTvPBT7L2on5rBtdq4LiRsH8AdQJOj/BfmDCfVURPHSClViGAV5Ka3pJ+lk
f1elqz6bDmpyCKayiXcczBY02z00umdoc/ft5VbGwRRIIfVJQ27nYZrGa7ZEXrQs1wvJo2aw6GA+
zA4j/lq3lOjg4Vs+srTRg8zqEf8Dn/3wrzdnxyhT4tVoqslWmGrRQiie+x7tt03PY7CdAgOB4Lbq
CmHmmmkOA293MN0lZS8OK2pSVaWjVpE/GwJEbQpo2UTA6QKl6h7Sir8h0jeXM1Uvh70byFKCXVlR
0Vk6SsFPcHoTGWarwqv9ZfKGc4ftCZ58gjmsiPG4Ke1KgGBDaNoqU9cCwKFNx/l5ymRK9ITMu3Ed
FeDU5P473rBFwndl20AOGOCPKebxAcV5mxovGlO0Lh/v6wr/YhwiAVg1MDqUvQ6cWRht+G7CO0Gw
brVQOwxv9TndC5wR1h1JJk5DqPshtuLVmaCClzWcxWOmQsTLH3OSgyg65d329M4C4G0nVOLa8NOm
dXMgKVOkgI4q8vONJ526hrTOaByS+KW0h0z5MXqtZkMBTX7vt5AywxHKK/KNi3PeSDRKHYppHmCN
oK09AaA8I7HtiuKQx1GVSGL75GO7YXq0gDb+9DOOUL7yqhRC8KCiOHMrJJA0N4Uly48xrONk32hZ
QXQDV75cViXZQNaeEOwDoFYWCGQvPhhsAdwxb9ZbZT01IAetGvIZWjOjHoV+gTLP4d3TaT9b6pxM
ggV6nPxUsl80L2386pJ0eiMlGCAeqrC2H9aye4hw4YJeNJtQ3Keum6nne2FMt/TyjhlT51RCtWzn
OT1Ki/Tw1YZco55H6aPfzwfNftRCh92dG9rsBe70VLQB+e9zd/hPVfnLYSKIS51nGmqPL0xmD4Wn
PxPeg1p5jrjj88uki7ezwp9VfnAijiM76h/6UJ9PdE72zO4XuR5m6fN6KZd2fShsUZfkKWV1vH73
gD1AhlahA4d5kb8M4XLqqrV4hlEg3Jcc0Jl5NPfX2ur0/MXcJNE4vWmHDxhE/OKsbvtA/L4YklA+
vQ7FmwCGoKZlWsqrcUDPMn3+MH1rrMfFmKdMtlcbnHAIpD33dCEVS98oJK/xoBnmCwi5p/kXg0Bu
bvmZ7N7VLFcrdWYPf56c/9n6zMJ+7u9ek1ipk20gcxH0j8QX7eSJz5LxyeBZuWJLBQ/ppKLCdxSh
5zrVtMRkyxGmZ7eKB6BKW3y7VYf9P9MDObTfAChFhftk6WX8acOzVqgjT5rugfANag/abfBoHBRx
sSnyTrbU/zZCsnqnQ+RPK1tz+18V3EEPLM2n6D1+mLGNNx/ONUZ2Q42S6x973KbwGjsCYOAqUjZI
/rOzzQRQuayiwhzTkvXX3Nv2b1QW6BCE5ltx0R5ueupQG5NPLjoAJYdULdeRtrDXlWNb24c4reaC
j6L6XxA3WC1LjM/yMOGQ8ttCX/ckuvdcalht2azrFa6XqAvflubgsNnjxlfBITMx25p7QpKh56qJ
fVXwiVfaKeyt11MIBCs5QZwjwm7ekmqSOov4JrQGX3ouOGlJTvO0Dk8N2gcXkoqhunU4cTk/yjmt
xve7WWHzCg1sw/1BL4uwFYAJDJAB3feWSprjwyJkm8UlmGRBGPJDVWQDio2WLT5pMbl7T0CrEZsl
OYWJxg6OXAJ18+thLDl+S1GhQ1+1EllTQk1i+yUQDoOczKEELhYfQj/uWL24L7hVfK8j8mfHOF3v
fSu0eKZM6/tcmXEUG853hf8yirv9HNA3gr93Vk3wGo/SfU1SGgFfRIzBaTEIb1aNfVOX1egBmWQG
meEpP8vWvkS7ZrExKKqsyXiX5Y2qgFJY5MBbvz0Am9PS377lhGSzLtUs+DbS3c85cDxokGaQIsbh
xFt1rgXvwZnI1PpOUzAt8Mt2jr09ac03svlhOsdbYb8Hxv+ccqEo8/0AOj9dygAMwm7b7EzYMerh
Zo81ZtGLZlX4EZE7RAc705AYJ+VJPCoxmibZw1zedaU3Vsje3wsuV45S/4rCAWls2EWnL+MLUbIA
7hvfbeKZQtebEpGdsp9FjBc7N2CyhgVusM8tGKv4EiYcZpU3/FNA7N0xkv93wyBrlOvm+WzuALPU
4cDy2v2rp584rZ8ywe5NjQirQOZHDdp8tgNCddtbLrz0Ywmt+M2uRU4C3bBDUUS6FXT8GgKvfwed
Flaldw+ymIsiXHa/kntNHnUVK2yOEILAfwQSr05ObY+Uk1lGGDc7Escn7GRDQrIRAVCmynnKH/AU
PHUGDbw2fmITqyem06iYuRTNRJkP+PqJ1aanW6twAJpXqY9AsXxIC07rRQuPPzoyuJbok12pODO4
9kSx4AfC8x+WzCOI0tk5xIp3MoLjfotS4LlWBTnpUFjLZL8HWzrjdu11WjZUOC99Is/U03r5hWPK
fVvjbLbOGZR1Yil9gQZ4nIbFVivLk5FjOeccoF/bwyzZuPRNUgSwF5g4RCAiocq1i1FUxNfGAzL1
8H+DaBglYZzPCbArbkFxBba7W4oBKAOfpHbfza4AWLZMNCP+KdHtOBL+oy/ZvgLRlhDHtIwTfQpu
JD8fqXaJbFqJpMshPz+vhNdHBWKve+XFQ0lKG9lHvCUG09Jav+V8SPtlSErkilcHAODoaG9T3lJu
RFPiwrRAaNZGz6WFNgyXRtEtGGKkZ0pOESAVxQN8J/MylTa9S98RTYxCk0IqTy5r0yMe+4Z/nT2I
1uwf0BdII1ojAbkr7so9DqGDp2W8tNBPUKJgDRugOUcIxw9y8cbUOV5WsWgm//zHTQ/O216jzieV
prVGsJeav7EMvKRYBTUXwEcSR87ZsMR14CyKEBBlMw+8ZHfDNg8SVroL/fETlGvKuT/00Tc5IUHM
N/T95NAlfqUlLKbmU5HmgoikFT6/3YdvvCygjVBtb6gcDw3JX/7rxonEyns2U27hFpF8tJUCqyw/
V/H8VEocW7Hgi+AWPXJs90PVpwBwvP2ckBQjvYFfa2qDugL+aDFliQhANGiPgAPvTi5SL7+/zlYJ
C43dOlFk2khp1XGNtHNcAMevVmDcVj34vg/Xv73MEAlzSTZIawKX9wNZqn7eh68/S0fGAZjeyk9m
IehjPFdbtYyw7XyVUyJq1Lz98ot7VgKUMruwUctgTUJQFJ2WX8n747qcmGqpMZZz/K8Og9iDr0rD
dAJBrfqaIr7sppwouIPqeyPFP8J3kTZRyauzZtlWmipg5gvnYXF0KZUNbOCp/cjxQXqHvCx/XMiJ
2cQw+hrXSGwsCmr2NXyLaOQSufJ3YUDBDkhhCzFFuFVUdyf6ZmBpoulfZc4mgn0Xo2JCOdKpFQe7
i2INO/1eI7otXrb5mzqii/ETFF499uaTPCPgTXqOciNpJbpk4/b5fWWWtX8tQVObRC93BzVxUUIs
wrSdVu/RC1z6tSvbwwnq5tAa0+36kDdAAFqeVcr4jiXngP46We76w3UwbuFDOUZ+zkyO8xOAR4I7
ScPsEG3Gh4ZvaP6qZXtxTo21Zy6nevp0DipkMREiWc2gHASXY/djk1UvpzgBggvRqMGCeOURGCVv
EcxssuJh82CdqmZGkdAwbJT+1114avcAUPHqQo1+UWyaTAZCsoEWVr7RjGXc7OTZyGMttf/vsM82
aIRZlW6eCNLtJwDgE/O5EXb57+Lux5eVd8aHfoXwE3gQnzMH5RWLxCFUThaiQz+c+LrE46dFDOFj
nnKqdMrECZasZSpRIbJEyxcOjAoS9/ezgWwjdYO2QXKc78IrgG5ik+OPRPebWO4lDTN4FFdKwUlG
Y/NXhxdL6rvTRggHdoIyjp58Q2OWGsMKNeQHJdoExd/qBftGUg0CTBkfjbYzS4DR9GfYZmAExBjv
Daf7fXCS1iHcF4/Ypstz88GN8kQpJbyrTohE+hjxWeJhCKUkYMERS8O9Zw1lJHjGcV6F9qSugG9G
hA2sk3Vb6LWxayHT6tSGz6eSnbF78jpuy5CqT/jxg7g1FDPXVHEI4Hhd+AhhkJUsrI85jII1Ofzq
5Ff6fz2/mvOncAJq+NEPRx0A7zBxU0Sn5OTy4KJ+kjUC6XM0Ld7vmLyw9q9dw2puVMRi6BDJoo8+
Dz5VXSar5ub1kYVdxDJZHSrKupVLPe6cwGYLCgJI8WegJtPwpFcBXmo1rDUsbqG1519LLw1YLQak
RrY3knbwx2lfcv9vplyHEPpM86IltIHlioAx2Z8j0zleHu4toIJNyodMuDa+dntyKxR3X5fzE0Ig
TFH2rw++hkPuU12D1O80zNkUlEM5FGz/9qbNVdbe4XlVmh+p83nwzjUzZ81SCFCFuzQY5QYl7jBw
elha0IaS0cS24pv2/S2jFXDhjuAkhdkiuFoombnOHYFcnHKBF7VsluR6hsvcVNXEjOrKT9AG1KfY
rbcphrEMVUj0cm8jr0ujgkctIq7Kuj7ggAqP4ZP0sMBPZYAXDWGvMfxxKsntmonntcRlNd4fknK2
0jQsiY618RIx98/TxE55jMYBwZG/t5SjhR29TktGU6nmKdQbSz35psHGpJjX9Q1BxKiz08dc/G4/
WLNmeycsqHhr3r2++WZkAFrM0qmAD3bxNzViys93v8NeZuotDJxPVbBvbTbtWDccGS0bkqrpHt+g
WVd3XBuj8mqFC9FKi6LMCClswqUxZSU4750toiXjtdu/6hFEoD6FAUMTROqJXafnAIOccZRsXrFn
us1i9e19BUSm5xLX3NWzfe5LLMfG7cE3puHJkvmJGvK43YNzjY0DF8AJkaQglaruE6ptbQbIXYpz
+fsmiLx+KEWRAz9RRwQRvQ44kp5Kw/tf98gDFzyFPvHo66C2333YKFSnSe/mGkcWCS5fTJq+29Dm
TBbeakRZSVE0aYFm7EXJ3QOS8WraRGNRKG82+R/858xxwFFHkekZhhSjk4ncQ/OaAucYh7v0hJqP
pYCzL3LlATkMLC/xrCUaq/OEfows5L0WAG+GUkxowqnxtWGPOvZXZhPXCpotQTHJzRN4NKUa4Fyv
dRZ2Yb5yNWdoCXY3B6qB6ZofJBKxIX4eX9WGebNB5Narsa/VvRCACSW3DFULygwyBIxxf4qkKFKU
5fg156ysGPTS/39+HuqdFPKazuVhzsn/pdAZ7iSy9ACUhLf6NpUk/JKwWnD9IYg9cKtLFqx7TjNB
NAJrXegDAUajOtxQzwdkRdXGgV+1TreX2e9W/voT1CAAYRFZPLZhlJiOUISLAmNuN+Z4RfnEo2EK
idzHQp9VQLSmFBeJsTYkHwnbSYdfbRV9oNUxAzDV5hwpEq+jDzcRayeZN3T0pXljCIpFulLB1uIC
kyC0UqcQbjFKs4WW+LClBC0fsWSn4z3tjHT62sbwJXu3MAmxizQmkAvxioC/IzhDygVw+VI9VRNK
tTEvDUxgl3hnYuOWV2RUs8R03BJL9tqAdutrkBgmroZ+7W89+8wRBNo6ujr7X3q6qCkt9kiBlTdu
+YYg0iixVEa1FelD++HQFDzsT4lJxATCICjckNwFNFFIozt+8Z3I/XnRiNtby1zBw5DvHpR32Z8w
50nTXmi1VZboCZsCJ/baLBiE9zR2y2vQ6kearHcIp4pqkuj84IoKCB12ufptjq7LpIexg/jCYTS9
GnWH+BXWSLrVmTxkfJP4RrI3oHjANygfA9+nHpkVCM6eDgGmUDa90U2r6WWCYJE3tcYpqveko5dA
CowT+BLfOdqK0XI205emF9aW7bOIgip/hTvvKSmWmTwlJq7CjIHOfgMA/cFjtY686V6GRpfzcReY
Wqg7MBskDnyOPSgOOYf43emCJGpIQSmTdAaLyYapngpTut/j4hEzJuiH2LiI0LK30BoYo0IEFrOQ
j40wyShsrEqKwR3wvxaB34iT8PxtGIfU48ULcnDf+o9KQThbbm+/IZFal6DO/7DyU7RSJ9+hsDxk
jXcZoQ4Dj3CPHr2hRi7A98ghqzOzAdjtcdLM/IAS/JaK2apJ6ilJY2CSfwM6//n/V3KPjjjExf1+
QMlFerw/O7oC3hGB9MJ34HuXhBAx2wxdA+fonvZiP4qjXVsEh46zeOZjxKc8X+RKkeaZ6xyOPJep
qcdNBNH9lYK5Iqe8A2BNTyGgkHkYN420XZaIH/Sc8z/ayf8hVMrmcHAz6cHXPYVotcTOl3h1uM6j
IxJNUE++OUGd+ZIj1QtaVTubfIABigRoULWMx41o/esIj3M1uTfADj4gh1vfvk8EFBEjOjDjoThR
J+OqJD9BNgZylRlqnA+u52kENd9uXp5mBYihUrRoG2MQMedzxz8e90xCAegRiRTBnRjEs1U1FbKv
IGpweYl0FkVK1mZfO2eA9PtLLJgrbrDBQCWZQg7QUpMKF2AzEjLDRvplXq51S0JGr2Mo6uYHet2B
HjKvoICsnJQbPcJ5NVsyfJSrZ7uLRjevqEqvh2Q9m/RpMybhVn7LJ90yLi5b3jG/Lh4YzlSjsNYB
Q/1/QvIOB20rBJvoCwRm7G5mC8iFbY5GKvzrRLU6jWPuAeKqvvM3GUpv6tMz3xxKQJv+y7vKfx4O
Wq5D2uU9PsQJQPxGr3jJfkmCTucn3UQiu9M7we4qYnWwn5U5MtHmnCm5R6NpWF6jh7siyupIBJMH
hrubqc84JOsPvS+Le9Xhlw33rnaoXQvUwqFdTCt0Uu5yVD4o3ACrAH9eeoXYilp0z2E3nBauebxJ
qJbNQNaJaZRkQ5TDICDEoMGbGUdGdQDAdVlgs5eUuFMgt3VU8+UFXu0Gx8kKLm5m0F5UDqFn5H6i
5/3d/l4DJChlYCZFKIbwgCMwxegAlX4Lq7nYMmfbsQyp1sBrHfgS17LMkn11GYCz3JYX6t76hV/3
vQC/pryv4Mr/wwBNYi76hrcorYvtAf86cZuoU8KQCM8msgPoPZp0USbui/yr9qbvLVgp8+ZcozfU
YjdMN7F8JjyCPdQ90+VLR2sNdOt26sgKSB8VClVF7eq80b7suOhY0zZcLcyLNThYPB9DbVe31C9F
TDD59WtMSFh/SZH6XDtfJzceHmWghEI8RqDb8QcOvM0Kv0kMyX5w/8rx4yBeaKLgAYrc1j37tekZ
sS48yFG1cCgxyv6cv+AlQyh36Kty1+bcp/kUh/C7QtNrXJuxyeBNYeIpCI+daXhp8roxNTIQAWc7
Vs+1kmiJ9a5vtHlnOVpf4+t5pFd5/MPiFccOS7OGPofXx5ug9BpCt5RGLmKtflbYz0wGQosGRJOj
mx+eqt223X4OXOknXpUZ3z0eawhZKH0eEzBlPVQxp35ni6IwxOFoJDhBmyBfNUrO9Z4+Jf8xjScr
5AkpPHAaB10AW3M2hbir5lRxYhTEf1VpOd5M6tLz+KMswVkcngb3oA/JQSZnaYnmPRlvq4E3TAbK
rCV5PtXQgQbGfWUHOB4uBoLO88WFJKCe5iSSTEY3+BWS/hpPXHZo6g6vrq8T7BKkWdc2EKCxAHJy
4m799xQ57dOzsWpL7hPBY0l2J3pguXYeExTg5gdaayofjtU8scS35qJTzVEVEFbZh0SmI8ZCU9hc
BEh0RIFI8YgtL9rOq9RUV4dYCc7UE55mpCLjJ3X/Uj2EEhpgrqxytZ/RSpJwu3D5p+nQzDOvxTpn
ABK6J9g7IFaFd4TX6BWyQYLVIqYRcM8LQFsFxDZvI4NK41+a0c+O1ReuKJ1G30uHdiw8jH/LOxZy
bVPJQygs/SKk5CqSUhBXglMiJXFehmVeakOn6cpzASTR7Ig0ND57oYGesrKDRQ+gZ6ZM2GWe/FPq
ja2cxq56vIOhK7Py91Q6vEtnzyLWKM8RodCyJhniCc5Y0GhzCPQuoneqJEbD0ZAzOw53+5h7dKon
TB+mFWsDu7ctztS0ZbNg8KlLpLpfrDKpEjd47Kpt/RKjZyxn1xZCS00qBKGMVXkeDIKkbPzxHKGA
Sb7CAB4fRJADjSmGMyN9XXvuHfSsJ/OLmSbjVGLHmjw6bfu14sz54nImyii1sgzcqK3Uu6aG2zmH
4HJM+vDVqlo7zT+amiXuMbeZZ+OQthikB7zLQ8EIi7gS9e3AkIEaiW7D890+7iqcUFoEAZFD1Xwp
owGnCoZJUXs1FVPP2QZxLb+wkYF5aU/nCH3rpmHAKaaBDiiHD0JDaJGUWAvxy86wlSA+MSbIWmqH
kTwJc99WdmRMBB7fTAUZ3FlwKc14+WucZ1NgDZuWer2HHjKoS3Quq1lrfV1rm5cP5MqifKMZILbD
JFq77ygIxjNqWW5ACrtumQ/+gV6I1YL9zfkqi3YILKdRCJY4oFaq7BUC2p03g9EHipTInYUOqX7P
wO78faUvB9qkEsUsrcw/VsUzk32kgfgvwLpW1xiNn60qQ8budylI+NYNursC4L4hAgOIUQkjqJwd
nyOBjEdfBp6VQI3ujX4GGs/22XLAFIzow7YSsD3v2NmFtNtrjzhp69emKfSl4xurykCqb5LToSGL
yWP/HqJNgNC6pRaKctvDgvZS1e+bA3sUcNkO97QGxMsLtLuxBKdlB1SJ9puzStIkzuXbKaBaU1Ru
J3vm0e1ijjI6sg+40RRerxwVcNSuICuy46MTI+39NEEQLnXj+lUjWJEDJBWJp01dtV7eqIJfOEQz
e9RxGt6uYYX/zsCqtzbD/3f0Lu/AyT/sebOk8l9/FDxkSdJci60sfh8IV4mcKnQJhXpAHl9TZspQ
1grCSn7s0vzwZqwa0ffPlD/xOTuxf4BgUUi0wlTJMGyuoGEaZcBGT/pq7S2yQN5Q018jEqKQSUxe
oKsYX+/QWZviE14J5of19AIDE/bBGIStI/u+X6bpynDe2SUnJipleWZdjqhtJUf8A3IMbqX3niwU
I3022UhZJvLYtpbeO6x+eEkdPM0GZXgSVfedNkgHC47FE2aiZutMGOX9yblnkXqeJajxxehjU1Lh
49aOYeA2ELnLUrX2pn9EIil9Zqw8cMUrlgyhImvQGUxyoj3leJhpjAayWjp7z/AaE0uir3jyyhdE
ykCTNuC4LdwGPaF+D2XwNFyl/fvjJosKWJAugcFX4cs0tROgpg3P+S/UvBJ1Eqx+gYtUe26wnBKF
uELCiLutzSzbKhf+idaNO7t8DDXFnf3gxSGHOMD57YtEZ8oDll60zea9ukaj1iJEz7ZjjwaRyDlC
r1igqFlhG1mkzzgtfa0odLDFgEuN4FWE+OJK83MkF69I7BV4ivnZU8BhhmhDv/WEDAk1O/naUEmb
BF8jUh5ZF/ruRrgrQab897Sc/KtmIWrX/igAkRKjViIBVD6ToTd7jjjPZJwNjdmOi+LaNTb3bwSX
t/OhKqInwFTdW78cSn1NCXnEPtpgKoF5eCa5V+PoeRDp2aR3NJUFhjRJqJbxZTXLcPWJQtBVCAoL
TOHpXYjYapsRl3/zQFkoHnnSyK65lHQ9b2WrHE9PQExmOrhMFOCkPAQ98DnDpm3yYq7KO5PW64ZN
nabZC6izBECTwLmSEc6xI+zpMAYfWvkqo5oIsCUdDeKWLSZktfQ1VgT7DzPH1kOsTN5xQW06Cq/Y
wkxHo2ZUJs1UDKY3D4If3UvkObTL2+0vZ8jGYGbaTkEI/Es9t5ubF3a9SbBfCrkdyFZbDdMjdHdZ
4ZtR2QHzI7Rf52DvLMtm2uvbyQik80Dst0R+i2mmX6sJOHWR0pMe69gQtiw3A8epkhON7GE1F9Kv
soqrkRziZnHp4wewlKeNl2ffPIrNIV7H3ITHayRc8oUfkNcYnPEP9M3KCnAYj9ZknygAd39PBLK2
FU7UvFRGb8EQjJfmTMVRqkVyWzOH/D0hA29eEnAesyqujTsSJgpdyD5wV3RvyCHOIpacj3hCwFL1
d4dcyLu5/clX20bX4Vx8lu+0+oHRlZ4bXVPPbCyaytbdWLfx/qpzVH95V2dVxQx2VlWYWbLDd+Wx
+vLfbmugric3+jBsKi+CZnRfCG3icG49mipQA+cR6iwylXefvWZoqs8qLt36RAMa+F6hO9KMlY/N
v8m1eT1BWFFjl4h46dev09qC3V4GYeWmBEucdVB5f0V9YzZutl8VW1NEq8LF8/FTWLj42xBoBVFJ
zGiJEIiVSTXmx8sXejYwozg+JuSW2Pf+G1zMqhf3dP5pPYqlEfsZZQTPmzsn+t7MEMB4DUAhOrmf
3S1HwneHCuL7L7kO8YVP2zpSuptqIylsMPdP1GjyFjTewpCpG4QP0Mb2aInD8cZG3+bB2+4x3Zid
OmC5lc87FWc2W7oNCqYsr9yBi4CD2n23OD1mjJCMVHQddsUAqKYgMQkeE+Drvic3oAAhmdgbpSbc
e3fXEeIcJlqD1ibs3i79XLveup9+e9P/e29g2ODx8kRowPZU1Qt4INgv4ypl7rTp/DmhqPy5jPM4
juB3HFYRQ8n29yzvTt5Rm4xwPcBj0/qbwVd+p+52RMnmICaN3yNnf2sVStK9SSpiZ5JqHe3i1nrV
Ety75ADSUDYaFjeW4xxOtIdTw/01fBHXSHsYrLQhPkvWa4M/i7tTGOePvNxRtUACr1/ITY+8jBtH
UNqWJN7t92VOC/1Ikhes7HqwW6kWJVeRfSwskgsGeQjZ5xReHuSyPKoIIH5RNKBVY37b0SC4NYrF
mpPEPsLcVpmK0mZ1jcnCYj52CB1gmE8U70q41glD9Q9iHsjBVVZPmkvnb2Nk1yHm3pNEq3AbJHmT
DzScCRqiSOp+/brxyvyAzyjCiFdY999CXOOvEDaIBnFGCWck8rFOB3i7v75GvefqUZ9rwT6vCI2M
EUk2F1FnxZzZwsr1/qwA8buQcC8fJ2Lo3SCDvPFmFY7/fHl2te5nWhnRugCcCEs/KbijLqFpy+0u
56pTkE25ztuHS+n2mEO6i7fFJ8BiYFF7e0/QFdBMfvCxUpO/oF+IodjUtdkc4dpr5eD5mq60plzI
J73+nD48I08MgxK6ct/PeppTfWuzJdw4zF68QtKJ6rY+2naKk6XQJPjhNy5oBjF+pt+xiuSStGaM
eFy7PxK+jUMVRuKDJ0ioh0goAYKAqrQfxLmhEQhlro4oaahzeDf7wa8E69ZL0dlMU3XF1Pk1Ec/O
MNQoJb4x55CbAH2ShK8x6ce0bduQL1IO9BmLVfF4gcCYEQ1z2j9NbqptwXU9zXUgptaYx75cBip/
ypuLo2JJ+buhLmJFTDbFkFY++6rvNwX2pS7bGS/9K7s8bqHR6BiH7Kkzcs2SQrCoK1oB0Y6BakOS
N/AuZryUDf/QWjkEXG7qPLobuK3lpa5dd98+wfz6NjvYzGweJNI7jMu0fnrYCBYsGQtrdoRKMY0y
55hHYj0w7gnNIqm9JFtDdDOnRxwyIC6z4IYJt4S0G/rr2jhbYwzTsHj70ObXvkKZzAvpee/7cQsD
zb/uZHpDSyYSJiyfmdMT544uJKCUCKc0ZFoeav0md+sZJXf17iRrBjDGCbNh0U6KLna1Jn/xLjcB
fVPLC/KP2jRsECf6lN2zG044EptLxcvr0wNT7ua2dMxd1Mxlw3vqmDMsE8OsjaXjptVl+d7PdZF4
EQQ40rvCphQyU+C6VsUWacFNcpTWTIqFJf9S4QJMmXihPtl8zzX584ry7ckGmeEbr5VZvgeooI79
g92+Q9y0+4BKT/KVX9yBevuNwHlO25IjEyvnjNr0MStCOAwUM50rIzkEjEEkdnHwG/ss3RU39nW4
xEEp0ar00JIOyNjHkCqNkKB1Zgtpyc6VptLRWmtH5n5rj3wpONN4U1rexomKbaAjxm28zO0Ldv5V
JFZgzvZqyfYMWx8m0RY3DEzobG95AzZYBR7NTiwHMxfterZ7qYMexsPKqrYGCYOXzobZITmLG8SA
tw==
`pragma protect end_protected

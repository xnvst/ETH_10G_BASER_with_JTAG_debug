// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:25 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BDPAGRNewUqVGVei7P0XmkDA0MqoH5mexCuakfzjijplX0FzZUgvnsRhsY2Z2lB+
Olco2N+xQ2FtrLZK21MzbDb6NYlqJjh8RCfxChrExzbExdYZuXBUuODy1isKELh3
RcIzJ+pmuEeutu4N0xxnnK6jVdZYtBil+XdP/C1jYag=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176912)
ar74Ln7NshyWVal8pMzuHbcD+cqRU9aHhZ6nI0VwiFhIdg6BpaA6cRK9cz2Qg1Kl
gwAQv1Ivo0Q8uCOfzJNtujJ/JK7Wi1cSeqRcmSSoSVnCp21gh6DkatmZCuX3NtwJ
xcjEe8MjY+qA2lDAEN5zSkEV+fsYvPueDg6g+YyqUKYLAELV3ljzUAqmf+lcj5oF
wjFPxIjbF7cS4CKsGb6+BG45AyYLepFakbCk3qjUpXJcTBUhOeLnaq9T3wcFkIp6
/7z5C2TagSoM3xs0ZVV3RG47oqIHWKjuQE5yOQGr56FSOa4tsQZm1NSETccn+AFS
/UjyMX3WXOeinuHMk2pjjxpEE0nK1FK261xMO7XM37uig+ZrCrxZFfnK8FY+WP0V
VeIISbXAtH+33ghBr/tGTX3A7zqqId9InvK1dGRZiIVvUJSprVeaShVpZyl+JiAQ
7dL5Ebni4PUVt8BcoX/sOUDc0aS5+sXmH3dJxh32QCeBF/6SoON+dMt9GO+MykAS
+WhTH7hyVfrik0txkmlAoY0kxAQ+c3MnxEK0ePdrA+rEyYXtQpyuTanyrvcKB84V
7xu8Ki9EF8Nu0q94To/2i7/7ExDLKyOmUQ61qI9+W4gFAku8FEduxC+d6CUbn2GL
VJC6B01LXitLJP2N1rcZKGT9vYWnqZcM3C9x8UlwrK6wRGyi8ifVJgDK+1+dvigO
9SqWXB9Y7fQ5w8qgVeECbp3T2cRBQXHLFNE4GLkC/DKKt3OeuXiOPz7+HW1NeHTX
wifCae3fHW6WtuhH6QhEzlC3eE2TXml4CYnFpjcBO+JXkE9wQesw0rX1WVOXbnDl
99Cu5cCzlBbTCzpOsHA4r5UxFRyvRXChOcQrDCIZku16fse1GziaUNRe5xvDKV1/
SybWJmgvn79DItx9Y/O3TjU6kGOY1fhCWKcdnEdQAuRkRsn2mV1E5Dv/tO0aZUzq
8guj8xbn0pzZb2gt7oXIX8uA82wmj6uhrTUpLEd/nJoZQBaAYILbswKYzuzy20MM
APgZ12ZNqOV1DGr3aHsx+vMi3/ECsE17jrk0CLrGOv7hF+5aSA8m+l52iDDboy7U
OI4Ns41+5z9RNQv2jUwacoJtdUKSLwFln6ozvI6MChEe/RSZtNS/HWaPhRa4DzeW
Cy1AekFotWDfsSAb3XTmfVB3q8rie7AlWIlb5Q0PPpf+Dr9kgwYAmTsr15oPQFs1
57Z4PyC6OH6ybS8xyb3QFgEyIzZpGk4HeiWxuEcLSxJiqhMksrFpfkQydOjMyz30
4TlZKxU1T3YKapXsM2QvrA5wJO3FX0LRj49t7bzvkEhFOwqZCXWBbV/DPyJ4JV3d
Xiw9XrkVCZ74wNoUdsVVQw9XP3VnO98k6SWPp4qGJoD5yIHCXVktEZIYH0IwNXbT
7LtZuXcSO851AlrH9RH3ybmGpSrjfQgpIVaz7t3xIMBXEzWXC8toRZ9YZwargTvC
d6pAod7kGRhUvcXpmrAPrqWgC4dZEn4eQ1oSUaejkuvxmq+o1W69p14cEDhaPbog
JV7Yw9AAqyqP1R1Yl3jIf3LpKEasqrzy8cEc04duNF3KfuiEmeQUXHvNq8wAHbuS
O2ilJAluywzXoRi2/5zQcVKqWNEoyt+6kyJN8r94VnyLy/xT/RTVBGsyX/kRkvSk
EUVmoG6CRCTVMC1pCYmigWYvnNqoDcK61CWaHRjtoaAhqyI5YqmF+MWSKXxP3KIm
HyaRgXdeWVL/yxkY0L4QS4HYyixpqbMo+GZUmaifIGzAZj81r+xS//SUcITTsbgC
7DiuxW80VkiCIWe9YsVYvYkNP/Z/lBkitCHYxsEyd9mUO4UqX/Ouj7uh3pJE3tgx
4REpvMvKoQ3gtPH8ohzrvI7TnIA8oS9SO8DN7lT57H73gR4hFTQRNfPMdjDCSJr8
pBWOmZkxRWWpjYuP2c3TvQvGYMmbmgofzLUt/Bh8G2U4MQLP/MWrd2LlWbcvKpm5
WseYpdaW7mmLe7N/jbPXhJY2clrV+XdtzzVmahf3Q7/AsM5X41Y5ykvVR8hPbRxP
fSyGqSoKKT9ZEoljlGlVt5i5gSjyf+gSsVljJUEkbVA5TpLS7T1L8+iv2jfNVcEF
p3OBA3mnvDdITygxygBd6a/hzMKb/Xc2RhIP2kJv9nlZdXAZ00c52vy4Gtcgy7Wt
KA7rsRcrrypJyYMUbZylqe1Iivp/iyCX8/dws6NMnGy7IAwfRlebHkM2eouftMdP
tTG34KriBd6PeMb9+AhtsZjbS325prKbPyetY2fcY6gP6h5GDdRFFihjkOvBY1h0
UjoS38yeNHD1gG8K/3yC85VAxPoe0x2KHtZC5P7hPnG21SyS4nEyHAStULt/QI6e
IYAIpbPRL8GcJ9W/RbdAEDzSvx3We7JuTIl8lgJQfeRCa6AwwqPxQGDLRfu/NGBl
Zn2RYt6BS02xKy6OvdcUBzbB3v+ppE/+DWAcWq0QoACBt6ExEUgv1/JXPWux3lu7
s+XVPaO8gGQTDmT7F/g3ZOs7eHhM58aa2/V/k1qz5u/uQroe6wLUu9MpQ+TNVuFF
ZEEhgKxM/tE1UZyMzolmwGhPd+dFv4YLHBGGY3iCyf1mL6h7PYv0DJdF8J1vMDdK
6uKnuEONONUSF0+xQ5SztorKb4bTe+EUI93eipHdTYnjaQzFPaQkmngxcDEIkE3A
JJ/CLaBs7G8gcFE3I/JjABFIJK5xfNd8JNgRM3S3UenavcY2mR2Pe9TeIcL6/K1O
9K5Au+L+aK9eSwBvmtC0pVQqTwaa9BhW9OS+4UKbYhuEJPbwkaTwxmojLPojRwSY
22xfhEThQZCzIh+OsWzZiKwwxq/WoNgLzsMf66mtqzNhL9XvWRIcG/FqazEswkB+
7mLGJiHvXFPO3soO5AMOB2EIZBcqoG8v5paeFqLx3nVShlVYvDQjpoV/UjUlV3Mi
8NNuWT18E55UVRs5EFivpOhSzB9s63sMwmG79Ge3nFqhcwyi91en5GjX3zWU4XTo
EDWdKVupQLXzPLuO22wHZj7GFc2OfHhi3D7/Ou0Oxoo/AC8KwYDF3VZKt4IIvJ4G
vc9GeP2iTgZyJcjhW1luvNHhQH17Ea3dv4RaISB2tXvFEBNKIDAv9sA9oq3hVvMX
CYoepFGGVHNBm/sO8ZopsABSWq1TqBMFTI6SukYqcGgMkidI1GdhK0P2FQyDaMzY
MEON/T0ZDV5XgSnNGB4Li5pWzm39OaLBONXac4KqeD18eBVOsORgJTe+qxRc7mZl
1fgBkeGehhEjKgTVbHaxPQI+DGis/yS6E2y48dUEg91hAHyjpZtzpGsp/CFEznoP
rGA4vEZ4ekojUxBhwp0zKepYy9zIpEu1uVhhRh/rzKEMthrFYzdbwfJcLj5ywIMb
9YfYEvBPuLxKjImSPy/ZrmsXsQgGdjwNuy8DVZg4hDY1efYFI+G8K/dIKI4aix6s
S6NkLo2f4CAgOn3j/zxF8qm3x5DhUcTE1gKx+2J1ywp69qQflpxCl78xjrfwBqk8
cpnUaP7px+wUe1CKf5oBJLDh1MPAZW38u25HUs9ruO5MBVB/EM0btVSqwQl4uMdK
4zYkDAA0g8RNJN8tAhCFmogYugYpAznqgcPyQUXTcdo9RkBL7scpeJuM1vD8k7Fg
QETFPom2S2X6ar5uTz91Z5lnU63WFBNnloVrS1TRiIoCDQ8QIt89zMhlv2+KVHAv
6dmQp1C371lP1RVzi35XjxCCh5tNPuwZwExrRrjWYpbcuOsPsCpz1M5VmotZfIIE
z4xgDs99ChVg0dk9spCCZ5mZqOkpXthZNvWDlaK9eHptl02mIJDlu1hj7j7Qrdey
bKl3zDn8yUqdTmDA1xZJ0mMsQrZZmyMdVEBVPndoVo3E6j2ufKFoJfTEcZOxu8wc
Oic78QaF5e1KWdrTedY6uelihvuWdiO/L5Sujfs2g65agVf+ANIWhbKhHwflMbK+
jEXhuC5cNHShV1DabCAvsrpKFr/J/1Oj7L04/PzWLjoiScFGx1I5w5HPFPlnDWfl
e0J/zypCf7XtAbjGzoenKIOj4MVKydZeAOHOrwp5LN/soR2jL3SwG94eeUzxWFEf
DuHuBjqASRAUDfiXVPWfjiMmzYpUmZPYX5qh07X7BKj/llxlue9FlbbCX+3xMGyV
fkFgIEp05hHxLimbYqW4GI+Xxx/HnxOEzQZyaz+sQE17g6F7Z1Dml7du8qbQpMxu
De8UiDNejb41TMXE4iV508NYTl96v2JU0wcpGx8BN2dzgmCmfWzWVJnZDkjpLax6
9tMz5G99A9Q8FIJtPmqYUp2VJOYDOVQ/wgxumKLcGV+xNOcOlEi812lm59r2K9Lj
Nh/WS7dnmD2gMFQqszGCWZyhAk40kl5TrpdhTl3PjzcVKkFIQ37t3MX1+Snq0kP1
nnhUpfeumOsGdo8lQmCvxI44Ojsrnz35QXHyBA8o9R4tO3E4/oGXy1HUAbh9x67l
epxMFLfdLR/J40nI53OmF2NmsCJ6rwTcPGxuVFH/XGCwZOiAjS5YfjvnBiRLWmt7
rZ4yCcWbZeHuzOEUVRjpYhe4EpO4vxvPT5uQ5MGljE+FOD9x0lnw9zFNpTr11rWK
erF6Z+Y9Bry0JGkcLRKWVYYMKp1ipUJvUhMpTMQXXSrNQbn4pQalRSRqNVfWRMVt
OFzpN9gEozidCxySh/4xEKb3MEju6ZUULHSANkxJXyEMtjry/onI0x1ZPa7hw9gH
dMvxlG4WjRUnh5eMFdQYgA3TlJ565vphmZfa4aQvxzs3qo25dZolwe2EE05NumJN
AvKFwgPsIXNtNouRc16J4pVG1RylrNfytHxd+oD4Pa89mqZJMivhROtqMgSihnEH
tEqmuaYd83lJMgR5EUCzWzEb+8nS5KK330Tw4tFOggVvAeBA50ICqyXtBNInUP8e
VS07T53UfDlpyQ1IiaXJnMqC7aB1BWqD+UfIuGD3mllJUK9xkjwLakrW54WCJp9C
KpGvPDU84CsV7DFwC2U5YefcGC+XEtm9xS+fouWoyEURkspYpV84GFuJlzablExW
XxObKSldsgCC1G1wNWI1dPoMT5i5umFLO48uHHKhav/MWamxy98dnLrwvtjD5VZ1
bRKAVPzHYOfq9ewxPUn+V0dCHU0LDFluSKDMA3LSoaJRbuXAtAo2F12Q07DtAZ7T
v93/wAvflLS7Ohzv9lmAJjecnCelq/+ZQrS2uS7niEmoOLSVvn8rLpK3u+9cMCO8
FTZzzD66H/Am1yL5UECTACe8JkF3pEDOdOddd7TMK5sqae1FX0T0DnFt0GjVzWcl
GktsIXQ46GoRc+WP90WeMoQX6ejD8pTpB6e2q9x+oMLflnVE04IEA8E0lG9/YyXK
XvydJsJF1JaL71QCVbq3wEjb1klpPGxbemrNL3eNl6FDjZwYrWvMGgPZLmzFVdNJ
YYqoIngGm6GVtpo9wZgpnsukni7ryFzEbIEN9pdPewc/AGHcYpA5NPViagVl0M6+
lCzMkw6dJd/COGLg1azlnBoedqVTdfuzYf6XdIduRy+aLmgX5MZzjQptcYuXWjDR
qi+3VeqPPIAx/1Sln/u3MdeBwEv4KKZzSE0XmsCHsxRV2/JotP0naQT22NZk29u9
IMsM92PLohU3C2wFEd+9pje9JqSfZEbX59ji8azaiwl2ifuP0TTmiwVMJ+gg1wYd
JiyKRrOdIHa0GOjg5WREXmfIasJVdXgrSztBGBubbUx3y+BD2ZgmPGBJ6XgqMbsr
b4/5kxgED5FCuRrcHz4sKIP6FWR21t6FVtfJ0zcpF/AICXEjPzIPVDVKVWL68D2w
eCTT63oOnSotuS/orRgFRrNLaXZvaZxPBOMDHB8HcPl+/aafpdHT30Y2+C7OCUox
XpDOXVE/UGeLRk+dRcu0AFO5yhXXLiFhCnsjAqE61bDOXkSxHNn80pMvZqUa9GEh
Ne0BJAebHoRKcVWGqtzOwvI9GzwKE9AY73+CKPP59AEej7lKdDEOxz+xmDo15FRx
3Oxsmi2bOVbAWzasStFTtbe1iWgejzi22AD+MoSD71+c4oKYf+2//38SLsXt6nDY
W1QJ1zLOWLMZ/7LkMsaS7tMFqnmmWwUf1/SvZcb5vVFEh62vQ1bv0rRKr3c250kS
t+HsRAfyf3/mwwt/XP7r92mPlqIi5dSr15aJl8hgLUHGsQXAFG5NXTBxT0kuikMr
qhwHA2zpwduUr+8xyaMUBOCxuzwjiVyCif47u2PjacXBjM9ioNVwkaDeN44TCxej
e1Obi3ZPK6Es+ju0phJLqattQG93pvvnJNyzfnszqUaZgnoMpZvpOc12NAWhJa1q
bnoC+Ji4r2VOOccbEzx0oOkQKE+VJS4SN8061gDmvjqrjniof81vejViV014JyQg
rcV4EBqGsSCZAn7FI3vFgSG3v4ZUsWf4UNks3PNvc5LlcCpgEqbvLj3O/Ec+T3fl
iaOwufuCaeXElmDxNczV8cYVNItliZ7VK1n4cAXau+L0pB2xSHjpsSymRf0u+7vN
K18EAkmWHNbvR2e0ncqio99eYMlmyMnegaNFwNFKEUheK5kgHrPHGcJIdEPXm1Sv
a3WVsqs2f+kgHGr7yWJ3Hw0Hd96a2H50RRKD+wY0PkinJqppni+x/Rn4WmolpnXJ
cE2AxuDW8FlAz/DwnIhH7FQSejEX63+Op5fx9FMIUAN/x2tiuyjfjKNyWdhQdUBc
usW3I04BzT8ygdYxt5WMwWfGHbhnAES5DiZKdbxbBlNHoS53LR/nrd2gnx0t+IMO
yuGnZplrYQ3xIBrlemawvBG04q0bAajQeJZSMd/xbOcxQmQojKoXvcoVFhf5a8Pj
dn9/dXUB/oF4ahR0RiAKx+g+wBeaoOu89WS4XqY+f4egJZklUMqgu756hMsf3uZO
1lcuwzcp0RwP9V+AZ3SsdpmeZxURbi3isObVFJ2aWJijf8bMwY6KrBlWILljqA+4
yanMGmJ4YEXY996m0P5KFXT++OSGhEV/U5kcSfzFulEasWZVuJh7XkT6uqddsJa6
DFDtSUzgdRWw8ZQCHeL83lUJpNpmVTA5fkG8gCIJbp1UCmJSxb8BlvwegZL1POpg
/tI/TOXelqh+tpf1oqOO07mIpAsxhPTjfxiX01MWnb6FBhBiYJQLWd0t5KCaxgXn
NdBZ+p2JyRSyInMlAtwqATYQenHXmiYy0XNcyJIR78sT7O8QWIG2T9JHOpPTEiY5
lL+lQcZkWI1JS4Y0GFNk6A9lJQnEGmxPEjF4eUMOv0jREBZERjvK8ba4T0IWapqF
bN/LOwbe8+xUzrwG1z6HlRq1+9kMFBOvfHJoOEWXm9WxWQSyoPslYpQEKng+kVNg
vcdy/R3kSp55CBcsxkclLwwYGDn5VIUgC77pGpsqaM6cULBjb0OO5vO6vqOTRRaO
5+43vptqkUPseXBZPxx6h6i2cVbeZoLPoGf51C3+IhIJzdAhXX0MZPTvkU0oM4Qu
4YhSMWkjN2ulK/rlFBe9TkE0ThYAKpsOuG6orkV0FVM3EC5HOpkz+DWRXZFa6S/q
2ayEmMMpNQ5D3WoEGwsY/zVl02JuaRjX0eSzuPLYpIA+es06rBfJeYkNRhLXhNO9
RTbpdmIMocaZsTOkJyHCyx0XbB6iN2DRY7wXetUwycC2dyJQxwEr1GiH7aWKvGRC
pr8fU3aFDTJBndSnWx3/NfHn0y4+hVzgcPphJ4L42jEljXCNBLFbff9IJac1d1IN
v8JBX4egkPubOMfIj4PkGOBNvr53NK+uqbDFOc6+WDLGEayCy3UFKLr+ZsLiSXeA
4YTkXNE07r9ZgXberT1mc7kwps+s4pEo1V2Bssg1ApZi2QuH5fc9ZNjZp2+FWADY
QtqPUSQU6PNg3Afc68bPYH59nlph2No8lXFtqFspDsegqvpdTlUED4IHUEVjs1r8
xwTY279wweTauWVoNkIFneKSLshDTbm0cFpPLp0iYz9Jl809heR6NTADNna2HSIF
prGbncCigJk45RfhOKVz2QGWTrExp6GAsLeRIo5X1QcoGRo+vnjaBc3lu0nK3M8k
KKbYrVwOvjdJBVvTLkfdLX54GC3ZgqMbdGeaFh3Fe6NupRDoSpzVaNnMPgj8ftDy
1V4OJ6464CDLEz7QxtZsfY3OJ6WHUj9GbIWmlvj4Crci/oZ6TgNU1gLhFUQUVGKR
g32/g3ZyE1iWcnjVezaV7kCK/ZbGLPUYBnQZdqayjZdyoLuZ0wrdGsGZvfYQ8kRi
7oJZ/qsYGJxLLjWZJAJyNurkY2GyoXvflLdoamQJuA16RgFk0Ui/cfhtFenaGVVm
HsSqICOfi7CuO7YrMOfUPmBh4xaDEL8SXi4MH7vDmgWFjVwKroWGJv26DooQn7pe
gUX8SgZOQauM1wbqFGH66OxdJpkAIWin9aq4STVqdQQlJpTq0n3mEAI6F+AbpbCM
GL3ZOCikdZzFFNTYzrbwJBGQtDA6om2WIE4FcGiFktt8EQTxVgNHqwOOfkrM6A1o
x6BKsBKxBPzeGvpjfY1k8Y0w+CdAXry3sozHRd1TeLjbKOq5r/tQ+B6e6B/lUPZa
lC4FY9RLzbq1pPAWpArFNtQgwtyjWto7r4zmOqjme+hz5qXf5VAaRjn8UzUZiJUh
JzPE4cwoddJWmTZoNcVTDfav4F2XCEYmHnMQDUarVx8PosZNG5c63mWDWvLkjbEC
5gz736ehIPMC47vk9UqTXuNLfMZxqaDg3Lc4mBT2duEOJoe67E7HahRFp/3k7XMM
DfLK2zjtu6xmLa/XB3o/NUt1bBPtigRoIL1sN3xy54bARbHoRgSs27Ct3p2RdhWz
1dObJ129EB3S6pxqPfwMWXvpEDZg8Du74oszi+1RyIczics1BFcdq5wa1t5YEbNq
n/kUpKhPc6AsUnG9xq35uywFqF8GRB6D19Xp7mj0XyiDCDPXEXetIZrgFrsyS9Wy
kNYE1/nQ8IDxpCJFQ6SkFmV2pb+y5TwIZnCM50H/uq6D7CXzPoXW4w6aeGFIuKhq
axvq8t+OyxmFYZFsbFdKDUrIA5RnTYeALyQGWqBJ9VcgmJKl0I1G0eNulcfMjpvp
2uzaQajlKFJT24ANonMZHCE7UEL/vuAdBlyMWdTbNRf1mvSuS4uijEITeiXoJXru
YTitTSU6NRzF89gHpJMxbMvsFxl8QHo6gj7Plbbo4cJWT+yA7ytTKo6Tz01zJTZl
h0EUZlRQvOV0nqc3P11rrlaJpi7w8SUgs4VCvnoDuPWrPxBkMSPEDTd4FLvtpKYl
Sg00LxS7YNplNliFS2Vf9BRcYtKBV5h+PgVjOee1LZVs60V7phAZqx7XI/5Plsrm
BXyxX8xLa5M3gt1WledwMb/SAHHZBAIpsLIXo66v7KUPeX3bWkPURrNjPeQ6gKnF
slZhQYMuyeP7MSKUvsz5oKaR0XLCc1WwQCHmQbScIuHP3yYXUD+mtQPQi/mUFckt
JCzG6PFkTOVLWwq8X7z2I+7xC1uhI83gKZrExQDC3omgb7um0n6HRqCIT5sgXS/b
zJ3KVjEIvVX16MebYP9kcQ9Lf9/h+n1bvZv5Cnd/qKKdO4IzP9j2GfKsxZKxTfs6
Wr/zP7DN77XvQKhM06HZD6gY5k/liDbGZqgi57DSRD+egiRoasvytHCqJVDm1ZDv
peYPFsbgZXpNDvv1C09FkxaXHgWpF4yVj1Bw1CN+OTRPmfUkFOHwYHGBl4y4LPR2
IZ6VrWXPy3i1Bshf81yCjajOvZxk+fboa1EDhRO3+d8MxN5t58d/8EydlznZ6Ema
B7imoBV61GguABje6GaXBKScRhT3Zxw6qqVD2lnThqoEqeEI6r5vE9nI3FRCl2Zs
gx0Hbs7zKBibkHq4+0eMFT++VkGzy6sayZKzgKDFAIsMNyuVekXtTn7M0Ltn7hiS
QPUo+6qf1ECE2qDsWII3d8lcjdwOM33SxItreSUtL7IHl6SHJZ+YZjjhG4kgy9YQ
JzcjchikHAFnVdJ8+b35Hy+AmNRqiA1D0JAPEhtVrkNA3niVj/dpiIKpSTpi+uba
3XD0zeIwZF3KgZJf2BSjXtCn9HpbyGOih3hmv/vmXJCGPMLMDXWc9ruZ5a7vOT1h
UdAxdEfi/2bwA4KNI7bEGBE8suSWvnhRXTrMGn9aSDC9LGglrwktVQMgcaE/dRfB
SZ7/p5J8U2zSup4sWWKZpl7HpeuNuq52ePiHT/i98703XsQDih3LUIpFORdd7Nwe
RafxBrRSZTcBX66U8nC2IX6lQT5ZQIBcUgWvtuIuEIKieLZ6BOip9rPfeFLuPfDe
yEn2dVe4vMhupvKVGk8y+pILwTLRfRBWgtSIhgdHDUTMINYKeigy0JUzDwss+yhn
h2z0Un/Q+6lVFfjg/SnuYYWHihNWE2Sswi1IE+2674CVn3QacQ3JO9lRQUnmfP+i
S0/KhSZpMPAAdZQMZsk6JP2+Ic7nWmqc9RTofUxZpvTQW6jCNCYPFy6dhhwK08yt
pwm0A93Bzsn4iPJldJIloSGW0MsnnKXxC705fPwxk4A6j1yibLzRlCQFFtpdIVef
+HIVeLdEVfQXkcb1bk3I8GCpG2CieHd4pnP6n6mZ5q77HnGzQG9vbHTB3wWz7HNU
m180AMauKD0ApuIUmzOZNzMCVESjV4tn/3n6hsEeaMXzHcHG9iTzwvNbmhBu3Aoz
wbhllxg/AseIUj4SF+I4XWPW3ZQj5yxJ0QMARO6rb1ExyWJ8mdbq7ABR531IN4iQ
+7BQZGQVB7PeCEucdkt82jmuRSEmtDsG0ZhJKPcCcXz5Pzxix5FEAcL6rh97CN8U
jMk7mr3fxGeMYrLrWEmgCZ17z8v9GcQkwXH47X5ukbvzmWae+MCKDWvRqi6i21iX
SHh811m5wZpoGXA0S5jtBMiaA7k2lAVZ2T9IK8kZ7ghNWdX8EYGl7+cCjy0eIqDG
nhAAfGwokNGtJRt98hO+YS99vIs3aOkcEY8hUAj+vTPe+FQANWFqvFnbrcv4wjky
xbWgZ3d82z9X0bTvKUbvHQw2q1u1lRPVRq0MOqCcsPWwchNLXOAWepy1HYLwG7YW
bCvtX3iwDVD08JLEiWoS4VWnW5o+du2ErPNWahgJvCl6R+u3vAgjmBGKCzQcyJzQ
FSfVJwGTAxCr7tEgW5wlEwIu+4UW35jl4gWDnWabo6qMAMPbdyczvhdvhGO2Ry65
DL4Fv3+1sd4hufJU3KcICYbw1m80HLx8Ahp2yutUyXnj67YK/6If8Gm97hTYGGa9
HuDvACkRjMe677LAyBE6UyPKlI5D5VoUDDU9XMFfz72Vv4KhblWYPKFvBIcESrRg
UYjsBikwOIbr9A9rZqrO8ro6WEfwYkX7WeA0PPSM1Hx+Km6qZ3dIQ4vNrn0AUK9u
0FJKGMX/iJ1vEueEGxoB4inqHkot0tLAZEvBcWEPdgkfF8mC9ve9F+ILCqN1O/zH
UWH/1TdUEqpRQRHlt2uGjRB33to6auHBiKRMnq64dERohBWKJV0qzlNH1k3IcPl6
UyX1FO83MOCFMysDkRaRnol4ZNw0u2dxQnTdsW7WiW3eDOjHcMfQ36dvXsUkydT5
hmBoeOorAbO2nK93TtGtHZbKGHfdksEUxu57IAuz6d6FKdBuO5x6DATPqXUh41L5
SWLki0vuoVRmPPFCNJQA7K+NXCJNtYJk+QvvmJMXv8Zup8VsM6WGsrKqS+37ybzG
qMZFzydS1EmJBDFuCSmrFwSUpfCnGIVKGK2Ptsok1lQ/iRWw2KSKQyfGg4ibDgOj
UL6aLq5TGYFMY5pKCPGZSZ6sV2+YJgm4NMQQQnOPCaJ6SF4gft9Vu3d8URCoS5bt
SB0/121kzdxawzXbHwqC1Ncz7IE6N0+w8DQAG0ozNaH0UQ+gieGJ92LHmQGvtFuz
6AatsNpC744IeMpJWj5gatcplFGkeLh22MgGhd8/KH8oCtRkAqqSBNwUVn74bIOm
ItImUOFC0VCT5b3JqYxXDopos0baBOGdM4+lQbjny8KtN6a/y5pQj/TEKxfd4awI
X1FDzqKfbKDnrlNaYBUGpE8+orfNK9Hf88TPzUvgfTtF8HePd3ZoaT1TYmg1kcIM
R7TiGpT7l9E+BEK6WY4U9nG4gU/3dt/xQo6OGk9rXasbDzNnTFEY1ZymSxdI2Ijp
ZJHkh7iLpBFJnHLNU9r5VqGL28p/Dd3PhCPSXYr1W64ra7IO4zFbpFvsyIPB9i01
fbevuZdjZqjLrghbhQhBzcG7liceDIv+Yv6fxUbPM9S1fh6W2CKwIfMdh/WgCxeg
uCgCJBr67MCwbUMCCCNKBGXGZ5P+T2oU14RheqLFcNyAStdWDMoCcTcZeLN+RO+X
4kXwvI/re1zYLLBlA+QdsIpuDJWu0ZONTsA22R6fm5CcQMIhCzWE3hUaLT/znfYr
QUzKEMLEaytNYXnBwUUKobO4MPRvDmBPWkh9fRtcNXOB2LfM6Sm0aQA+OFlKKXKg
W6YLR7ZLpCtzqzelpV+r8yNhQODduK1nr8d2IqW1C1eBpbkTfETGvpCnWQyUcQkP
VyQ/dMB9vsvGkiYfUC/CSEOmlCNZdyDdlkQvRR35Jm56eYbg8xIWb9xOV86+8G16
WnpgFLZUS2/XAWBflXgyQHzmVeRm2eZTnmrCLShOMw2eYvnhT2aDyGWG1dW8thdg
gP2l9btMzq3XPmXCp4lU0XvpZPDZqDZSjbgqtr1996dgGL+YZJrwfZT/6qsb8UI1
031QAt4NLmBONyX3WmHDrxrTwNDnOTnFdGZalXeCuuEn3uQYGQNnnnR7dMofE9Be
NfENL4tTyQ4iB2M1ephOV1tE65FexSqcRt5LZlaD52iJOVp+twO3p1Bv+Yel2MKU
AdZwSCn/nmsEOJj+Hn0RYzeqL72kCZUx7HdFkfcQGplsVPC2G+DzZ6YGyG7/Kwm9
AtDm9ALbysyYeHoTT5JEXr6TNEp7D2e8wfm+Xl+4DVLagNL+K3XyrNyBuMDyQTPu
/op6Y/CI2uZo/zNf+z0Redy4rwgz6aEgVNG0puL1fOZDrSppZoL7pjATORriyoqd
Ac3fLAs8XJOlOYLeMkJAQ1x3JWoJoR8Va8JvSSeaj9qlYvDNCCIk4uaISENsAx6+
C4ECQIkgIUWyojraDDi+3ZR9mnH394SltwyenI29X93C5xhtcpHqLqo8Q/+zeXKd
yX98DIQ7JO+8glH0udPBIxs97jBUa5nqTwbTH36E30TK2/auhPtfFROP1mmuhWvP
z/YVUD7xL9TymqMdA+w0y8iJIusHsq8FbKBnvxxi1ia/Md3aaDvRKSXvvhky/ktg
8dwXhV+72entqIHrt/Hoa60fdutv0OAsyvOOkLA83W1VUBfJF3ItXRLlbvEmhltw
K24iXfKl7u7Bp+kb1hxjZgH0dNcwEJ+8i1QSUY4aOIbAt5A57NJF+AATXrjCv+Gn
VJwPMRp28Q2JIBBZEIIvuauiwSfsu82sP1iZkK7fprxwriEDGcaW7+yBLnu6afqf
PI/0kbeE7gc9/j/LbwOEHXWVAre6J0bFqaz5YToW59xrzz113hh5zXCwmpmBrPj7
Mm3JaSMNn0wxmSNsxJlWvz2fiLfxvAIoJnSq4fML7TCWLqIqQLlocV6cMyGMEjF2
KIRuw1DX29/nhl9e00sXkrCyZFLJVV6sUKs+jnnLBRMjAndPtfqwxjXxTAX3nIta
39DqWzEJSLbXigF6UHRGLKtsPxawMPTvuW3o8O6xoMp1xlnkVjiF1QLXk7pfzKdT
zMk2OreQm0s2bq6ZfTjmRzwgI+SadWS1WfkDXknfuqawRJ+zU7evinE1hwz8RVUj
VHTm6LR3Ce5Asr0KWHEI/y4vK4ZfgIZi6Y61Fetj2zeLcVav+FzjLSCx5bOKvXuo
8LFCiHxgITaQtNDbmZDZTa5kXBzrsW4KhrbXISybnilKr38+6xOLn4RbxqYXGLuw
DDhyytn+nVAU+UAK0qMd0YtKmDE3SwaFO22pJiLH3dUBnnq2mqHaZkv0sBZ4aEej
Z8jTbsvjHH4l5c+MKJV93/EDYv4bqPDbC7Bdz0vTdHAAD0ku8jtOUU9nPz9CTt1i
n/WWaWZ8oZeOIPJdhiMSeATA1M2fBkRGUHEfkD7SHZmV4tjAgdSZBmBSyBbZ6eAJ
3zTdaJqUpVl50PSZeYfLQxdUJwbPYAcEQtTufe31aEkqg48clHW/a7gjpXrfSVZU
EZT/QAWfFycZGsYqo+GIhKhpawNSKpe1Vuw2eTWOxCX5wxwbfYVy3bekkI7m2Qpx
Um6wCGS3YfQypMo5DwhoNHRB0nejaQn/LkrXFWhr/KB+5dR0cFQk6BeuG5NAMjD+
mHedQCCAmSJcO8mWJryvJVIxXLI2kqvgbCCGbuc7PjDOxZXJAz9IbjwiKuBBht6x
Cov5RgUyXQrDb8V1VObhyEYx428g0GrXkv4wvQuT3TmqTHGCurvmHVaUNHj9r8ZU
N0PiTIU7leQCSJgRGOwpN7cTPa2vf8/zSnsgCtTkKkRtprIe/z8CTNIkXddZ2iVw
3uvqYn++IKLoznBP4MWqzD6yqdHpKAXqwgOzHH+PXzdZBSN/6ysqLb0x5SS7htT5
w4VtO2cgkKKShDpJmv3/+6AnR4TvgJDy4pP3o5A/jcYITuBXSY6lg9ZqTY0samRi
M0kv3c/yd/Z9igS/wZxtRyC6F0uvm49XzrUo7bkclA4pvk2quc5iHU2RAYg6S+x3
0BpaQ2eJQTXwlcH7ZtZcZTbKn79mnciZ7Yw3f6zR8N3TKQanzN++u6JBa941nIdC
KQCT5fnVUctD2WfjC3y2ajDpTIeTW+j1oL2NnRlacbdRZIQkHx6t7BQGtbe2ECXV
hQdb6IkVkblclBlZF9lwFrncYxyJZMbfr2zfU8OfxkiK8A8iAE3S1ywiehlp8Yiy
hSslLMIa1E6o+Awkf+r0YmZQA2g/s64atHqafdgVB7rnmVpDOJatmqSOE4ACN/ne
VDZjvbsV299+gVgn5HR5nlPBA6NYPP411xpIunUi39Md7nvKgEcmkXSVBw2sMmQh
HHpVvYyutcZpYMPtkQbXVAfS5fY6v4lj2pfAXcBSCz0qM+VvHyE5LqnITdQFXCEf
FeGPmF8gn1z6ha3iorvTdN4ceYVuCfcEMRsjF3x4EXr2/a4q3gancGmlV+/WlE1K
MAX+L+wLQlfH3VN/7xZxkHrQZMDJTxPVsSGjmBHXN4ZC407Rd5I7vLVm5eMOA9l3
I5Nx0/N9CSAeXoh/sZJhMPHVVz0CxcnvoAehLXZyO167gnTvtsoipOQ9zHsDSTsw
nHjU98R435zH/aX8FwZz/c+7yFHCS9N3IradoIliYtIkftaMEn/rIzBStZE0rdS+
361pEUbf+lQbw66EiXwRR7yLeUe+9/E2dSPstIug7HumaauOaqn7c3ecTUNVyIoY
n4947i2XkjXfKnMNFLK1ng3Ao6D6BCfoa3Cs1j7z2MDy7UzUGzajkjudK+dnv48X
AZ+y5alXNGcAJMQB4kP3HxlMf+WoyuOsm6I9VFh1is4DakxtcMlHYdGVBCbBQ2mU
QIqvQkpN1ukasSDQenJdCCZbU6g9af6f+uNWCmFF5Wt/y9xA1MC9ikVo1+0hjoJJ
47EkK15E00jSsall2l+CHaSBvr1UtuA1LnHLszmbzWwQ6Cn1mkj3UWCIK8/lBKLR
yC3F+utf2NNKuTnvpa7HX1kjDvLX1eLeRaj9KM8u6VjGBqLfx1y8zrxa3rt9u1oi
9Int3nYD3NFHIkZTdySiZ05IAqHE6J7XZFABzguTB6sQ11Gcbry/wG5h31jqvVKz
n5GIAYZf41NM68y26gSW9eqx6iwFb4NkZNg4o/a6c5MpyXUlACxcQEBtmdWQlbEZ
y4JsECbZq39voXKkbQIwT1CCrreC+k6l+0SM1UGIB1ysbJ9cbBNA+SEcg7rBNE/B
kroSSuV8up6ZEJUN63bEkfSqajHUDV3bpHShDEfhWowxxjXErjWaQEz1Iv+dBnDZ
ue25SScDELqcwp1P4VVr8BTJ0gl0x1tZ0uWmT/wmDNTeudnOuiDUors4Hd9sU+sp
sbjfvcLYY6HO7MwO5jRVeXHey3SwufsvXkEv26TLJWjBdOA8WWzakRd6nW0zOK3Y
GFQX54usfNBsDb0jWgyKgJOs2sn+5uwbkfww7j6qoHjcOgV5WEOhbevKmJ37RNyn
Wo/m4FI6H4oIRG5GrM0x78wJNRCwOym1eeb0q7VUyV5GTsTQx/qDMo0JijMyWoF6
Xg/BbSJXYwOz9abaPsJgBbgaUPnGFbY/lOCv8+Z/a6Y+QW2FitcRtK2jr3IyeGLK
BM20Hl0QMXFZColCiTi4BwVb3YxHJB1U57U4hRNFcfdRJOeKnesCX2L6sRfd8Oyr
oKo8WG8PPbaAtDyv0IwS4siPMJayntRzU0lH5hy/ziCFHIGFYkkfYVUYIqZt/R54
hLHS6BFBJfH4p0/6vkDGIZ3Zl1hbNu6CsHI1JZEHZrIia9Td3iPb+Zpta468X0aM
3sKTQWAYR9DHAYQ93p0LGFA0fcGcytAHedrkqPzrHSU79BmDrYHzsnAquIHw7WZw
hd4RPiMFW53pne8rUHIxrbUN9AHAVxnsfIqQbiS2phF7OHgUZvIWEA+uopza1CXM
a/jlx4h/TUDs+NPx3noUrMphGJ4pAhrqHkifwm8Ir4thtshP5aUbMWDdOSVYxVEa
5Cv9jQ+GsYG7X1GbOXrvwNFf/xHxZEhLehicHFy4zBN8D+KW04873Xtia+6K9b3l
rdMHu3RKQogUzN3nTlbkvewg9rbKOkphpWf7/yABPUFjDfrXaQB0SM64q/6PhWgI
8TtGGWfPWaKzF0DWOTvHfzydAoap057Wavx0tlp3UM78SIoy8285om+stv/mEJ32
n6aj/81/jLqZkJk5b40nBiVgeBv1197aM97exj/tEbUkwS1cBIF2YL2RdKM5QyXy
n3EjD+msUsVwX6zXwKLqtQ/n12pMJaW/g/MaHjcb1XPd9y1uPZLdu4gHbSyVmTIJ
TvZxsW5pbDB+ozbIQCmzkOVVpVldbzoBjzQPEAlIpAxczCpO4jSv/ock9HVJIduV
QQ/MVZeF08wkbmNzRMorcIwrzENZLaKyxP9Z0c1NrUZ3+88mJaYdcTdFrd6Y8S/v
LU2uNxd/OXYR6J1Ag3JPcKvpFdXZaORcgqMgyXfnaQQ3oHPh7fi1B3gcLbBrCAGs
qAC0e2S5KuXwAjQ+vSGrlMki1l4fm+3dj0V9bW3ypWbcgqmNnWy1TQV5A0QW8eOb
KEnzYhSOO5fkLuuQP5F2bi1YvQUjNmS5F8EqXpm2L+Sn6t2vIZsZywt09+Fa1xuV
+AewQjSEsOR+nDLJqWGtX9Ghsdq+i03RFL78UFEupr5K/E41rtKOh67ZquEekpRS
5ZNNH9+LeqzQftZTzuTfXl4niDl063nrFTpme7RC/qunluDTjFCKDFQSDMYDD0CK
5KuD9RKums3U4pXmY+ECKfg4+a9NxrCZrulDYPQvtktlFsQ13C9XDdbWrmurWtAw
PhExZS/xSOztV8Kud72WJOyx2HBSXqIsyjGvY1sjF2p7LcgOxXdfuPrOeSUR+YWV
GmGTLy4cFu1a/6w63ONrSo11PbaejbMO1cvFLC0RQecYfBVzRLWyk4gpr4JWUom/
Xp6UXzxOP68CDCIeQpKWvtyuxJZwT6sGJeOHnU1qqV7pmRo/OnwkxKC8RAjSxlw4
zDEZLYxtrdWic5PDXp6yIfnJOVymGtR5Pk54dEBg8+kwhhFIMVdAVByl45AORBXZ
KUY87qLBvXS+4zrLOJmlVUZm9GFerspafTYFDq0l3ZTIMI1NHGqsAcMIYOg+zUaN
5vZTGnYcAp3pxzAUNslbsnh0z0a4Sw9VG29gvPj+j+52phQENn3tOK8vqRwSXMFt
A8278q7x7aBQIr8pEaglyPlg8/4EbpqFLhxFeXfjkCWgJ/yQFNT1jVL75ih6WdKG
7DAg+1SxD2r9wd2zzFIcgtOhOwmt0hsd9so1K1IgDjdWGFoTy2bRF3kRL1jhX+E4
b2saTmMg7GrTyNXldhGPJVv34MBAjIggIrFH99N1U37JRa2xcQWbOUHAu/wwtsyc
ONYBLtLlZ6N+n9WS6QKBwzFVAKvMlxR9nABotI6RKqvuxDPByy0SUmMgbljJCvKy
3MAz7badQxqXiK7Im1p9msai2cnsIeweV3eIZxBXOZvhMs0vie1dE5iuGmyxyr5L
JN+o1OO2zUa1zoiGUXzUqLHxiDr3lBn6Uj8teQeZXUO8piZ45DyOEFOBbFMKbU2c
MWhisQMtvfCoYZIjcJRQNWK+qGrXvCBPF+K1DKe8+NzhT0KDkGS52C8pUOuP6KCJ
1nUm+B7Uc++qz+icNRGuJbqNfjBSNVtE7UExT0FNcF3fz644KRuUqZ0ZvIb3BIgi
g793VXHtavHqL5/uTS/W/MOsNR9SjT1g1WqxlBXqGB2ekHwYK/C0lCFp9B5LXIJH
QQM/le/gaUPTsc2FkIGK43j23nytbWTuR6c9929zGzIZKy+F/8WwVsCMTpn+7ccI
DP3SkrPIsNGFUJaeTVyWRXT06Pc0hIdBQM5ymypgrJwQm2c70xH7fn2p5Dh49S3k
FfIDaP9mxekqx8Gyg2Z7Pwo301ngt5wmP5rfaKqkyRkdlKn9JT0+6V6NY8S4lKJl
4wGPUZfSLtMQiiuZhln2XtaVz8KCiG/1DN9ELKajpkKMgKKFfHYiEudyLvDuqbLv
MBrCad6mIUzDJQYfMrvumk9xoI0/P/EGX5rkeJCiuGttMrS2W+KhROjt2vI66zKp
Ki10lHt7Xz2sDoynordWKjkJ+p0J2pEQ/wLpn4qauvxME9xlRpjjaL76k3HC2hEq
kV02wEgBfZul1YixWAHbLKSZ1yLHNev0xVxGcZ0o6unexp3UG7QzAgfmD5sCKDEs
1zjlLS9tP6/YZjxKzHvDKBNaoYQVZbfHto2hXXGfR/Wj35dIB05CPjAbBAr37T3g
X7lTiXTimKDMPQSgCCta5Ff1bzuHktjL4JuIzaIbZ2K3WU1b6cIZro9Ni7GaGVKi
QXfnU4xVTNNiek2L1r1xpaAEIkRjNwEZNTolVhxxYKFg+rjEK4OEqYlW9SqWeBLp
YMMFSWGFjLlgAid7XdUkXGhomY3YXIdUoy1V2esKulyYezEY7d+zwIXq1S6TzAAH
jXfiYSK3dtzkvz4WTZvRuE8ukFRozkKsLMigwfyLQDS+kSH7SJf/c3YPVQJ6CKI+
VFAiMJxuF92VVjHlH7Qltir+SYftlFAZ9q7snh8wXhr2ggSEXNZzVdaLQfGBrt/m
KbfIiTyEGfpNp4iyigIefxH476xnGS1MTxLVnB4e5SKaEioCSxR3eD4b8QN2debw
TL0y8SsHigfDKS9vh2oshjMNgmNAep/9zuQPplk0E2fZ6/AVieQApuAEf1ss63PW
STtxJkSFD91KCvcdHF4pCzbK74uSmt069puyR9vX0k7hJfnaktt7jTDnOhvPS3gE
wTCqESqQwKoaKyn4SnFXTYq0FYCpjRwpcYbLBIWtQAYO+lfcdPrVowQ9bJkeE6Mz
Dy8wu3CMWzgOwyFaQujhxwcDgUJAFOScPYSdRt4V8tor7UxMNhEDDZQ0gSYqzHWp
0lcE3QRIgc45svESx+5Kr/Y4rjNZadlFTeh/e9+H4pjdSAD9ULF4bMGvQ+oRp25G
NMvqcw5/l1ofsjOqyQdkHg2xSa86gbIrS67eM+1xCccweh3NNN+H1i5FJv4HlIvE
cENWM9wSgYtDhffB4nV9In4kdhruHt+XMJugjP8gXwAxIWpaieEb4kHpvdrJAlQP
o/0+0B9/81Hr7+OBYC6bZ7M0CdzYPVKiVe87tLXzw0vTIZDLmxBEcRLm0//mkRco
InndDt6WCHDrkSVcSlCMJHtBRUETWj5LrLib7iZdembnIjdrbwvgXMXEOfkDOxCa
M86IenW/P73Bw5eZBCvZ0BEAJOnYtIgCsZVSqJDYLzxc9k4tuhrh8SUE+3lxifBE
1e7Xc0xCMAa0hmQ0Ax5IDef/yf+DkETMV9F9IS4z1Uc4aSqiseq7uyAmq1isuGa+
qmCEymlyku4jLogqLtYDYGaU7JfkUo5iP4sJH79n67HN0ONd+9FVjuVvBsLPwkpS
+/4toWmZaZjNCe/PQ6szbT5JV54GW0y1dUHPv37opjwwhPjj2k59D2PLATj0Jt8Y
Wdm3yhccqJUO/rxwzSUsPrn6ZvRMKCDU4jO1RI3qPZGEob1CJ1w74wNi3K+Bo1Lw
m0IVAUsF8xVMusNq/YIEql4+DIus9L2BcA9RWXxVVCiv+g7LbL2kqY058SL5KPow
zkil3fuuA1sF0+I2QzqzvDxXkEkv+WtTMcscZNPydvT7/XdZTugValJXYCPs6wXM
jI1lrjBUZ4U9jtbmflOmpc/62j7DEWLyGaCIxKcsQUvup/SyikEjhYoNMRLegeOi
qk0BZtkmkZF9vhXdNTJ2NSWIdZCT1nHCvrJrr0eUNgC7wnAv6YKV+ftTkVsBbFRN
j/FkoVqN0CjK9EXCbF2A9snBouOq1qUhg6qcDF6KdrpjBUlc+uSGMaBoUNeyh3lz
RfY6bSslboS6/xdzdXPUCpdwt7dnAxdI6SyoNpc7En60hDZZTy/esfL484ibqc1u
35DwfxMSLV3CTy2WQOwQVNtmuKoynTuBnJp1Wx3k5KGyL7l3wcDemFxj0E/qvkPI
QcAw2hzCkZbtcA3EPR2mkJw/MeEjzK8fghb8nqlCOPiXb8K3AwmadNm6YxxNF0Lp
T4AVWdFl/QuIxLTNHfbKiJlUBYUjXou4cjyPXXfsDTDybLjY7Nnsh5AZJtZ9Ezfy
XXEpkRPpYqU1WVNQ9Uv4fYyOmO3OCabpIdqyYRVgHDIwDFRqCWIVzDrlnCs3Mayd
ts4aNLZLC29dkcuBTvp8uw383l+F1yR2Ep2caLziLtOFqF7xBzSxaJrGnpIEIrqP
Xcf18XTcqeRhQKx54RVEpXX5lDQPMn3d4ufBzcNrNY9K4G7Y6ytYjFf7eGJGFEBi
rHocFkGmlVntwRICKMzMPkcIObA8Sab0I39tuAPoVJTZBlrj0Ck7pEPH8yeR11L3
0d2A69V56C975AIGorzuUHBXQVsVY4P+xqjDBuJ2PFUGT+3KEgAahvmu0iyrPF17
sRQsU8PVB+wi7VVyrwSZVIzsgQnBc6Bu3WvEUeHgFnHxxd9XqB5+Ok+RIDXQVYaF
7TsZElCm7V56YfKQpV7Yn9H3D/scNDX+uXP7iYHXDE+nmnDqdyJzaM4PDeKQfbh/
ZOK8HQm9oxCIJMN+uWbiSMhXgWiFcoGPDL1qK9gpYcd9o5CS4TIcTq2ZE0ioUQL1
YN6YBsZdsPVQ131t04dwPWY0j8LJ/2F4I+TEFsGfBsBoWjEvFn2S8B1xLUtzbSYO
7tlOp5820h7kFKV1MFYybpvZjQ5+yh2dnp+ArJt/9oDTGvOgAUxGQbaOwA6uyLPc
NLTW+puT5+O0JAADKlpGuTpzSquFvaz0XPHtAQ7JOayewmNXf2uRx3aeKZcOV28m
fshze31+ElzKtYlseI429KkLuzOe5kp+9nfeiEE9xRAawhlBcrQeUnlZ7rRVEXgJ
KGw9il7GuuUmYCG5pefcf2GiRS8JiCa3Hy5ULvYI3N6gGJOojsMjWyASg8l4yYfi
x00Qp6dr2BoefXHGsm54WxAH2+W3xsDTRXrtqpm342oUTSvnAU0Swu0C/L4R5pyV
Nrih8S7ZVJSfkwCsmwy+5EtpQRW3RS18SqxPMz7Zl1vXPzhaAruDcGCl1gqLcD18
N1x2CBQ6/IoTkqjx9EzCnyXa2gRLmMazt6tUMCC4qgmXBWm1lvS+cRS0QY/DCjgd
ArVp06DKdp71IbZPbMMZ9EO87n84yIXhqWf0VwMa3n8yqxvhpyEBKepmdpi45g5l
nxX9mleM7azopNc2Byar/N7LRix/hly6pQUXtRpPk5NrSXRJlxRZFdvG/tdygf9Y
Bscm+YvhyD/HnusPjTYxZAqrfsqDs8zTIhq7jIYEutkO68EnbI8lYOzEv83Sqqqc
5dkmtSiGBsgcojbpy6ofY4031mFbMx6Lvcdk6rr8wKeaWw48qxeQO5ClRIEVYOuz
Y14BhVZ03WAARipApB7JJsDUf8QTFVP8jORbmumYgWHumD+jWsR8FrLyEeeEX+3M
mAAjGEssCWAz6w6BJUtNTJH9E2KSTXBGZ2eYQ5bN7/VoW3581CBbUXLKkS63XybA
pbHZy8/imA6P/f5BwqFrHjwnlLC+amj3w2d+lTvlTIHS9U6oGDNU1+RhJxbhkBwM
Ib1gpBQA70nKHY0umMQKDWYRDH197h6yEiynPLPO75kcjOX38/l6BJOE/qSELUCJ
8dNEtOCxWDiFaCb6ZILD5RmgQY3YhZbmaZZnAY0Cd84CHsO+qt5rpBqfTefmhfl4
jaLeH0sUwWlA1pVUlqmVyGS7cTdOMxtVUNyYXktWYhiT19RyVodu/TqHd9lwcerT
i2CjGC5TYsVTjnAcw4fAtc/e77tkRixEGzggDjKlx4EnqCd1KYquTYVLuKn2ty0y
mAByfbLq4kYD44yyVwPVhqqHcE9LsewHSxMRJsAmfwcGJS94PMaicF5kdtVPIqF2
VFwNy0t8xQpTXCKJR+7LX253CMPgP78yXF8LqHpspE7a1fYp+X3pyRNH5GiRDR+L
tKsRwRAIa7MZhWdu716wAmBQlaUtwYTglxBgMA2IzGgsjkxeweXwdJqMRZS8jupQ
0KUyokUqW7jgEhXTN8H4T8Tz1/ijvPOw1YxlaNXB3AL3afvovo7M47oU4eN41DK+
BVIhncl0y+TdOPPNv+lC6nko8EBxwSzgVP8zEoqXsIZg7pe+fo6bXPHnIPLcaARa
Nq6WlkcMd4rjjD49mzyxA+5J8nTNjgC5EOdl7yWNjdtYAXr9LpAmeXoC7rN1KO/q
J40vSFUPqLd5GutVZ/e5imyNIfTH3xEAVxkZqCNYtqSx3/tqIFZGjMHBnX4gzZ9p
SD6CrHyEkNpZLgSmRxOwgqF8gaTwhtPRqrLDF53fL+oGuvWjbw2TLG/0w1LZfAD5
kDQoT5R9XJ7sNwQx9K7OsSlLTGBBewVh2P6BtKQshrYs6UzQVXSS9XJKhb+HUZFR
WQoQ8tdoEYWOOLxZiAqZLh3lblna2JpRj1AC6Y5t7TqWDPe5pBQIwFs80VKIwEGl
6jjTKdkMY5p5dy4Kv8yy2Q/axi/58yJ9EVFM9gwVvTrW1a8zkIEauGaXSJrO26W8
7YmNGJkK/DpeNhg1OWSdq63nUISXwln3k5tsSO7PWkF4gFcEXJM0uCLYv+/jMWF9
eEXpwMWS9o1dfXg/NlGjnJAgQ6eGFx18tsvPOn9uu/5hczW3sl8cFBLtQbbSPwoW
OJds9xUo+yOCpz8DkMi6MNfQQCT73tv3U8g2z9pNecdLpjNDkTTjjXtrOb2HcHF+
/t+/LbZb0WBDzGtGumb1gS8mdo6Us54LPo+UEFJmNVVQIj62T38iFdPDyQ1r0g7j
VqrxuKhhbmVIc+A6C2owFQ8HPjDyaWbkEOL3NOafQCnGnnAuoisj4U7wPfYBF9oe
wRpY8CRfo0wcPeFhWwAy4EtmZvgHV4svcWDqMEAcWK0UcUJ0FNzk499y3lnO+EAN
HspDPlzo+J6X9xG3IzFZfvhQtO2xsSooVA2VgbBdxOf5dWFtk6WPMzF9emW4b+Zi
V1eRlDxgDju3OJp62ygmiyJFdTCXPpwrZEsaDDbanUOFV3/YhgRM8Hg0ap5LtvTq
5xJOzdFC3fi/86PpXT1dzW+hhVcbSCex7WNPGS2u4CewwP0wrV1mO/fByzQ6T8Ln
On5aYrcAQEbjtg8L3vuT08mGOW20Q4BjN9TX2lpyrTUZR65bkn4fFibcOIHBT0cg
dU2OfKjRVEsnBqrkO64GSalm3oNlQw6w4xvpJw/Kcd/nNek0w4bDZVtfZuuAFg/2
nL4n8byu4nOCLohxzxb9+leW5/nnPHvp5nsilcbhE9K8+zCGFIfjKhI36lbCBU3j
+AgBVaqQIVl/u9X8TaQgOsJuu/PJiZaL6QwRYh5XLfkOrc+NGlaFCXipIfWZaaT+
85I6jHks84koCxHdmV5mIhzTJLOc2KMKhYq94x/+W+8KKjjyUdn0aufJ34D8J6xQ
N7A+JlBde2iqVA8A/3QgQZ+sajElj+TTjn1HYrR6dE0Uz01oUchpFq6zGv9o/xmC
ER9l6gpDTREl/00eWBPLIm/CqVfkC9uzsiimcmE/QAwbAkzqSD+b5U2kCznga+v9
FIi9wBfmuNbs5abWDjgHWzDQ3iY5r9ngfsgJkY4ya0nLbbR+/t5bOp58vz52ewzz
umATfSiNgd7vQ2/+NtqzM7F6acTwdJBn10ehKG7aRW58UDUa88AIgLul8y26tQRj
IK8ESzaXFQZlIoGeHCHxuTS2xfQjhHj5R8xGSMj5OlDkG34oWpOSyHpQmRh9bgTi
5i5bWFV8oYzCcRYlwTlbHGqdSILckmQJO6pW8WmvOECCFhWjOmSKNHa3OM1x9rJo
nLEAlYSBR248XaQCyjEnPYlm/e9McE6tB3fnolDyaNCMCuPMQs2H2W7tQsY64kkU
yu2in31mdMRuu+PuIpfGWMs+Nh/cY2NYDek6UL0/D+HOOTB5qvuJa714F/wB5z0M
xedS1DXsI9HUYZ7CfvVMIDgza5SOJNB80yZEJizqlCdgeWuKCTWvfM6yAKPXlGQc
DRQ2GsJS+u6W9jjJlEYZ9rUTMsuNibXoMQ7NYLMYepB7DaK9c4QwRvqrkrUy70bk
UcPMuXAFn7Su77NwIuv9CLVI89pJ6iOAMIhiiURiBUCuqEfx9FVCv6eiNaAIWLgv
xLTjlPexW1UZ71cyHegX/jZDF61LIhEaCOjXNke2ymPqzhz17eWSB6Q1D08AkDU9
nHkKYQdhjoBmy7qQhXXTBEGmbH/gOVf09O1i37deAYPyfZO4s0NE6a3xC69dWx9k
jm9cGOqXJSq4pPdh2JuPXIV0C6BGLCf31GPDU1BRoVim9ZSIXIqN/4+4wEmEJtZ3
z0X2DdP+2l9JZXrAz4Sa2Peb0IRwwoABRkM2LEcjPYyqNFE4UEtNoEy5TLjfGZSf
o/JYxQkseLFPmkTlKa+OHD6Z3ajIldGbiKO7CNmrlxytW2NMknWL4GkBexOqced+
ZZH5vWePVyf/F7tNy3zI1CS1aTPPWWOYfBERMnLxxegan56OsEQJsLrLY+8HASYw
y2Ac1TiwqtkC+NiUpVcB5MYr6NIoofIpUIlvP9eb5H3xrgx/3weDlZRx3o8UkT+G
uT5ykm3JO6Ho90gekJo9gjhYBx+WB90sT2rRWVw83QE32+CHM4bCvdZGQ3rQmaFQ
DIEc6AUCy/E9ZzsYJcCalVm0VlnFc+4HN5ZKK2OvBFybkrXbb1FpAFSAxrGBZait
kD61RNolV0nJ0KpkCf63UxHMW1i18aquXAHSkmVpVMAhE+UzIuqteFmY7IsfwjpC
t/ZwFCEKp0EXECS0+6f6qDW0T6mLdCq8Gx+i1/1F4sBszlJ5jQIvvuOKG+NQpe9N
BHhmeLRR2FUTHi6HCxyhGRWJ/Dkiy8p3PsaouKRJCSVtV48PqJXJLMTKh+lqCTBI
c5KAH0HtSAYN3vUIXvJdxY9ExHrXGFOoJCo37xpzbRJm1VWXiC7dweIujW5EzzRx
OyVqC9UOjTNRm7K/gtvjG0Nei/+4P6RPwQub+iKAZfD3W3OyU0bbHXaxya5FgqJ/
jGs7/VRi2fsLQSxlhbmqAeHUKdohh2+U6WAn8e8+bgxAypphrTf2FW1lYnouKnbb
psXgEZb6xvhqbHcbwCgocAv7koH+CKGmJZKSVmRt+/y7EwzpmoKh4954ShDsT3fv
uAmsQWTDvnWqvPahTepKvoOiQb4hT48FOieiIIdVa3HRpUnDuC+4hqUgC8M30+FS
LjXpkOEgEFDbWg+O6liotsBC+R/zfRauG3q0SrBxwtftN1gWt7Cuu/yQAPE5Rfy2
WF2nludsb1hoNwmFS/n0aNifkfUlmraVb5pKRjpP6+cFp/OyuqGhzDRw9xQAjY0m
0am6FulYlYm9lWLsfGqxrzkzHZp+UmGbZglJT3g2jEtOIIyF+MdHNC8mOv4Q2Rer
K2PgLQyp4pSqLgjdygUvrQZXHEIhbdNNX7isiDfH7H4oOV7X0AtoiVTpeckXHmKI
JIFuV5GgoyFXabMas1j2f8EoKxAw6jp4y6tT7aVg8CFM8FybFVILfar1LpFG5FbT
0vkmsHiOr+xO39OS70nJ2L58Z28Y5lvpAeZRQx9DqvDCj7FKAEBWcYrdPd8L0Ci/
ZyqH7QN9PJYwavcxLRxAS8m23ZlPbiI1JyrWkZvSLJr4y9pGX4Z2A8mdAOwC13J7
WNLgChqgQ7GcN0sXg+KfBFZM8A0bwP1xjmW1NvXSo2chzh80vm+PWUU8T+NMUSaD
II4jm3DTCsTRECULhzOu89L/xqHrlFkgIVnPR0maJPsqNFQX0AhK8P6VKuX2r03k
G42N/Dzc3Gduw/u9Zf/0/hHYjWteSW/rgqhF0OiCTvBSqY9Q4BMyakJlCCJQM9Am
N/sJ97YgJ1a1jONJIaT1CqnAJG8KoHRiXdMynBiZDfLZqvxa7uDNrrSz927xMkno
mWEalGFlyNpdKF0V6KWBuRQxIS4wwrnuUBMCDB3H+ElFJUeBGuPGF00dRDXFAwQs
j24OqS7W1sE9XPKhVDcrfXcDoCOwEmOH+f+tbxKf9JfvZcXguC1+QDAEckpiPpzR
hERKa0cQrp9qlgFQvUUBqPLOIhA+7uepmcoBWKzWgQQLsy8rsxj9nW7rIbvLlg60
7W/Idx9EJhxK8giLLxQUpZQM+A3qbjOj6Spk5q85OiRxmFTt8pDgUcaMwy4yq9GL
8NaZsP6A5Fl5yQirN2dieXvcX32xB++b+B+Vr2btQ1v7VkoqIYY38j+8KDhTtnD2
o0oXhNzNuWnD+I2/dJJ4uL2MbfrAMSYkilCT+1ie2CJtXy7ZuMDLpUIHzjmGdkem
Vu58f5Pfp8iNSaYX1/KhHAoEWN99D7wzTlbrducebDSrGOC0D3RYu2oOC9jxJBuP
nzCmAsK2Qz9OBPIqkEMK61Y6hFzrWk6gJSoSNirJh2Wehn4lB0dQow0ehLkGKKXw
/yyumO1BBMqfu0iKuUHj0cD/A/28TOtyLBIWmbGCeCjBOgyW5gKwKtvMpsLAes7I
d1Iu5FAO0AFUwWWvhSmxHoJMn9BYgzD8y1g7CFJwLO/oKsjubbalMBqIvf599r+9
LSPNBToK7UtWUG1m9zMt7a8NW54FsBEt3BajpO1Q64+aSwgqOO1xZyEXnNokYoa0
i21uu4trFKM4SQBXP0uybs5E4bRYaAS1OXgpVZQnaCYi5rn8rdwKEdZGPh8u5UBT
e+yoQSM373w/DIiJYKAVQ6gpmudvdVZ8ja+LFMnW/EhNlIvqjqHU0SCZ0nStgpbF
r8qpmxIgBHVWTb3ndCkD+r+SNuvywKW1mRlyms726jEch3CDEDU+EY1vtWzIxlO+
mHq7u3aVT77XBpZGWdhbPj73EZ9V7p01WFvpPp1Pa0VYyPC6CZ63s6YSvSuFc2Ma
a2ZYTGi5EqkMjowPtAxaJ7oniwsmJ0+qyPLiTuQ8vOtjGyb3d+uwKUZ9yYpVXlXp
HZ9BApWW4uA/mJg/kxsDjfxedd5t58udyQWyKLWjOBwkdPXJPFd34148URcF0x6k
cwP8GgHtvAOZNjWlin7rYQFAmZOsDf8pteTAxlEX6DuTElIko5eeSqyM9I7Rq17U
+Va/scf+C5oBb+AE7cNsgGE29uDPLFl1ohd9sAQvQA4fywu4IYa/kvXXO3A4mKEG
FGBmIrUCu6A/a88XdmvVpCXWKuGNdBvF7yRCFbbvUg6gmAGWrSFhHw9y/VIEwX+R
64LfUespbWPtLLvfkc7EviIS3If7Qmx9Jv1gRU/AP+H+z/y0xf7gsWjr8gHsN2r3
4KBQYAu5XBvBY6WCzcjGhwoukSxJQnGevPpzqQXVjvhmMQYTs2TuUBSGPpBLoJky
T2nemfv0yBXeXA/m84WfD7GTtZOQrrmDDNvoYtB5XOaM4aOyyM8GXVoznjS3D/5d
0W1LnEahLvAj03isLyuTBmQzFdpFcJkLXNihFGczo+p1ABy3PdoW7wpoGyw9yPFc
0KfzRutMfpapAnrIkIm07sEQYKOS6KbSqEetBVgTE5rZ/uK/hM4y9h3z9lY0ycpu
7+7xALuFmbe9bvlKEswGoGe43YMuySlvEMVNz04sFiLyISp+T5zkJUndNtkgzpB8
OocVoyjQrQMQ4ezLp7jQjSaslOLV8lVL80vj7l9lpg8BMT5uBsEDkyK75UGBf2OB
3GpFl4KhG+icqx59jiqKUSUekECoKhILfbRV6VU8J0zZsheTj09N5drUTPFl+rTE
V16OYiX6hmzaX+yra1VENSbwj71v8wPrv3MIm8Oh6Kd5j2E9MobpdMR5KZw3Z47E
0qWgGk2roayXHo+dJZVfUM0O53kxqi4WRaPd+2o1D2Kno3q0AEIuVcj/1QrNZVj5
pFirhQmx3a4fROPXR/Pvkk2lfcSlZ3RKSGXJSpSMAqZZBDAzbDM0YaHN2gOth9+I
LaVjssN2j6BlOLposE00+7XFX29j7Rn2BPtWPYhi3T9OtO/+Mn+dFw89kKxiwXpi
F5GQHbURFZteeLEKdK5uG+iXMg++NTpOxEJnritrU3xJLw8uNZ/lcPZn5pr/etNB
rSeCFjSFBCKhx7Lt0NyZ3t2EDczaCVlxKu4HQ6Q0LWoARlJ+5i9yym9UYQJjIANF
lMsJJ9T3My7tXXeuW16DMMCmkSKVcx6SLXgfsQxD8M7ftVjMlb2i51E0XTYewaGC
k6alybdPaN6+EA9DzbdXU2I8hbemn0tSis5e38ity3DuHMuzr0aGuxgpz7ebZ8o4
8lFftBBahWsMNDFkCC4w7/c4bV+BurF/lXcTqeS6FzekmEH0O6oDmdXh5W32IWSd
GXuG//gyMRptGjfkJrYs6rV5Xr4hQdc5ISyUFHisuyWLWNaQ8FmzYZb8Iau5Lgia
KPDvSsnCzYnVQGO+cv0jPEpCx0wRk2eGPFXN/z08VgJ+2KwZYljiWZ1lbkyZjCXY
MwYmeSx0pD5JzFCI2soNpNK/PRtY5dMkZvKc4H0BkE+SIbVe/pM1Kts9P7c5NPCD
+ibbOd2k2CkqH9mBq7oTgMuf6wiHE+mG093F70uD4qN/0H3NZc0VWExYGMYMPb/K
3TYHmV20f+sWZ7Yk55WyGrLInauM2KJtuArvKQ8CDE0gOLVov2o7Y6Hv9fxQVukg
RDQwhf7dcyrRRC2mltxVtQsnpsrZXlkP6Op9DvS1kN63DEXW3zUxUfHUXiOZ/VX2
RG9ynEEsoiDJCptq57+vpsRpyty5Zo5XlYI1SmWtN+NopYu1zwz5rEJVXJrvEiIe
DAs3Y9Ifv/U1grA1B1cU1oGJXM1N9zox/1zYTE5kHSiThj8jhEbqsdi7zKxvU2v7
DIFXbxqc/llU/CbkF4tRapfZ6fsR5wU1dVHS0FM0QpzRmgv7/5iHAQe+KfwODro/
odDrAOmO05iLMRjqObMIoZB2kCyUjoT+JfKAoTnfIb6QybBqYCedbbpeVCcXWj9e
fHwq/iuqTAvklLP4tVaHqaasTELb4V8sCeMqpZPLRItoqXfMLHNLgPjUuilT+Axw
59uSDHXBbL7TY4XCkCkFyUij/R6GmGHxeZ7e2sKzIyK+/N2EMj9qrR12N0V5bAQU
3/+EtWm6ninu5a4cunTTQnUabjcFF0diHxalFCwEsimuCoXm+pES8tQtQt2hxZMz
NdcP6gOYt0+rLsQrXWcfC291ELKJuJbHv5+78x551dLB5KyzE1Cc1pWaORzuZmOM
EBq8kdYdCKSQCQ5uIkMhApLfoJijl8jICVa0iJJNkqzHd2/zOjjCrziM1NKcD8hQ
tbNF0kd4I7PkpcNUf0Eexxgm0OjE/MOEVDDnUSDZdrhUrqj+l1MZXrdEodF/8Grx
a6tIjoYDsyGrRXyofcOUYV3d6HTYChHPKWZuQq039fc8rFNFqbCaknAOq4XZQ6i8
j4JtVsvxb1n/JpVEZgsPaZztJHb+S3H8JP0M3jWyvFWaD4K2BUBRsv6ZEnkn9iz2
woSOqkAgK/JA/0bh04UZT2X1YW0XKBc65M4wozSAdUY8rYxfH22/SazEbVG5cYP1
AZ9RdHM7wDGg9Cd6tgKO9JsYK7G6wsmbndcqWbAdKYXlsgivKHygbwPKZnOwXZKi
5hL/0EYMqI+THUo5vTLaTvskurRinjkYbInUNyNRolj8iJV4B5dcubzm9dfzqcVa
hwvG9foR0KwxBUbaXOFb3fyUcOLeMfmNeVl9gizX1B7Xkdjt0XITVzAFYejRpC2I
bo8JzB5N289LJByw3pT8qUvwcPNaupxv5+1y5vNJMpODPQSON8MfVmdSPyipmBLS
kvPAqQgwIvdqFDG1Xa7yoFprkvo8RTPhG8HsEep/Tb9IR5smlSJrTLKC4vEy7sx0
FaaRYqPSFbt3sVYFgX12Ivr0RC2vB5bl53tA6zni+sMCH9nldXPE9m/PO2qRexMt
tCzyaZZaxcbERP2M8KTtEr3yWJSXWZWkTQgMwEnbi/SdZUGtnObVFqZxJcjIj69V
Et1+Xqzbiozc6iFG94OFsD6rVgksCffCCcaQlc07JJpLhMCsabbOleIRKhjHjqoJ
5R+du0C8KwBPtY+5UimMqs0fmyzcS18eyPCjGQD5XYnODY/aR8xLYnv/Q2syvKuF
7Su3Sw//cOogaStd6GQEzA5MquwklnCPpad8p92KwlNckjpP0aLWyp+RnxLJ5udL
b9aPYOAzH2l0jirJi2OLaWop8LW6ltff4nSOkNoEtnTGGbpFjn25XkftLn7PHlHs
E3oLRREVUI3iRPPMNig4pl6lvO0mLnLdDIM6JHQ9BVLqgby2EZVF5zeLg1UVRv2C
x/5Mx0IVUhmMEysOXuf7BmnWJMeUPhXct4nj4XocNe1neLlFDXz+l16LNbZv5GOU
3TJwoehntb1dlekyxJECqmTJOHHkhbZM34PSySK6oWqX3eswDjfLv0KFjXB9BNdw
2MY9XxjFmWZoglUVigckavWCjaGsnPQ4IGLG4oRhPbTv+sxUpHll4dP5XxJBx1Vp
bnkmWqpwIXrH+h68+Bfj9mTlz/Lzwpk85/B8F57zM4PQYoMfNk/cbHunICHaoZf1
ib9aKI6B0FDDHQ7P/2zi//g+cvoc2VoH60Zn1xEQU3OJZgXZuJm4uSD6tr3yndC1
8LMMpLZWdgEdXWtKvsC0SYimxt67JN4FwFZ/Eh6Kw4SbI1bwdX6fsvNxPvXZlkXP
AbjFMSYndxZ3lWL13TmgA0P3xDGLo2o0de7z4RmRkapU1fUoVxX5mejQL1neqHuL
g6/tQsc4v98OkI5WYiQwKmN2hxsn5Rx1CVIk1qY7/SStW/TdAMNTXTurC9eMfn3B
IG3uuT3U5zb/gft5LEfzJ/ozGK4pks8OzJj9x3ZT6vb7/gOkOyXqiJ2YzDR4dBly
md/MefCQ+5/BOQ5JMttBMyvlkm2uPMD0w9dasRzCc7SOxzFMHCEyEUFkA9EVutmq
IpYlvV0f1SybmUCzH9C+A336Ae9Iwkwov4mu2FuHC/JDY+MUGodmUiUDKteDeoTH
7sMhYLUKJ+cAQzlp5qjY0SZCI2pZoA81bXzM4bCX22OBL9zpbdjBRvqkNzTxOCvH
fDiACM0uORnpaWppugUj4QyfZNSmw5V2A07VtG4lEkXG7AdHyEJjiRoQflchprOG
AUKwuHVzmzRzHAQxaKByao+BObmUqSOwJI6u3PCTUEsMuM2dy4XcMH/z4Q+HRmEc
mxX/T5C4dZcAKAximWErMMt2C59QTzWhkhY73RHk7v+pM6iMFgTZdI6v20lO4fTI
4+BUGoIo6nz7xvgBJpD8WejQzcvqFeffVUFx/1vVhvMUoCq9+Y5yWve1rzO0DFv+
COkWCivSi0Go5vMMRrPY8ycsqLdNJi5MAlyTN6lEQsF7HwfoQgVGAUckl+VLn8iN
aKGZB+1dqTTJ3eC5TtvatSNGLTVB7N3gyJUC8Mk1gYN+YKJQ9F59a6mClXpTHSOI
/5bfzj88NV2ulU4y2LTh/LXgPp0NTMCcksE+Ozw8ErTbL294fkDdbJHnGmmpv4cP
vjyZ5blbT5SRVmhByVkH091FRpF1p+Nj6aki5F8prpJ9z+9Q2IqWc0GlbuELXF/3
fuzbdpj5YzkkVcnTRDrEq0+q2AO8m+6SpOnALCTrcjEup3ertlvL0rp9BZYApzrO
L24gilcRpfM87tTbVZJBW1KLa5XG8DvmUMCEpRSgBP5ZK2HNN7B53jKeXWlFvA9J
q/icYnRI/lRd0DglOrgyZX+XVNTafBHdB3FiCGcNMgRkCa2/7wQSOFL5VGq04D23
qZqb6jcORhl4mfNEgC6Xvt6qHc/uprPjgo9tffCVYWsI/+SVXCsz4wmeGEoua0Pc
Fibzg6FwZi5isa4hWyCZ45J9QWte/dA0EShwyEgeXNZFwnyTgzgBaPzv48y5Koat
toMVo1g4R46zn/d1Pzjc/ao4ZXumbjW38595/YQiWOfFBZn7wWbY9w5U2+kacfPU
y3EUCzwNQ2I4dpaIuvP7fo7bmYQzKipKvFxQld+DMqsRJ6VoOXD2NPJFqWWTsQBS
kAu6kaagttbRdpZSXRcEeV9UPtBR8Jqpk0QXXeBPlfBDjCQnFHcs3OpyH69NkXaX
ySk7ehQIZAFOUVUp8ZqZNfWOEsvixWYP6uZpNUrv/bJQYXzJfBxVQCAc/cdUXLUC
8Vicd+9tUjRAmr0Rsr9seQI8S2vjOhMdKO7Fcs+6QiYNO6lr9vX/i3Vg0+SR3ucR
TOp0/IAOYivnj1fwFjVk7okuhJ2Cn/wp1lFLA8XwMwvt6v1eHe/JN6Z0Od7OFfgm
c3zsPumQGQNj6+jhi33XQjByVLqfRaMGZBMImxpqx5gsVHu4ME5DS+DOHetXtqvc
jnEhsF6Q3h7QUKxMYPSVz65iYifZcqy00BqoCRnaajBWIX978WwhqKP/bhho7ClT
hXd1Mn9G3OSv+S1Pnm/rqPm+38sxM4lfq6AzWe/66ronRKZRTuSAXwLzedjRKsr5
NzXEGb6KdhaKhO8hXaX3UPizkVazOAJlaXMnvCrCuIAGDFDcY+LlanOU+P6ryX90
dAfV43MfJ37dCKjAd6VzeYoGx2gFfw6em9eoemcC1Fbx/tAYJX8iXm5+20gQA9/Y
GCksD7dT+ko6E9+RxumbEf1/5v1l0Txl5dlay0FhtDxHBm+I24ARD1LzfIXuvGOm
3y6ELVliWO+KsUEf/pboAdrW54GEDhkZ92rz5dVMNP6BlBbFn5k12viigITcGmtY
vBlAryN2X1n45zb7wnJtIKDOoJ+m0+8w3UOkTj1jr0eHaR77noef16EyucJd9/+y
b9bh2y5mgLd2cUqyVkz4L5bkRj7DFK1omDj3z7HVGgvc4EPfc1VC3LBQGfT9Xuk2
l/+HuRcy0nA2XWtD1fjeRM49xtfDo1HWsK6xdrJenAwLpLQzI3DTwc4rxLb6bFKu
o0sgy2RyY3GSiEdoCZqdTHkL2yYeQcQwrCHOvCZHDl5YZMZ4nDzBtdqdXkYT5RgH
QXR/nb41JUeA005X82GEcrC1zdYp9z1QTE3RyUKSr5pCi4Ijqi2YycfLiPYi7abY
SfVApbMkBbUFTQIYyGD0X2KS7951elEG7VmiuHAWVbCosW0fug68TYvwWSYjzDuz
yZKYdrkcWQnaChHu1QMNaYQRa2EnUkJZFQgqJBCwjPlfwmVMQVwwx4iEqCx6/TPQ
cvvari7Of7fYCnMpYQAG+SZJTiRiFJYk1nOsIruWyVp631ydsBKdU1+7cIbTiERK
77F1f0PRo/O8Oue7ZzmKEt1MWKYgR2TyEtzSxJZ7/S2CYJBh9J/5vWGCV/qJEmgL
oQB4WkGxEqQukxAzPM765XhGCV8rfb45Q+mFrRWEtG4BJJCge9ZUuHpmP8Sly66Y
QIb2T3rKJeqg/gbbZ6Qk9WVoR44bw0YqQW1UZ5ddovOek27WpIs4Iu5SFRENi5Wd
KOX4Yma4iieEIxJnqp8V9LBxEuch8zUleM1dD3dxhKWEIxTLM9lbX7dymq0Zx3IH
bExNX19j56/PHTEBsUrE1Mwye/uqHGmy9f17HyJBf1scfDX3OJf2rsH6K7faoRUS
NpeQE5g5UkR3c4q6o4b+OmBf4qK8yjUvnC3ZyiK2XPfLNI3+JO4LH7mngGz6k25H
f24vzgesCxAlbDiCErf6u+cYDnaG0WUK/ObXXUPz0UNkByzJoxSkhDZ40RSSsVgd
rj3PciW11wqs7EMtHoC/4Nsrn0QyePqq2zTYVbuB3ficB68I00dL8+A1D0UFMAUv
w+ocDZdJPpUG4XqK12JeoM/F34JraNfEAQomQQn8ROvLWy0oQ5doQJHoDcAm8zZ9
uf/KzGKvbrwqTAPTdizeXbXSt8dWsZl1UUbFG+/+QpQvdaF7YUgsgc+2LtaFvj1f
r+xhTnwgRIDfAKzxAQphB4jTjiwpO2CMhZ3LIZK4tTusqiP+xPBJmL7RA02axl/i
fe312Y3CkwwadcOwws5DEktGwybygRkdZjdbjYgxg1sJ/zoYDdHJU92RXfyiqzJA
nq19tUj2FN1b89m51V1YoLEkiT0JmwFKZ1eDJvv34T5wputTp8NRyd/M34loWX/C
x+jl+B4qlZ+OICdmHjDxAqP5ZSCnJ+Qmk9/+wgyOl5tOTq3jMj0exbIPzeoAVUE1
y1WFRPuJXoCEspN8fp1bA0abcIHxmH4yqqz2V57p6xsaVDglhksJA9tfY7Sz8xdM
/H4YNWTO3b60oqCpYigwGas+Ygt7vJI/iCgZ583kuXQ1y65ev/dyL94KZF1vCA09
systdVXbgQ+rqaa5kTQdlPa5CtuIkTIGrtMas377tANcN++bGQo83XnG8x2XKNxy
igjJqRlgFNSgDyHR4EDiXA/0NNSieqYGsb/llqcTA6jEZXSrtgMXSwEwTD+FaeOn
tsSf2+O83tIzGV+burxaXJitqbd5G8NdHU+QLpMk9hkPkQF2P2ynkCimgjBzXcmb
0WJGhG/nvsnwJE704dX7I+BFuZkOOhptdDNAULS6oQ7FquvCJXhdXDlnJn/3oBQQ
umYDBnwbebmgkYjle+tz5++qYN4s3IXAVjo/uqJf2jwjFbzW28qbpsZZwRfxFp6o
EscF9ZuwEVeqi9oPAjDdRbVaNfatn0LWseaJMsA0bo+MHj9Cx2EN2qC/gSQYL/0a
VXTFStdEKAGBKeajSASiiqDeJI82bz++cEvKAbS60kI2s4x3I5EyP8XL0HUsH6xQ
R3AgrHsvWSuPmxdCLN+FAqbZIyNlUDSONannXNiYsnF0SqyyUj3hZgb8wGkgDtLZ
gdE51ILOzRdXzaRioyL3Th7trgtorgnwjK+zKhprGpuItMziDUNaarrwsH+RzoiV
vX1Iz1Dz3EwYuiIaUS3QlowZQ/QrDHsMvgO7QQES4cRi7pi+eCKL4CJzZZFhBy6Z
nA/GBUc/W1WCnh+xztMnegrwMkaubZCB3kHF2MnT1ejYszhnsMyv+B82FugJo1ij
7QbyqhZ6mzmQUFWgTXVPtGKDLyJqIZO3Rq6LO6Bg19S/6gDt4UI48WHhclA8agwI
eF3xUFRxvlKKDVSkHKlfE1Gd/OjJzbrqzKj1dN9WVPjqm1d5KLzh3uGEqYdfgFD3
+Bf1r8rMrRhWKAzLwJnqr1VePD62Zd2dCMwWnYsXc2GzEt6oOr5wk5vq/ooJrMeq
snAN+11RNau8rwBdek/5TI7ImOnG79vY9h8rr8IANeTrIWIT+DQX5vErVo43w281
JaWt58fGhDN2F7f9NAaIYyo7a0QNl8bq2YeQX7+IooPdHH5vw9zqf5dVpPStJnGc
xxQwi5VLMehuh/qmHzwP6MgsLj5OQQmLDWTLekVeg+vopLrfPZlCIPGsZNpAQYsx
VW45v7t0M7HhtnYta8DWo2hmXO8l1jP38Ydf+rJYkZ5+18cnVuAwihuhO4bqWBEY
OGZtEkirDHjPcGNHYbJfaF7OJvtboHcCvXMV5Ske8jGk1ALSPnDjEYpH4bZf7MgK
9Q3tFDQQAFiKcu2HweZLzVbPnhfUgHlZVjEv4y9Tg0byb+j5+ZjGHdaIZUAwPmCA
5Dm+trSx8F/7ic307Pqm5UstTYfJRbSzc+aPbHueUk1XM8a2c/8Lr14Vf/0iMFfm
E39NSxoUUUuQpYUQ45LB1Pr3EJFHdf+eTclxAIKaQq4V1H3i4E10If4djm5LN9fA
3rBQqLBjOE2pC36gaC88SIkHxlfiAcHyhFf0WlaMsDhgKNeSXUC9ham2t+oYdDgE
4+NN9J4JuyyIqtLUtoyMGnP2DHZXjtKkaNHKy0XoD8J1nSYoJNfSEMBla4DXA7x4
5793KnE9ETr4Ynomvkx/yNrSj3M8IKLhgmKcf9tqHywvPsqpttso6TBPrPzSf0Mm
2YyeQOIpMh8PmNZL7VVc5jI9R+vxQ7GVIixPzz+F7CHq7Y80GOVF0t2fxThqepN7
XM8z/K3Gr4YiFzDWANO8U8M9oryoYGscfSDzRTUWqHn3dM4yxslTvqMRjL+j5mXV
wFvtilwAxnhmCm15CLm+gAZkgnruw8BEqjGIOfaaLnr1AOXOCoCLgNVbeGC0VSQM
fNT9iqE+qh4oVTtrgBoc1mFLfi7ZpFREzUU/7qwAjU45vF/Z6Vc3i8XIdjt4CNol
7xfVZ82vKn9kY29UHkmrxnyk+4ifIAk8f5hSSTIPmDLgWklgM5xw9NA3YHerGONl
yMglCIhbpvVB2pzODG08wETquvNod13vWqBs9JD7tWmBZ/nq5HpNzCXO8zbmMmys
vrlZmHhS/cRzeyGiBirefPTydolhayuE79Ynh2oMlCwO9jwtdWexeBx3h8tE3F5O
dNkWtUMmmU4oA03mEoLsET2YCO1WAWlYbFMIYH9dZxOJkafx7b7jiOhJg67RdL/y
X75nVQM6I4oIJzkZ2VDJnJN3elnkxMAgpJjosQtOBD7BeXNcCpYxdTjsIT/Fx3Zb
B+W4I5LRJjbYi6AZFN0J5Czk4cRgX6QaGzuSAslTELWleRo7O9+WdL3FscjpUC6r
dExds0SU1QqRxUXb10q+BPolyuXtSfVUzrqiB8lpynqIBIcEoV/wZKW8VVrag8wQ
sZaZYrGelXQSeHQXFdJnPo7m6t+/0zZwbPaEUk35GHPJMtrW7biX0Kf2cuD4ojMU
LGhYxEjEAMcCDSPPDIH9T8xnyuZjmYMgEIeM/6cMzfwVxsK3cuBwMMVs0Lk2UCqx
uQEqjUTC+EPrp7JC2Wb3+piy2wWw4ZdRZ6aUnPU2gQhjxCtDVV1UAPb0Qv0y3gle
uIbzBoKcP3nASUVgjJMrzdQYgKFupu3iALXJhHtFerel00P9iqfe6J47g3xC89NS
Ja7XJAer6pwTVq8QnBe6jlkTLpcFZiZM9F+GON+GHqgvqmHEEjohXPYvJJX12Z+p
93GnHPDoUtBdhgCEGFnY+frD3A0dQ2nHB/JqiK9Kjms/36mrQNCPHTKhD67QZnfB
1JUQ4J1fO3q48/kUIrYWGHLiVs8p1iQT94AYd4Pu6wXryCL+gq6iXVfMDx/HAg+o
XqlslJLH2yiWjDBKXE829i9chK/x1fbVUw/coY1s7fMHOE/KYNvRiUNo3yX9OihP
NTWUV0xVtathinlJ5Hr1VezzfaivH0dU77/c4Ryk60fAa01UuLD4oGWpYunaTiF0
bygy1RO1UqPSU7cwcgvxvAhOH7HHbMHaw7GYcXQp/LF8RgLzve3E8sN5XmKmYNKs
vaTiAIHzNmfj+C5Wh0is84gJe1scgfFbt7ILNjYPAl4uFB2m/8n0FYsWX6hjle5G
ieyPtpqtGQxuSt008nEfxnAC8ky1AdYTB9fOHIkyDiPjJz0xglI60koEtiaLbb3S
sKn/ec9VdtRF+Ck66iVqaC1RaRVHGQ7L391rdVzD+BIdTi0m7CJ6f80dpleb/Vzb
TKQvDTOzze1g3H1cuCVG+YaV/af1J8EiK31mvfHtSEYGPLjlLTv9b+z5nJ7WJySS
NUrFe98Yalvo7JLSxbESZ/dEdzaurEdfKz9FlMrHh+yVoa8xg5f2st3cUd495Zzj
9md8ga5mhRtfKqgSuX0ZBsEQ7psfhBo00lUwFUlz7b8gUB4iy2dNiqOKffydITNN
yNMDtgZKkCu6K/8FZ47d5ev8HZbARwuFc1ZMJmDvCud8kUe1/E85pfZa2r5t2UoL
pTnQC7NksqBkAlHfyK25fGFvlkdP3F3UR3f5H5oF1EO5TVxgKhZOkivDFnnIsJBq
XtkaYA+A5mCJkuEpB13Cp7siFuaRxDd6GXUqAl0K5L+pVtuL4ZXDJIp7l+He1CL8
UbWuGvFZ5vLNkn9NcSNTSLjRxX4K1N5RnAvQOeXpvNcmojl8ri/2G0HWtQa0/cOD
AYfILzpzD3e9uIW7AXf6R/jl5nG+i1wBZw+5+fgLQkfqM+cow1Aw+/fjK7xbg/Pk
/p8AG6RPRf8ZIUxTbnAwkB+QUarRaTs/+jRr6H7tkiX5WyL7KFNexvUPN1VmWEo7
N/pl9eDP7M9HWZc+YM8b1ovTHzazCnTK9QGmXoQO0vsCbkq+mR+2BENVPbiCpiST
INkYbLox8sc6IJYa6thF2/8IzJVszpiE++59lJiaBjY8UtT9felblkl8R1GoUZ2C
CrWBlpg0a1mfm1WNnIp4ys7wjzTd5FJF5AH/2bRCg/mc9L1gz0EEM9HIcdyCYCRi
rApHQzh8G/zhRwd85+57qw7qyW81zJbk0EF78zqCdsgfiLMlTajgf2PC4BJuM+JC
YqAKd8lZDQ1x8aiygctaGwiH9d0YXoxj8hemh4e3Gxr9CVBNhorNhrSJTfHiDCTY
cMasc4EiLFkgX14Mbzp9Z3O3b7i2yrVBJIJqRoUdX+i6z7VMdvFr5rKxcvJjOGYp
cye5qELtRVNKTNYb56XG3+TLET9GAUxx3hd2RdTEMwnQulP6AXEn6jOMCasdUYC9
TL9yvKWVNlmn65pqMLfeK9hWfI1RmAwN4Ae0fqm4lJz2MGb/dbEfuuA3uQziWRMp
qXYEIuXLoiWjeRqwYxGK+oUThKKB5jywESqtSczUAqvwdmD6oBc11+lS7kVSNhXX
VvyKGiVLUIoqPB5qhRwQ55hvfd79QyS9IeCDdLO4HJUlqAj7kBNUteD7ph10tgVb
CIspSU4hfPvLA0TheAylRXXqE18G4i6rYhxZLxvbHvu2kB9yU2w/AJUYQ4tkdGDo
q7uqkp/WKScYeLP04z20lU/kkTwr/c7HUAyMXP4T3Zu+BgqwlCKdCGnuO/3auoah
pRSn947KBrwGcjg/ufYWYAenGZ2xap664Dto07KzRMfowYbUYGHvFTX5QeCpxoJL
nFnoOsDzSQc2AQ9N3El5rvIY3Eq6ZXQYGLLA2SUv2+8EMbqdX+AXLIy6knfexq/2
jMXn65aM6Mxxh2AmL6FyuaplPVqvZGk3TU9SkpeUJv2pj8IMZHtiyfrEZr007P6h
PLKeX4tuInHnG9F0l9/xvqg4FpkX495xTn/hYT6td7XRqUSXv1qce1gUv/qrJ9Uj
2epZpgIF6ahgZDrAhxGkOhrNMPa9YipPdvaRqCHb/3MzkTw9qTEUhofubqJolm8K
0NehqTg86nZHszKlR9viwdJxMtRwvY05QUgX3f7gDigRseB5i4NoaFjTOzT3m7oG
k2nZYh6yT197QYuqUOPbz65Y4xkYvRwKq326JZ0PQBE1LSL9GvfYGzkGOp3Yc00l
lkaLsAU5Bie1QBbupjG/4J1OZwa3FUDUwqaiJJN5mZbtckQ1jX90FENMK4jSBDY5
WdjXig06pRUusiuZsZihT4uzcde1Spp3SStPl2CZhq0v02EoNp6q0P7EfZD5VWyN
wwE6zyJwmzbOI5mMleCu96EZ+8QmHF2bSf7yTL31t7twtnk1s74elbQqGWwSDsna
3Kg7qTzr2nyTWV8P9/JZiNeq9okTmvwJgGGR3sBNAkS0Frcqt1YMKPs3qtknsQ5B
GhEg8DembyRC6wE/nVOECz6NcW+bPUlFy4nvTBt4IENCPeVBHpFVBRcurHglmybH
yz+6ocm9dsrYYn8ulJrXdVUTtIlJRqurPVu/02aTD7CZnZ8CDOsa7cFmxjsh30VD
45sFtM8UJaCCvQ2lYpafl5hem1yHWcYHsVuLY+VVFNESYp9OpsxWtsbVfBZrmg2P
JZIFUkR0vTdpG+XB5UgQ0T77xG21HA/O2fDHwtJECSHE9T2Ihg0YNSUsGTkcP4sG
ZUZOqwJKh7X4jjOmRvYDFNym8YZE4kkXeeW4J+XA1bDhAS3KZwKvS4m7yKxcwFc2
P94ZhZKhTpwfK3SLgT9gCL8/HtpDsV839FWMLvECN9Lh91OsQdMLKBzV1MvWXaCu
PwoEATOIoHQoLfzBRirkiT0FyIFT2pK1kzkRtW4dxWhNmRegPSB93/F1XR/h2g8T
2LRJ/lBe3zTPEYzc9DYf14N3IbtUxMnkJsEzNA32q3RHy1wpaQBuPQx8gULjrMrE
YS8lU5cX1RpZsGFeyozjQ1/XI1Of80fxEBaMhP5zDGJqtQR7rq/ADoQR8H1iQ6pj
xHSWOJMaruoqo7pPL0RdNBYvaYE6/SCm1F8YjAM0fBUKFoBIiGygkxiTYLzhk1VK
3Kk7AYssr8nToKIjSNHainYPoVzUaiuYnym2rSWJiu8GG0yfIUcBIJeOrzET/CnZ
ifr7gcW0SOyx/5ohGjMpCCMJ7O8zcKQkWUhcvEAmobA+Cr4QpLYsjBLoZkdTGgK8
R1d8FNfWGb5UEBEw++FqyGKh4CiwqMYGxw5MrdMURn6zl2Ayb3pSX2NB0shLmyrP
8FcHhG6EG9VanIsjYD5jehI0Fi/v6CuoFLSrDtI3PSlcloe0q9R9jp3VV9nA+CVC
2h2r6G3QWWaikGCyNnRHo1U7yAHzehVvqeiXHTWRWvw8zX5TaJORZooLFbw+N3Hi
aTAZKER5b6OmSHUdXG+TqYxrcWcMPSqIHuBuIsJ818gLcLAVzctondMSNhFR0yLq
gUlVMZUUK1343Y8G1FOE04fAlJ5KaAsEBSCoX27mtiZxtVJnpINhRfJbevntij0K
78TPa+O+QcbLD+yLjxBckp1clWSXqk273/1RuFbY25ItN/uAqsqsj+CTY4NPQZdT
ANtySszRTXAQqv4imdyKf1wZhAElhkG4zGhSXkb6J0T7tZU34L2LkZYGO7V3t0d5
Vob0eSz4+ULSNgyQoGkF/FB56/CbrAkCbQQTihKfpYlQliI0cooGpfGlLv9sEWhB
mmcX4gh6dcd5WvY38f6iFXb26YuRLY0jIhABYNdJK+1gIj/NweaJQUENUeGMKdcN
3ar1SWBg4ZWm98S6wDDVIV6qVfkrsA7EuFXXgpcHOFxBgVWjLUim3VOmB1ZK14jC
zoE9kqk8DFYNpqagYjmc0NUyl/+jiK6DSvbJ+ElJFc+EqzG1WwM3YO0U9YJ9tDcp
LtpTsLhKhVdQSB7NI9v2g5wHByOr7vdS0N+lGK+OScMMIE+2avvrc8472lvkCMPZ
IVu2ViEBurmZB3PAKDNJKdec5bOfpYsfRoVv/V91vUeSSw8adUjmz9P4Hf9N7LYE
lcRw0wLzS3joG/2Gi6JqRT9myFZh9464t/Rbfy0WoIIMts3k7VP1EFxeDHxcUFAy
X1a6R7SefgAM8YoxRQepvlmPJEvBrpVus3KRTaZ6bddAr7XbDNLYEMzReXLMAEiM
chUoBrY+aap7vjltg8i8mgqcK76EfwWwoR2fRbFQV95TrzRCjlU1LO4kwdRqTGMk
oXSGmMxFXpIHCyhtD8m+cwDvfLYxQYJNE1yVHFTxCLCIWGY0bARvxhGpBZABP4Kk
GCDS6C9v790dk28v8M0W0Z9jZ6KSaOAGbVZaCW0VmdLAusIjhW1nXP383SE2k/Fg
Exg8jqpuCO5MweajoMIRtg5z9HMbNLSs+nqAio4LJ95dBTth8sBSx8NULbTtOvLf
mqGZ5apYvSIMrIG2bMyYql/etzlSZ3T74S5Iw9bNVayINstFRK3UIjdwwMe84kaX
D9PVb0kLSC559VfYLe8+xn6fj+7pAByQm9cBO7WbrtHmpiDmhGuzUmzwg2qv2OuO
mui10YmgtbH68SZ+KzhRMWJmoa7vAY9ukJ3mGpWBOPTGqWZ5AvGJU3diJU7Z2nYP
9tJEvhQYnfkCfqpj8qU6Bg1f1d8W+af/9FYxmsvgNpJsiP9whDc1ukb2ome4bi/v
C2wkVQGnwldBaeZ693r7fcxAtRFNOn9NOjW5MspNhLy/kuF7PuofjsR24x5VW2NA
bHq8xJykoPgusm8igC5k3bw509/TmqPfxxhZQZgSr1bDQlWesY3Aru/aqByonew/
VQdz6RzIDXsfeqpuXS/TDP4S6DuDOUuJn/c9nZ6CUpaDYj7YoRjjyExJGwG+QZqi
s2xueR/Ts5oLVFaD5bF8jIVLH255YpGNWLTjL/qfdmGnPVgonhpZfAae+C2UgmpW
JMxPsktLXyl3KZW8N2joI7KeJuDTZsFAN8VShk58H7tphh10NrFqbMpT25JaGZpD
idmUR/5SuH+H78OrPT3urTgKRSFJ+Fku7LHv4gfiCSCT1ccT2nFS4xZeAZYOMdJd
mJPvCaNLA1DyHCOWhgghWFJcCed3EcFBRz9BtEI+S2dIuqJBJI75J+kFHcm5/Kib
ixaNDCXUOGF6QvLovcTUkTwIlFhEh3pwtl8BjO4TQx7vBIZDMN4TPRjBKwkylDAp
SGtnChWlIjYAR1P+xKoHzwzNxhHkVbw2Ws33tulqrMZbUaXINitvgShu7w4cMQCq
SQA5HEO8PYFkeJNLVVVo7Hndb+0KxH9s/0IR1srVuFW7GNYjIIYgjkwZouw59RvD
1hhZBi0JZCb3bFJkwhhMCnPtrpkG/tYAvaw6WXYM9D1cvQSh6+oFTwSpyUuoG8Ie
uVkeC8v9qZ5WT04wOxOw8iHjsxXPvyvppCFIM8yag5hmltEFZeGdniBtRrfNYMQz
LfzD0MTrKt8Fx8dF739G/I64ekHI5rRTZxCbedMmnCKh6VeiGID+H6P1OKMc9Y3L
46PVqlqzDR8C6D2KWmJZ64vlFEAGAc3PuYQN9Cq6pMeBZrFgcKvv+nrvAkypPrgZ
AIOb+MZYawDJXYsY5dJ58crdZ99NPeMY+tk5Fjnz2OOpyojGU6lHhWzUHiur4jhX
Pdj+a5jhg4B0CU0u/ysivBYokQEbByLNXDAeyQZBWJ5w8S7rm5Qgq/HP0PRoKr8B
mMApgNjU07i7B4crBgcpEfr4kbI2T3rLv4uYTU2ET4FSpf+1ydd8DGcKEb/uiH1t
OPqu3U/5tTJ4TLgDuWcb34jRzwqvEHNl25RXDQ63ALATSzcuYgx+rgwRwum67ACP
5MZSBeK5XiTgjvz+U1jFsfyk5t5y9qFpfmFTmvkTHYwrofnSwme/yFveHk2RqIJh
yRljBFF5/Y0acOO3+V80WwMC3oHDA9S/EloQndpgimt9s5q6wo+90M1iW/HdFuXf
vJdp8yTfHKpFIjCz0r/bQe5pkKubuHzy+6p6b2y6ix9iO7qj9T02lhT1k7H1wIlC
LtTRrMqRtTRlyCqUF617yUXwKZvQ3sXrFVlP8xeFvFwVKTAkzOdySYJfk+2vFFZp
vAeznLgHvcV4IC0KwcjJRGTIFhV0aOo+fNERGz/r1jJgbECSK8fFRzMEQe23BaRJ
c6IN7MBXUQOKARRUeXRMWsqswSB6tcrkdjodU8z0ceQ5D2FdNZNBm9aRhZiQ9dFB
MJAFVhwLTvTwzT0lWz/3ip4SYQ6EqjTTGhPImf2ozVl9SCz983R+lUA4iZlabcbB
r1YXsUFLneNsy4by8wekt2KB8ZBzOcYMGk2BTZxg2VEeMQqsc1vRuUqfnRv8kibN
t2D/NfcvRbgLi1XaP/N7mBmMIoViR/qJbsAYYIUAAxECl/D21qjve9HLGkhLBF/R
eb59/AkZfN5cmzlDpwtyLHZQ7Pl8yEUQFR2BXRXmrsKohDk2f/FWXN4CEloCEwOt
cGe71WVAGFUrqt3iHUkbocBX7SHbIqxhEtYerluTjR9dWr2WtFVW6tWw6kuA9zci
4slFQRIX6bq2Bw9XT3zOk0w1J9qi5xg1Aode3SrKY1menEcEGldW6S6aK+wfraXt
/3VPk+2yMvS56HL2Gn/vYehPGl1ETOH05s9hjEIY8Lprt8KKa4HPMJGOF0fOXfJQ
GRREq6EcNskNvCu4lsppFrUMdugnkA66KNZtyZDZcb5RZlRNaWNEAplFpWe4kdA8
DbbEioke4jb8oczAmEfbdV+1Riv8Y3CFwR/bz7KhrHQ7fIcY20LycV+/gvb202vb
W9MCqkbvJwdHwxJ96IosItpAY8tZ4bfPtM1rUh82aWWLpWzVpdmwscU8z/6t2tdd
P69n3+uzODp5SZEa2G+5oymLlPEC+fKsGleQQFfS8LhQ7QAXKaB4EyYlMs7Q+hIE
IFM339tgkM5/7hl3cv4wlkkZgDhBSvEPYyMGFxcXfPP+CEZJS9TdVjt83JrwrHZ6
ZVFwvlqjDuVyCGUibRWgbnCOjzjK4itvgPFM1+8qqBwVZdWyT5F19Hhzj3BQL5iJ
Fsa56hWJOpTyJgSlnlDTdW6RqizhuOIoxGjlAEvLOPDTKUYQlAeszVNn28l9T+mF
bd0BK1sbAFxcYTlD3tZaL638A29m0SHBSt5ezZj1XDGGv4BAeFeLEQl1gdbYL3gg
TKTHNJan9wsiffjUurouNMqAVIam3iYIGd5LF/xMYsfEm0EqNDo4BQKbsZSqExWS
pqmT1ekaL0kvOFeu9yL/A1Y83iIBIn8Twu9GvGraVTDy7+ooywzfOSNXV0w40wyo
zAn6RGjWVuryNlwB8x2kGPN/7FJN+gQHkey0eYTDu5ndes1RVG3mNlC5KJAAYopi
JjMxXyKnMBSVqoV2O7kvbkEqqr8B0a0ThbnARu/D76/vZcp7YljcL+bIINKFF2G0
V0HOogqPikHCK31uvdIbB7Pa8SZa3JX5+2tTcHlHHpaG/Q3pbUR7RvBWlwLjfsav
j+L3A3vM19lrYujtwQb1h/syfBvoWZYPVa3pPACEL/W1/+ASJ8vOH+IpduDFDmNT
C70/QJe3GzI+izZpTSl3gcPcEoPPogUapnyOBtM98NOi8731cjVhd11hnnbxhWSV
asg+PRfZ53hGgtS4ei2moteEgYgHHyzdSv4GibNLTE4dVy+omB4UegmjdMqdo+Yf
Dc6NEjoc4USw877gGII0gGjB4C2EJYHqUXSiOzXNt72ioJm6F31w3BoNDyRfLxEw
7cHmCarEBfAm/jzo7ctVUUFZXIXNiT7hr7NqEFwF/OXTW0RSoQWDBXhWtQUa96u5
lPp1LflctCn1WmABsUryddHqscsOGcWO3c5miCd2Btu4qbhuB3nWahzBAtvctGcE
r1O3WaXIOGgJ8+vPgck4UjH8k49cTrHbFpQPlJDZs8t1MRIsrLPLho/TFHPa9pb/
0msDjRy2ki8ZiL00mt+MtbtJZzXys981/yggVazo7I5zGN7+tnDbb1uxo9du8Ndk
LB+1jZLcC3tYbH/Sap3MKd+5gFKWKQLnF5gpoFtyqywYZZFhl1GqIL3Jz/v7QHZX
XuSPZDNMjP0zSDXYuyHkO/CADeo7uVlsDbZZ9iJjfjKbkk7xUFmTihpmpG8eyLHQ
15FXz84Ak50At6a8vjMIoj6yqUqruFABVUTModR1wMbc+oTd+HUi7s6bqo4sr60c
b8hGehoyTcpRn/fpDgTLuHKrh8arDDvdVI+kIbYZTHLJZ9PCRPlyStF9F4VI8SFb
P0dqEm6NAkVnedU1kv8e2VbgZn2a0K+qtWBXTnNKs0rkmth20pwLPucrEqc9qge+
4Z9Nenfmxt6F9KlyK20m/iVIknVNop/SVA5MC75Rd+KFbzOBqvcGDP3w/c8rJGzG
ZHrZThSGRmVzFwPJLbiQnD7KVmyZybx++tzqWOOpBOaLqdhOFnpb6ZZeHLyTcNkv
iVIB1VPlsy7wf1dBcDRKJYrNqwcuSi6SiIXiRBwLymEHMUD9K/7R3R6hUShlDnuk
v/QCgIpPr2Oz4oNq3DXZZItUTDJWHpNlA7sm6vQFFGWJySN+WMecheP7/Pqh2/O6
QN/ZU4prYV8nF3qV7ZJ40vAUQB+bmBRhamMkvh5+7XbQnRpBH+BF3Ena6Z/5eRt7
zzPN4wfSaPPNJzK9cJz3JuZjBh/BUlvDiUmMgEpcElKhsJjqraWHIFaoMf/PQ5tX
GjHbuV8990ezl2pXRr49Dd2J8ZmMsJXyJBumxau9jrITK22LuTIcDWPp2MohSVg0
aqONIx7snBq3EoGLrH0ZozoDSomMW+gbGzYTwOQifRRXPWjJ8nkQh1ufyOj9Np+C
1uIv3rovYhQffe6UYS2CECpdlifdysexg36aMVsfcY6K9N5q32wMd1lB2xnkig6T
E9iBGfN4sNO4m4mHrWYe27+duP8aQjA41zycVqhC//uIT03ikFTv9F2QZYM9OKoc
DYKR+hwBKRjUvrCnfkm/cHYAS1SUAYOzXeb0qR5/kNg9gZ+Of4Ww91unM+soCMvz
JqZLlOyx2BrpXUjtfQBWQA2ZvdbIAfZaHNi5HNMLchjYSOzbdcSrJWB0E4PRusvk
afyPDOVPTBB9u7FiubkTnjqoZSH55Pzs2ET8mwbzQ/85JD/5K4JfxYhNh6vkEXgn
4BL7ImHFwaLIGDS5QKbOMieTI58UXLBrSVWlSLcmY7NREmdBDcg/iEm3o67JqQnA
gvD3rsjP15Qcgc3GBqBihX+qSOJp8DOLzMDA7Bf4OU98wc2HDUHNZOuQbcO0X6ZB
7BKOGF6pxLJ7IoMXiCS0Gr9jl2sl2s65Eh4xZ81tNEkmhNk5LvhVw5SRZ2g7u1KK
xVYbHgx5rtn7fMP7Zab+oVErNqMqQPC2+xByFR+goLBiD/PInCH4h1kpDpHYKLWt
p9iQ1l2vECvCuBtDqYxN8uCL4buLc2bK+OGbfnOW1rRmW2ZbRhybMI4h/unHLMM0
FQS9ntMvNWcAGKzZF7zMBVprg9nNH5gZPy865dHN9FIkUZlemFUx6oFRBwL6Mj5L
u3rlZHRt5SDY91VvB8G7cFNHFMOt1kIJt7a/3q9Oka9eZozySwReGgVlfXJLBjA4
uzHoOus/MiE88R72CbI2yHVDOoh+HzTAEqGKrSQfTu1+QAmMmTQnLms4HERVuLJg
iZw5FBHrsUwA5ghNpPs8yvQ6f5xHVWGGu8o6uRk/kuqSclvu58LAboFBSEsbwDnl
MDQVmDFXHjIvyY4jHNGso5yH9y1mq2prXa2q788xD++n6RFjJOiM4kCUZQdC6Gmv
AZpxZeWZK5SiPZR9Rc6jD0k8v05MEjjnqgYoELAv4ujUy6+win0zXq+ttrbfYl9B
lZVDg4DEkT/Knuc+q4zeKrEzl9tczSJsTI0X0UVTCHFnAfW+7uoCyvnRZzilelyO
amQCSdWzZNt6mOdRireTBhZ42o1EiUJwBMKMrmiDyzYoO3Lmy32P5zfU3O266gHb
anrtN1AmFtsl6ZKDcGZfWKQwtMvrnM5nAKyk8qd6a9lQRjEpgDcJS0n9tBmsTp56
aD69ARhRRxyZ8RVHO7GkfzMPY6CPHntibfG8if/V7FexaU2QbWhvZdcReSr98I88
I0zxlsqb5FnSzzecYDVx1v7CxEcH9TjvLFTCV9zIFz0DSa8u/+l3OFtYa2arRAY3
zvkxr4xJr7V3QFVBZsQNJj21Kr68VYJqUJL/vGkNruWlPSTHMIaY9fX6Jew5CzFX
IcSy1eZONZFvAWPKDtTwE0DBJaeb3Oc8SfF6+kQrd0/VAC7F6OVPWO4CbPGxlAXA
Fd3c6tCLkRlUDgq/FIIDepvzHQWYxXyBQmhL6jB1pHGTGABtt3hVVI0zmJ3SUQYy
NY2g0ZVZgNyiA2Yg1w2rHvgsfyH7PB4iFdLUEiMjtKW9+Qfj9GoDYkd2blPA0MnH
5oorGozu4RwRE+A4sqIMY5RdwjncWM45q9UAtCOnu+O/3BViP0dWpiSTtHHOM9Sc
b7W43o5L/VPh5xrOrMEK0ozTZ3okfd3IYE2VUwI/6kU/VZK5ItJiK3wAfTrpkOa+
5rrvBENl4SoHhcheRQAjznXCdRvEqnO0WA9VdlpngnQLwDR3dI0jFe2/+aZmQil2
ujOvT0Guv2kwrQIj0vbpGxWuCyY9jol5tL9qXVkYeo+hlACIBLysg6ahwYbS6Xv4
oEkvPk0l+Q8sXA5TKVC2Hs2nPajcdud7/TspVHb0doZvOzrcbDWYz2atErZXLak6
TDQICsFNZlF5kAwysfDZijuiryW7atN4YHyolBkcxq/wbFWEd6ceyiGHRu1VzR5q
aJKWIEFgPc5HD5yqhGMqY7qpGRh1KG/TmV32/3r+d1g3gJxHvcLzpOyJ4dxvA9d9
JFTVIlnSE97rukIhYtTFazOmotJONxxqJjJdd5Ysybu4IArjcZA0TOPPWKFdqRaR
MKpuzHsQ8rlzJfOV1hUWORIM/EW6StBfMGKFjvfWaoITl89gJV1b3osD2jc067l1
V1JPqSp1Ho3chZMg65dDZhj6A05upd8VOrni7tqPO6vac62biE6CbZCiICgAyNbC
AMWu128gDi13KOSQMRikjNzvxeGy5PiqW/DJktP4t2piRE6BDDT3eq3DVMM9oWBO
FgmaC/BzVBJ6KYIp7x8WZ0gqxIbnkjJtW2yARyv17r2vyariwu8h6fMqwWgHY4Jo
1l37RZtiuyYWDrWQY8EA5P00krShCxOK/vPM0v5vAHJp1k9M+SJBm8UcdBV7YU9t
slgCs9QSzpRkk9qUk5UQ9tVYv6ra56hJxj4RTtx29gPpergq7+HehaPOZ46mThe2
Y8S5zGAC9hb8WUYhHiYA3IcAxvumbPhfdgbWkyajHhJ8AIvD42m71Px45tD2UISu
AoBkz5KWCqadPy/8i8eGoFPPFfR+AIkOSbKEcx5R0wwa088IggaqHCIKSTErrBQ4
kwPz4xQ8cTF/L3fZMUc52+mk7ov2nwTPpkX5z6OfI05gvUdzT3yS+5WP57gtF32Z
N+0H9uJvIymCpPJ+MUJx6P0ZIXa4d3Fxoced2XB/HKAT82tH8i6teEPOfvrPE5/3
pKmk6qpCu5BBviPjdzrv6tHbGG933VhaOk61NR6IHeUXyO+sKiA4gyPzA9EE6VOq
evxUYz9Lexjn5ZWQdXDHpmtT+NlcJgbsgZqDmGeU93ZdeYTP2dIJg3QPZ2Se/Wt3
28TLkspcDwp24dFKHPavwz54YMX1xbyf18cXzt0OnyyEQXc9NKhAA++/snZNzv/3
w/glyI0rrOjX4PHnfV+rK9xUEI2mKzWGB7INZsX+1e7IzDciiX107gT/aImrnYJw
sshKaWf8VnJfmu6rLkn2FA0QX2eK/B/LA9O0CvZvJnt1l8bn0H00NyMNPt4hpBXV
ZSCN1MPa4F3xS4bIQ9KeKnIn06lpsEcFFkXVlC+d90XXrdCSOUCoIGNH+yGduQgO
kfxSzmqp2lk6TVHvT87gi3JtqqMo4dUNQK/i4AIuoRn/eUx+szTFf+TQ+ahtOngO
oouKeHMDZtFKL3+XR7vUPKcC3VO69Gz3vXPKWMUJMwk+X8C0z+Siv2zePn14AStW
Envhs79Wj6MEBZTT0haqQwaFYo19FpbrmjTw8rnN0wfX7LHQj9ojpCY7whEoco/2
3EHv1qJBWKx0cLmGOd31SDG9raKHuDHxeRBsrDIc7HdAAOJ14EZJgCSzsYjqdguN
t+Bj9KlEHdDFWCHCdplxJfqtJWwWv9FHF8MOS3EsAvGHotuqCuwhAAKcKDdEgqDo
U0f1imEezaV806Cjw9eYWaW8wiCulIiV+WFQ7n+l+Zq/aPz/FmyO6pNqFUkgtnzi
Fzj5n+ognqLKis3MUwRr8LnnYahJUvuomxaBH/JBsDrZFzyHOvRZ3DESVs/bcp9r
5Sb7Gfrmjp25OgSLltPOwdpKBtabT+Ntz/vl+d0TgYdT+CVyYTKGjUcVX8BnXThA
1xQD12nIlB9XOTrwmWuSyV7lgDClKypczGRT5+2S267iin14NfptVHSX1IODKQ/j
es/2i7iiSHybZesDgimgh6PyNp68AuGy/mspM6Bn5tHl3lfaxd0MvX+KVUSxV1tN
Esxlq8uK3Zmg27UoNXTpydgwCNGnLCxX0on10fJYoVJXzlNZziGma7+biuTGuhJi
AqtfTwTiPp1HqyNxupbCXm+msvfWF/r7I2y8mQawHIpah/P8kmX/TumBWThWuOVj
GjEr6ojJsbJdQdSoVxrrxFsAGkc1ddXOm5+r1AGAJKzJe7ojKlaP8sKo/0P96BOn
eRiG+p2SSAHIBgkJRjdiMDXnpXe3mAQcabr6zdcgajuh3wnXFPaY9Jt9w+ZUkp0U
M1wC4AXNKc3WDhHOz0KYvjfDGQS7pZ7VCvVb0GnuHnhHvTSr+vmfUlBoy3W2MZBF
x3ihIKrTzFrUhFtvUQuAHrQ8V9Tml8cocDWMx1qvsZRNnQymDkOk/8RKSDRSPq6v
7tG43kibUaaYZUynZ33xoXz/5wUhWckvrgkVNhcklaXOsUa8DzeLohkJfleTVAj3
96MXwEZ9S4F1kLMnZLZJDip22Kg0xdhyuUYOnQWnyiX7vNFN59ni47smSwLmGXVv
U5Ey3y131IhauU/XOLrGi/qYR5aFeCVk/4EBp519uof+lTNrcC9K8i36LN0arg7f
uioGQmHPdR6mSOKFjsmAS1cdUjj/GCvbxD1Gsn81vt4zCAyIbyEsO2dfT0cXnbk6
NFBhivvTQg+8Mkw6iIf9PocCxF78x7OArRvIZcVPTr1+BPiPUwVxOMaSJvjtwdsa
PnLT8w09xkKY7nWZZ+lusNFtZX/0kp6P4C+nfCE44RKtDYJqKYL5JMfeDc84PSIt
HvAmCSDeLlUgaoO7Gq4YVnDCyPOM60aYRrzkdziAVEOcQkyFJDn9nJUTMhCQ7mmv
djZsv0b9viIixHjJHgrbwTdbMDPYOjlx7CaGzDJMUAi4K/zCMppzGI8nq2zdhOTn
pVOwVwesam0Kw3keBe0iWU2Bj9ZqHwlHxgHuDwB+inHK1PweR+jSuVOvPngf9YTt
K7l+X+bZOSQtSzaHMcu3LB9/B2152Q8iy+SRWFntDI8t0D0wRe9aNcb0duVfMf0c
on3sHF3sWRuXIbgtEDxhStCPWbzDjZ0lFW2JWHKHQhYUARt1LS7SeisT1O/Lx3k3
7SdsFR6qHFAhhgpZGyxvDBgdD5vu/oRn+gXaG9YhrTJlyTNSGop90gNacBMjLcVc
zT1sbCQl1sxJM8PSR9eE2h8UUW+fyVKecYjncBkbj0niOTAVGyWgs6QL98EaCbRP
OBt0TipcAeeNWNHSsq3foAV56JuINZnssDcyV/zBDOmBoZKquw+v910e0yIWUxGz
Zoj8MqSn7xSRhg9v9unwc6WjokKBXkV4r4E977Qp7Wy5rAC6gV8+XCrT6WzfvumX
CpM5K8OlLxyR/rQBoLCYKqKhJRGrFz8D0STX6EdfHvOJvD4y/X0bYLgPy34VB5q/
CMmKRy55PhiIyFR0vr+AmvH2WVzSkpxqTPKxOKqYALcAey2C5nwx9c2B/zSuyo0j
3xPTEbZcE9Kn+XBKQHu0QH5RhS7Z8X9toTerjDIztsC0sMEfpH0EOskAKAVmvjTj
EWnK5EMNA32MFn8q6p3b3UYCdchktI/why91Azu2Zc25lxe/QokbHOorXxQofBPr
GJM8J6XRVFuFW6ZLSKF+lA995qMR35s/b7OOW7aCTYZoJSoHm/wuX3d2FdtCfe8T
8/S8nT3Y8pslyvMkdnZQhBhcnlVpOMtSMeBCM9ZgwrEhf7N3EmpSpI4M/plGSyES
SzmXap8jzQKRWXJuEyRlVkMXiN4DuF3WsMTZ2ABFAMrjg/FREJiWNYct9MGwzNE1
P4RYgnklXftZOErN+H3oM3Z4m7T4SPAHi/cm1B55DFyS6jhLj6a/S5VwwH5TTtUX
RFtFEpTvgCkrnDHb0LdCutdbMLeunUh1zanZ5+ZXPkRydUECdLp3ICEJDsxotESP
k4Y4f77/y8tmg0qGX23Uz0tYjti3Azwk++WogC+XhkH9B43wuPJo77LEMKJi10GO
5agHMKbNS6O0lEiNjpYkdumDhOD8N3pI5peK//B3eiT0geP6nrD3mu/aVmxKfkSw
YLWzZteSsKy/A5ryUGtHkPAqmnRthRxVrSww03m5BfCKIxjYYr/785niOLr/L66s
8jXfV80XhibP3Q+bQM3yNAw4FNGoZXT9J4phsrkP5zT3jU7DG6psqcFopT66h00W
cJzokcV7iJSwIItcn2oHci9mBSHqxzw+0yopDfUxchzgL5X0boLnLC1k6sdvNgLJ
DzNTas3MOxy1Y+Nqm+TWA73i7wGdz3rN8qWL/6xwfCPSA93Nw2mvcCLO8E//YYi8
c1MKNzeRIdCZewmZu+/wX/7lYqJDspAEkbK71D2lr3RcgyyY+WbfJoMCEK5thuc3
u6CV+m6xHPA0gcxDAd2crDXjp27LmWdZ7k4EAPXEx/yurm7yfhyrpiEsW59HL2ua
FVNaROChIMSSX3At22mmw1QKyOYoQ4nSmpp+Kpels0himfYWFxpUNxWolu+et1j+
NC6b+2/UkLg8XQ9uhRsQuArT/cPcVr8OlVOa6O3a4g0c+8YUl19fx9/O28HKdN+o
FYA5w6QdhCZvVaLPCm4vld+IbtQ66D/3RQkirorpe0mW31BEYUCmV+ulzrM/4KlA
qPU6+TZBX3gGmflbC2GbLh3VCIJqNoTmGS+RtKyKyOaSPvD7WXbLbLl92x/6XnN/
By+jGHsEMM5lph3VqPaUEKUsN4OniSsvTN9igoj1HeVKBiEInU5N/qf7Bc84pvn1
f1jEvcYJMWIpArSFaS7BPEfssMyY/AAIkahAMHycjBj5izy8epw3RZ7NnlLwPLq9
nFnrkhXVQp1A14NQMkcUd8mC+OA8WK0m6txs3Ft/69MQIVuoJ+ou/0PgPU7oxoK7
1+7k8jwpXKtS8akyTKDtb47yMSU+lHafXqlqpoq+a1vFtMDkr/McEYQFUthd+zlH
6lnsbq+CYn1RHS7x8JClDyQi93FLO0eVGr4t/aRQEfOkEouKlnDK5BcvdwGI3VdM
x4Z3srhsAu4pU8cNPdhd++Wgq3cp5Q1HqIiFFRYnBwVDlHGjOjsOXRrs1jK5pkEF
5L8lsgOZDTiupo+P8tSacMT4a2VLIx5RcMIpwJs3biJ1C1MDoH+mQ6lGyDQ0K33u
e42IO1QToMaiNlRa0/ZGnY+0s8dRU6mSW8k5zp4Jt67E8+K08stAneW9D+6s+Kkg
eUL42vL5v93ywRTR22WKHLDZl5ECJO1lF2gxYt0SrBbcFnyTrkQ7lSxPMjItulw/
CrSHVL4eyKwdmouhr7nY4vwOMiJVoc5NLE4vG2k1eTFB00wnbQ22tNrkSPpaJZ90
+JDgGUBDZOQqfFcBKfZqRAAJOeXxSfvKvJXGBKaic1sjX8uzOyxYkk+oGBrzQIiG
esK8opdimHDe5DgvDqTjNKO3xEgIVisL2+HL8o+v9WKLWNHP0D/mB+RJzRTbQWNv
SmIza2vwB6qa6nbl/7zYw4KHhKZukDo360X9YaI/343iWOfRZ4yS7YIA7XtcTFo6
3XeACuk61Z4vqt0yQGG7x49K7ye8gzcQXuV2qR1N+u4E817tEyKEpU1cxotkawJR
tQdDFhMmciDnp7BNq2LS9QyEo+MkAIsL1ZGpMavDeHQyI4e16Cn2m1WymNttPebF
C7cUwB53NiJAe5ghGc5X7KKGW2Z1BR8YPm4qeebU38ZqQCpxzlvVUcskRsDtt/lM
OPgTa3Mknham+rcPn0GBtSclUF0F7dQcFeCydBdIjN0vHCsTy0s+jSe4ENl8sbbp
hUDBlej5eg9ExwQhYFjszPIwFY5SUlKQHIlqOHurKzZ3QcIABiCqqM3fSDTSuzro
CSYtJU+hE7XYhE++G+Xv2erw+DNF0i8XsqAyLPndmNVPGb/1xrrNFEqvMr8sAeB3
VJi2+UPTJgDg54TqyY8DbSc/dVi85XOV1MiDzsuA2ecAKPUmofF8Aik2yHY2JoFB
XySqAdFCy1TEDBvcRcVwCL9E4ItR8Xlyv3UT//7hCseQYnEGlyCiiA+eyZtu/CdE
8H+YPUppmvrQUpP4wciKLXvjJ6rSk1Bax3qFWw0GuWmRjDqAJ8Cw/yjlzxAHY2+e
4eJywzinkEG/HHzNU4UX/hAmtdcz/ysqabpUsqHuOqTjeXNB1vCFrV5OMKUjwcVy
ARgSEXrXKBvekXzp6jdj1rp1Kp8itE0D2gkbsxYr8/MGQU/ANk8kPUhv3VvqY/wD
7cGWs83ubdZByiJ1JvfxgxAzJxmW5ZIC5xsnKaaV/ymMxsFM+h9NB0hWF4fkiZOS
lYfrDxJ/e89Hclb8zx1K20Y8L3MA4fF5DnFJASCjuILqlO60I7A5JfOpayDsl9a0
ODZq0GWJamyod85kTBq1yrzZkhntsSvbUhpafBaldY2C4WrVyufB0C11lb8NbFqM
J2evFkDY56PKxcYdJUVAm7IouuGwosDX4YcuJ5kFTwfH26zcl7nzlbTBVb0zHZJv
Iq3aO2/j27mKqLR5j+XvBYfVNubkAc0XHJwTuO2wm9/ElFbiVQ6MNImmys21tqau
G7udA6hFNVm8AlEbRHYhM/ErVdZ4zFTWqEyQG8Iq7NjcMjoduGQooxQyWRzt6yw4
ZFU3zmuZ5UjnbmaAWH6pcoN+LPadUIOQ1noVvHRiX5CWD30RkWllYHcstdPugEZ9
9YFFb1c8RaHpFmgAjo0TjsHsPcAEZI8GzPbnBveVKioLGUOdHE4wjLQ3VpfVhYLH
p3iFqLtrLMxvu1gRz/nCnBS3OZVEHHqCUcXZALuMcQRKBmsHQPmOoel2FFTejBeT
PGqWaoyjEY732B6Q+7s416KMDGMdOiWseaYRVgwewzWvwIboBiFfZJM6bBMAjAWE
6kuevMb9EZh3DG7yTSdKrYqIHdpjVTeIB/DD6sR1gW8I+bPHkWzC+0LrDaLfddfq
EULmF3RUPOO0kV/RLTiA0vKo8kSSuPNXmS4ysYdt2t4Nu/T+N06KuBvMI0JC7Lzt
HleCrG4q//oRQSKaFbSeAfv0aE5JfISy3D2EEnW4VviJzCKMVJ24YeWxh3Y7Mk+6
KhoVZVb//0A2qH/czxoMgKlSZQfjgPvvoREeICJsJi2wy+aSjKCyNAR8xeYz+vWr
0PGy7eTo01xoX0GONt8tyjrkXMpLRFtzCa8nDlXh5tLhpZQnLIav49PeoGV/UcTd
hZa60P4wliKAfx9FLVypKPED6snjHwat4DQtIioP9kyr0qIshWnnggenLZGniQUe
saA/M6ICsDOEXaxPR6Y4LJgWsNgkxsuWCOpGapztLX9LJKgwft/jryUfwI/ol2jM
5v+lxKOm7wL9S7h/jGxw6PajBl61yLNbjtyCTYQ6OTA582dtTgPCZlPr4tbnZY7a
qT3Xvl1rBM3ejxJgkQ0V+2PlU89OxGa4tdaNmEcU0S+X0EWkFr+XnysReJkYQzkK
rn6kVr8mMaN1HDJzP+3BXfa4SPbVrdJOsPaxyrdUw1BAqw4s9AVQSCSfkYbepoYq
22Odq3zddMNQq5h2h4MuMCtjsbYatpQ07r1hm+2/G09PRH/ey2aoZUC0L2xG9iGZ
5lcdjlRIL7b+zqhZHP2Yn+7pUnl5NDMo7BWrgzzSrGeNIY5iOvkplk7pReLbb1XN
t9qq0G34tNzmUxUWYIGUhEL6xB16RTfFM1F73h4zyYTkevyoVh9jhUA/K8Y2ZgMz
g4Ujq3NGYX6vDCTjdd+dRKa8zOYQH/5BUAH9alYQMq6cJwHEcfbmgDcpNTQvPSZ7
bpdpcmHKo3TRh9vSRcLR3jALdUT+Dr5H8VM5sp9LUUirTpS0Is/X+seUZlHKQOWs
jw7jeXoHktbR/xveInyLm/pyCuFUvx4L28Obcureh5AHPLnsy4pOjI8urn5cpH5Q
Otxr0mY3NBDcpC05ZOXsRmH5VLN2/uDiFE7Ruk5sG7+3e/URSd4aY3o4vno4M9X8
FaAoRzhX9oDtnqyBjXa1IpcPDG0I+Kf3ssXLWOJEzzHenXEVrKg/jLLycS7ru9AG
+d7r0I/jr5Q4p6PnrPojsGIrif/yEcYyLEYO/pLDPynJduYtxvc+Ys6pJWY2jXQY
pu3c8zInkCuripyixfGI+pKEx7INjkVw0VAlXIjbyWX9S+znpi7YL/E/82mgnKtK
dRyx1aTQij4Kt+PokyDIk2Ghhb3p/CZvXRekhSfVmgDBfoOP2wHiXQl2MBcsMtDh
Dhrui42WMnHKcQY4RWXI41vn9n0Y5IvTsZQicGHUbburft56SmnFdfNYpV4rSBm3
hcz0hIpgu3Yc0nQ4DKIROtCBWrCwneSs78WQROdqGfNDN/yvOE1dqCtRkLN/hzxC
aiemW6x19E+sJvT5aiwJfwDl+8XCvcZEXhlFJKhBQ0wBKXymtEoMwSt9CjCQwddw
FMGL6uXzmKyGVlYRnQdIQNuceqMY7pPLdzmBjVm3sU1QtT7CcdAvg/KDQNE8DE/I
YU5tbNBMdOHtZm4AJ8ADnO38fSaPnOyQhOHp4KDp4n8OKi/RrrB4oQKkTj0AKV1R
k62ECqaZ+NtGbUZgFQadVE+PXTuJeruXQptRI3HgSh6ig05BouQwKxwFVJesbaeq
mSwH/LbfWxB2HxBhUVNx3oHTb3ReELahPDoTGdwLwfKhso/alntObFagHfKVxLh9
F8aXRXOGGWi6bixCVRH3BDFAXQkqTgtBFm97NxIX3BrjcCpJBe6Z/cHHWB2N1HpQ
xP51T73upmHllwzMsOCxyAh0+DeFBMKEr7neenrbrmC4itm3bflVt+RbbYLMVnLQ
B5JBTAOgkIwbyNkwkEaqQhomL3uf2gHkN01lUJ/Kj+hNvwWAHJpDxY8SsKl+GwVJ
/ZIRZKjLdANUUVtDexNY8Ori8mwXMjHA3bgAxVBCcXeYUQ/BsZzS94tRb4glKckn
W+TvpfvBjc0NrPqB66u+OAd+R8DZhIkWIoNUOxshWGM7IbtjwN7mzgLXrK7a31jl
U3a1d6yY+Ta5oXdpQdEtCr+onjm8aPa4fo3ayhObRk9JgR8T/ZYpTODicsQ+FXan
A33BKvJArNL/kT//6Aa8Tdk81lHEpkKLX1EoyZvCvYr021iktez06FTOjqcVE1HQ
FvuDtE/T5g3eYpGVp+7Oyd9aeFmOH3UNjPmCvjIQLQfCl2uYKphxYBOeW8ndtGja
br/4xfF2lIRysDy6a5nSjIL9PJJRYUJSG6oFRBlC+zTaxiaFEaQ/ftQLhu6r/pl6
ixMOfYAE7i91c1rrrDN6TVVkW+2Km1/ClqdyDniy7OD9guWKAjqFzZn83k1k6CNl
Ppe1l1GDPktRCm+cErWSNmPZlff6h2o1qjfm0WECTu9c2JnKXgNSC5Orh3DPGc/B
qbdZKJFrGEeVVr7T3fYsviLdKrvSMEOm0qZWZwkCZvzOyGqoQ/3jYhb+jlROnK/B
eT4cNK5Q7WXjM6Y0DfL9agfiLjhCIPr6zN2HMgqi8WFXUyUDuh7hnsMkgfEFM2Ib
00oXMslJ09UNnCXF1fCZQwjztn64WRvB7Dh6NcFyEYg+0iqacJLNx9i+WXMeCAzj
+LQG+BXOHup9b60S6Pl1uAxldAuNlRrTO7LR+IszsHTzmKYpMNRlB6U1fuezCO6Q
ayMx2bAfY5h1evkQHBEC4UOxdC4QkC/QT0Csyv5d5Z0DBuz5s5YWqH8MaqMj0JrR
BF50ywD4OlRpfLag1oZVZ5yr9L9C+XO0DEoSo0EaxCQWjao6qOyCPyEL5NEgkm36
uvqXJtSvfN/81oaI3ap96yLJn8N7Bepr/rMKlnARWsbdj150n335hzM7H64xOinF
mJj1aP1olg13aTzOmpKBnxdXoZ+qkfSR9l4cJg2BhBsg1BDYAFPrSLoubFFrYDVy
3fMv4Arvtw7E8HgLtYrAtogDYEnFgilEMdeisLrNs0N9yt6GBSQUbN4NjKQwJMpI
fXMA58CWX/H1UsZ+nBbvKPTFC5v2ERP+I5/riF/SzgtAbzQdw8TVXqG2OsdxEF16
7O6XmyYCHH8gSyDbkGRElpbL6Df1RdIQn9sxo0i0HzITg/wcMtS2gP1dV570d01i
Cg9rQei6sOWClK5uuCXnw7FkTBbQAyV7PPztjSVsY38bRTyurCKi7/AE6WmvgPoM
Ja20oPGj/1TWEQzDj1hZcGXvpdncbXvHYu9GtkCwLPWfxRwfHd+3Q3m4nKCmGzxX
LCSsdVssszJTL1TECVnirXFVC+w+QFGy/5MuKu6MupCsVko6xpkQglXIusrc0hBD
d6EkF8ZSPdm/gV1MCF9gZSMmX23Q273vAekDvqiSQYgcMJrBREZwrbVYq78v34wM
ZAsyxG/m2igWNsfCDI5zFkjEyOC8kWMQRVMy9mIG82oxn7vgG7iNmqnq1I1PFFPx
GEcRi4Al5qfVRd6EgteKqFrXUQiLU0AvzMXggCyPIKMRLb0phgP4XdCxEcunU85+
vFnA42tPZXREMZQRcGgmYqxeBwAFU0yW/Szk6UGdVkwEWlFbShIRRVAmmS/n8ZDE
uDFXB5vAoZtytzrP1bE4zqw22D7xWMVCRcNaFW8NlbZxtMxB9OCFUkiwN6tSKelv
3+uZTOFAbeZR8iJ+nMn8fGc3EdQ7beb1A78P2kgAp43ygQKwu2rUDCCmWPx9nIBk
86lwTB4yJkNhFqjd2IfR/vz9psVG8gC3nicEc1v7JaGSI2MPcU7dr0VkMhnBThHp
ox2nySCaIHDltKLEu2OUhoeIPNT4dhIoEgtA+mRRB4TSARRktr7rjxz24jAB8C91
zrmnoGZoHHSrnxX9GDTaCMVa2Ay4yKVnlaC76tcen6NkhLrt4YgDzzIWCUsoNCR7
5Pkx0uwfj34zL9Fp76utODEke5fbdnk647395EPH2a3iIt9UO+DxYuUeWnec+E5w
1AVPWXx2T6+yRETAuwLZ+Rn0d2HjT84qeE5mH0Oebs5Z1XrsJqXbKs4oQLh1xhws
EfKpOd8U1EX75uDXyz9Hyd174rFVpLDvxqbFF9qqRen89NckJlKUAH/fWgEfMH1s
1P0HrW9FLbA7tAPrehLoFmNRsZsGE6teONBu8MVkKbu7CkIkpi/ukp/CL/3n5WEW
9t6hfiVj7HAmi4yo4LUmyu2J6K15l06Le01yWvW1ovYBhsf7XVgaFt+6XqFRWHyV
KMI8zdNkfH84Yi0XWIxvR5fsD0fbuBKPMrmMPIvk3chihg2y9vs8O3iQZ7ZRIXsu
dcJITqDX0pqv4gdMvoOzuVu0mWgtscHjCrhYiJDda8zTjJtGLQOZzYNPCZOKvh+2
ZWUR4wcoXhJd188ZYVxbAiciA5PND3Tu1u8ez9dMlfqxc+hyLXI8PIUkCEp6GUL6
66omw5oSoIG0MpTrT8X3g5U1AO2p5EOdBhHVuHcMSLrWDMZ8u4bas4CLcaAI47Be
RMRP1dtxFp7b6W6DGZYwx2bA+clJccEQGqAkLIzHYnQXmMWc6bre7ma0QzPqSpzF
Oc45en0sC9bUNHrAw4l4sZyEJZ8UWv//rkPKf9+RJI8Omb2KwRXygmtDjnWvobeL
znX87Gw6i1cm3ohhLZgdKRqs/lu2pbHDK6R+PeW+tezh+l+/0NwX6AfyVXqEblO7
zN0A/dV++OTMOAjPRhVbzFcdhQ6BH5+BHat6NwUIPcvU7FCPboUzAVyAxeEzWTLn
9nATvw8VfHIpbzCd+b5Rgs7yxEDD27iyDAQ9gQRrxRby+5ylbcELF3Qai/wyRoMr
7E8S6XVtAw8bTa0dYE6xXU3EwuY1aTsg0eT8c88pHF65MR9/YJhejh8MMdYPqHLl
qT+5eXHNYw2obOXbQoODsm944y7eDHwa4XPsPZFEBnV2R9l/4SQwQPpHV+XvLqpy
ZOf8auHjeU/ahqjr5Wiq/5qGXWxUTzjj7BRjxr5IAx4j58+P+2eGoIkVuwz83p7/
qFYymnIfT0F9ZURw3XLqtrccegzAaBBg+v6ddPmkDagzBLRoamycKekvzw5mSokN
TKV/LXbTOFsFmqHtfvqE5tY/Ogm8u5IuYAejfxoXE9z/Lm4nDPEuGroplAwg5N+Y
WxIsIfEjqdFxfKJgX3ittqeciwOVg2HaFkPsiw99H1fSEno7nVc5i/vZLbuRygW4
k+IMVl4gy/byebPXaTeDeOUZySiJrGHQ9pdIDmLJcLhjZLNzDkTttXfZCRy5cgKo
PwZx3A0iNHNLY6YpcF2XINMA6CiRlRfjWkQW6nBvSv/f2JCXqz/2yq2ToRQfGsLL
TCHm4/T9bsiYbvkcuOu3ETsvzRMAE/X9ka+xCO+nqX/NqYmWBnKJ+8aFgnxJLiYW
Xgn52t1v1mt+okRzVfD6+s2oMNh03Z6D87HnOgf+px7dePL5oFRydxStwIy2vj4b
4OCQw/bzN0NITm6a0HGnrqF6lTpq2NzmyDSXSiM+88TlgXdNKH3lDf5acJKiy3KW
TAwZ8IxyKYNaZFWKxIKQZYLeakF2Rpp8P8DQmFso/ZH/RBTiopMbQn2KVYT74l3E
OarJfhjehmbGwaeLl2wUv24xsd/Ef7MLmklszEjqcOZrrHwJy0fhHMxGQo2oC4ut
ooqAfzEsxl3GC3Hx0kfEjWRzTgEHMaZChQcaL1S+BrOCBrgCO4r+iLs7Tn4GLEGY
ezlsMT0EZZ23cI9WEv1nRD6Bo4Q8xYvzgZ9DMClWL3pTVdM7VmbK0Qy6e8HlmcXe
ftiKrh7rGbpTe++NUIfJEdF0y5dOmUgz2SZZLP10hYjCjLCSGROTE6VnZOEytqpH
qdX47K1GSOUZayxYbIuYRCZ7y9AJBTUmXT7AucNoc3TdRLtcc7E3gIu5vk+2d7xQ
FHJ8iLxcgsMPFsEmKPZb51ysVVwiY47jw9uaf/hPyuKmfmca+gpSEijddTsJv4aj
ODNj+5Ow8ZKbxYJBLxEdPThrjfXr1qjMxt6sVnidKz8KmIFtH30kCmTNSmPxz7O9
GCFKdRlNdWBxYvGLmuTiEHxFMbBIZNdR2yt020zNQWRe+xr5DkQ64t3JfUSpGjox
bkvSpiFPNC3c4Hh9MiMzEjYYa/LWz+Xq8uviIPEdYOvB15jZ1WUg4pRl4LI/xFtK
dKEM7bpYtKPMVcJ7Vd0B/LbyIQgXZ1rO6fZ1G5QliYSVQURXn5KjF/NuAModaHuI
ylOtnCmRIDZ0GyXgWLg8HPzufKg7O3lxa8HR+yyTkDM4VrstFDz66CaYLClhB7ww
g7cAZ6hGhN4TZeNJveQEFQ9nP+Bc7bRhxGxWJLXXsyHpz0gtYCels64Sc8hoq2d6
jYeSz2ot5ifjVTHm7jvz00E92MgDSRLg95CmqHq1a4GSqaqzXvJ8OkBQcLZ0Xkr/
El3JE7JZfM/k3cNoE0nNmoxpBbe6Q07NEvn1h8J9Ez0CyKNNEBLhx0pDmTXQOItZ
Cw1JO+Tdm0Xu/ZqxjOy5SaFsWD5qPCV9P/SzTEXEtOuNbLRTXCwtZOsDJv3RiY7i
ktrhAt5hBt/81sMhoecdKTimwQex++SbJAQxeLakz1TejhVeEdEs4k4EyduSO535
3w1+4cO0aOZATAXagzUu6tmKzVQr7230D+xhFLT3F4k0+QwRgVLYHYMjPLzpyvNm
A4GOAhLJ6yScgapKBuf62RhuZpJ8FYeIvx/dHQd37XH5vYzTSHNy01fvyK+bLLHb
dUmYOV781jUdpMcbAmGVoN91ilsQNQTLGd97ZfyKSUGjf3gh6U4U+oe4YjD3ItJa
nnqIcDyIij9xwbhRZsR3pPjZmdO9T74KezqPvahMy1tnsNH+ay5KxrH1ttRycEV4
GtJhM+Bm6YX8YpQUjRc+z2J9tiJMrItqw4GyY7K6xk44AbPnCVCWLRArKqwEWr/P
QBxqAKPd//swdS6AJqdRBevZ95yYsHFep8oUbcgcOm9us3smtHccyy7Hc41WMT2p
kIYDim4GBY/sT0eOdJRZ0jOtx+SopsLv/nK0Y+aU/xAkc81pWeO2vP9AUMENG/rG
VlljDYQyzcOg320FsPjQf8yNiceERnNTHDulSHN86ORT1TuAKUifQtOGlumrV3vD
Qt2kRrs9ZnGW19WbJI8c9m6znwNtZx9vUu/pewZIrOVFYcw199E42gAhxmOJH1GD
neFsdeHV/Up/IVm7G07X5zYOlUGpUzMWYCWHX2Jrcontt1GcBvqGhrGaCGi4wFiK
18K26zH2vQ0JXvz8e4a+DAtd81BcqInLo3RcukMFSzrtqNZIJzahjYBC4MGxuJ/h
82Ext8EtivB5DRzyiv4Ad856/jtjLi9ONT7fVCBxu7ghOnZIes0FEZAFQl7sH9it
76y8kBoXXjn8qR8e3L3vLPeDwcOenxaQ3ivYopv61ycMzcqi8Qy8GZrcZUUJx5NI
dRFT5GMa4YiBUazGmLP+DKEzacqxVpL05P9oDqouDWU8gs//JmVsp+n3iWGJhYR9
18Qmt5UgBLJiEkpbQrdCPfKWakXE0h1o4clpvIGp/9IKQ0qmwlUeJyHOwwPVr+Nj
VJTMd8k1HvCUJWglCRcseeYQCYo95W9TdD1hew4uJw1DPWX5++6yWS29qJpZE1fQ
47ijOfDgvzJfmt0U577zh7Jtrz/TUuPNJj0VEnVW5lcV933gDMCxIsrwsZmxwcrN
NapJtcv+xiSUqh3he58Wyw9dU/xs6CChzDl0mhWvtkBTWQ4N7hwJOC/aTYOyWsHd
qR23nvFDXMA8qsX5lqsbotUkUmA02Cccg73Bv5z2MPFdw8CPBOhUXxjLXKe0gUZp
N5PPpP5pGH5NMgL/Sz8CEehQ/YIt+EcmxGWCD0a8fyhoyHkQ6bw8yUiEv/TUU2QC
XojaNMVXaQkzKp1tR+fzntI126aSOVSedZec20RyVxCCfL1oT8HUxVlQHHoFDO+y
2KfJI3ezbWQZeVd1Rp0gtvV94HaoZgpGHNzOjmv72EBBAv3jaJQShnazTpdp4EeP
SCDnPC+ZpT3siE/eXhEa84qefJKrL3n2fNEzDsDRGTuSe5TijlI3t7RMgj/Ec6hd
R6KyJBEzHVujSV80XuaV0lupst95XV2D3FrwQzPESdxZ4Dvrqy5JWFHUbdNO1N2D
xQs+QfcFHk1spdl+JCq1y5ZaxZMOgEySO42IqF2nIpKl0cTWwVO02En4evNZkbHC
hTj8LPXxN8wCQK7ur8pLyexRri7N5Ik0WXtxMUi7EGcASwU8Xc1xW+KP+Nmz2Bcu
Wj+K5xKRSLLHzk9jaOqOtmzlBmDphPvy//zvqdrsaH7LoOk+n2BNU0E1K6MtMnk5
dPuCSyRmjBQPVIDQ1CPH3oOXrtzIDvHr93RRrGrIvAhPBxppqSc91mb33KAb/aDo
eCAgumWIN/nvs7UIgi0MxG74aGRVbE7IY9yqKzW56AE95nQLx7TiJ3rUScSUkS9B
ePrtpjr8GqF/Yo+d+Pz9yaD1l+N5+h1wneYUy8TWQtIs4589FY2ghN4wGZdBCEXh
VtPU81znm9pFwruX9/sqhGgi2gduE0ZGfu6W0eDXQDFJ6+HoGdBx7LKdCjl9TVjN
bAQ9+qa2wyVarHSvTrmjka4WJ9AzElQzoq67o8XRE48+3xY2mew+5jxrNay1sMP3
2XCSEsSp6no97PAbzE3cqpMGaOMhNgMLJ5SE36/t0w/LsNg4fQ8YWdv3Ffse8ZgJ
VQVn4aItnC0q401Wziv4FuupoL7Mw3hD3OEp5fbxaUlOt6Rq4I8zhBLJUaC56SSz
lrJJxztFUKTlnFK8I8B6ZKBKhGrL12d57cVK4pQpj+t8uWoPlYg39jc08qnME/mv
S/dl6M5a22ulCWtUf9TQpFTzLEsriXCyRPSEGKTbG+MPhdr3/Xij3Ow9DD1vd65P
KmqcLfXCp2iyREIxmRVs22dxd0q21cDmXA/a7U4VixtDsqGKq92Z3KOAO3wGBTan
7t2iYyVDaiYcEifc4d2zBNm1iJ8NmbpWVsLv28DE/H12DPanj5BWcvHxNg7NPfbN
SJlqV67O5E3tA3uSUf2vkL6ijYwVweXDIsZIt42SJBbkzP4kVp0bA17waDz/UDYd
X4XvbVKvXZSGD94O6xzQl/wA61hiJBRFiEuE2Yq1I51VstvQuFJNvTYmwb8Hkaf3
R0UhfQ/M7JapgVbThW2//GVfCzCclWxSKtjmqlpstu/j1lFmQte+hbTS8KMncSFH
tlDXT/SVM1ibovJwPdLlEGDG+dQWOsg/sQ6BKtaASyCX1M9u9oG3JSpgGIeQheSU
aCWVZM0e2XbgrDTxwg4I2RtfmMY39AhdSwzzmxHb8+0UOyvspQST905Bi3RCfRTG
FgQLBy+UhFMMCDFSTB65xmrKpTDk0guodCWm5uuCIZh32EYJuwmGI1DFjLE8OWZ2
TblFi8PTrjeuBP8lm8Qt4wHx3egNriiYdCaV8h+DpyJL8kOzCi8vwJtkAUhDq9tO
gsOshEv5W/kgKwzEzxkUgP9vyD2pfSsbDEN1SeibIrEO46SsXxx0oUl/Afx6IUHc
idxtV4jsX+Lp/dwQphbL4uCxW1Tzr9z/mO/zxP1sBDPWbormkoDc5hm34PMIp+tl
UeQJflTsbSl/X4VcyhBcaxeXk4dOQJRKiioM1Kii9aAawKkcUjSwNRbvlB1M/6dK
ADQdmcRp7OQQ4NkOrNH4twIor5mfzS/9IiDsl+yM9tpnHaAlmhovU66Up3mwT+KF
rD5ySV2QUcvelCahk6fu3a9igTaO8Ovuzi0XN6ianhPfwf14UC4IcG+FNo9NCV5F
BQ+R6F8DpMmlCaj6ba/n9cP6wQotI2EICDSXGeBMFwQWmB+n83qfcIlhJggDc/dq
DGW2fZ8ifb4Nf1+JSngjqI18eYFsG0CqYX8rviMrVt7J5vObmzVjDiLpHP9BYxEQ
hZeJQr/Qg3qKUZEs00gD0GCncR1mwbfwOxRh2lOs6IVUfRZ7xfUaGdhyQZzGOE56
yfDxtNi6+9KnhTnLSvWKKtsYXKG2YR/9BNPBvmAHBtQgJbqK3eHuhI6paUx39/rf
r5/oOoLzmuTwhOpunuWUDDZ24wbU9BSzWkl68Ga0LT36aC8uK3dwohKF1lRYJZco
VUaCo6d3u8CxIs7JfsVWpqmtKztV65D/4iS3bqOKqXPlJcoc/bndYaX1mUDY8Gam
ylt/BA/wAyYbF6hqKMD4iLEZvhBNQH8ICGHycxzfaq8y8EyGYd7mtvxDeJm0NtGq
gxRN+dseJMj9a+NpILqoe5rP782ClXGkKv8EDBzHRrmu5oyrY2mcKwJ0LEW0ibSf
1gDwoyxGx1oL39ew/lo7XQv9S6oUpbCRDF5QoBND8PnPW0PP1qm9GhokM2isL64w
mcvYcNiiiW9S53BQ+cJlKizEcxzAUM4VyP3SgqY3/cR7351oaASTk96XfrEWn30e
UGvpys6WIdz54cTZWc6ZlPB44oqERY4nW4f3aAS+PEVYV1K1KcagpgoSbBs/Bw9C
ZVfjbBWay63LkTqtotXSbzgoiEFlokyJqskOQTYoxV2nShByKC8XOFiQCv1TuKXb
sjqlBb2U1el5kjzvhb0WN4IBH7t/eXRXPehZQH2MnRouWpiMX9EbzFkOs6IH0qQw
qAa+ZoAqRTvD2XyYHEe7uhVnpTJfeFFsHUPEUsACpLWVjlzN1vZuXnQCFf/HFUOo
vJfJjtlT6XpjU4Y/l7xCji+hfc7YQjaSXEDcq9Ch9bh4qibXXiZcoOFY6en058dt
GieCTCWkQx3w4xwGUfRYZnwNlePyKd4xD2kkmi57HsqBbtgwXyhT3e6HwM9yEDA/
ND7s1JF27Jx2tGznBYkjhuBzLUNYvtpduj2/vxZWz4kr4Bc/9DyIGJ3hilCHrUB0
LUfJaYxe1dqwFKt8AmJD0dK0KAcLTYG36CGMizf4MAmbANy9BnIq8gnShplFZrfe
8lLUkOV0w6W82WRiWrlmPeY1Baw19Vn/uQiBTL23UtBU3hUEbTM9HBowSICZ5vc3
yHhKYjks2GbVfX8B3Xikakj7bRA2AqMWSUEixV1SumpyqrogzTaQVt8LJVWTSghR
pm08Km/DQJBokraeBArkqWrg534aVSoknkxqI2DqaoSTkkxUrOAW5TqPFQqXjDDQ
t4GKO7vs2kwJzocFkOO1TvVDr+1kn/KMWtgDwQPXqO2QikfpkHXh37ZkBnu+iUla
z5SU6POMVU0GIVxzRHhGZP0zREjxrtwgyo2epkmwZPzmUwAX+fmkjRMt9oZ08kNC
JDbuRp9JnX2Zf1hfNeUuI+EdN76PhNPCzzifi9hsq7ccpCC5+qT1aCj69G+4Tjzy
RF2wOJlmNs/W2tCJ8x1XceapmmRQXimyTNeLITv58jkmPZTU5TCMtzDt8rcnIUg7
iWm4Ec5c4QqKrYpRfTOiDV+OeNKvE8vI16loZazShdQYrqK8bPosTZQrUTIS6bqN
Ywi2aTMACwG+MewqoehLlS8xW1Fte4v5SEF+lfP7ERYbO2ekkskq2B2tclqZj5wR
OgzwA+VuczDzmdrS7z+HUCU6HvQ2P6lUE40oCn9KQ6FMuHRTkLyXE5iRWoDJUjvm
Gc1QSK7FvfPQXWyo8aC6wsuXIIfCfACXzBMKDAOIh1IGCj+eob1qlnVYpIM4TDgI
/8tltByORC1ONdobKLkuqO5sswyNsVe5MH5jmD863JPgUz1D1jfYVh146tca8/7i
sr8rX2rB/BaS4++29RUHzAseTxEE3JYMHXB9XtNzWU3j4YA6nBlD6Kx6+Kg509PZ
+363myPvNZHXozHbX6Rn7Gq5amRE6cBIi5RIrmXJORNIEKb5BtipVBt41IWJ89zb
UI44TpaCGwAJbubBeGqSXbqptCv3edBZ9GdAAIbLy9ssLxj6BytjWyt/J563ozc6
mGd4d+Op0z7ZDdVp1lUT50r7H5oi9jGTwd38U66IO+nUf/kYd53R2ZHku22Z6YEB
CfMRpLAOKId79lzM5r8beUHStBuFy4nzRqbcrJ3evjpv/WNDirT2s8sYclOOSaO8
KIE25VFeHF88MYOckV+QRxsCxPdB27908hxP+A//6HSQ0E6c4wMINMUPHWzIlplz
X/BNamYfrR48mwaMWBk1xZaPyfl8Q86/I8kVTDoI2LJ4+uhqXumYJ65IyXnbDU6M
ZA60e02MMvaSkVMAK3APov/Kcr/u7+tazzIk6v3N3RP204qtWbuPZjGtDWe44f+k
C8om3H82f/xhiNewZhU24ekXBI21iGn8q1MZPwjashaL4d4EtiWTjw0bUj+bOzmL
5ugcvDlqN2xzDx7MxA4weJlcnuz6UCV7s+n1lu8OYsw1rp8OnZoVNygGLjxKhjC9
B8hBlgDWEZWj1hn34s8df7NRKamg63LJmfiKPnYa1Dg/48gqrRioW6lOD3arERPP
8cFRWbt3Pdis31qE2OEpJ/Wjnht54832PRNDfJAKIVsy1bs8Cw+Juc6f9IlbYPq5
yPQfO5qkPu9wYba/2wYIGQQQopo9MbVmrtiq36if+ufu+vT+4DWYTZNYT1JjUsjd
xYYt7FIzS+kWSUavYb0uJtGAs06It9kFjSvLP7VH0QU/Xv9tf5Mm858k02iPVtPr
FzlHwnzbdKMdlJn8bKo502UYDjAHKsmpH0CSCjxLEeIWiBBI0QfT6vz2yu2PWVuH
UrHyDKjmazeQjkkZD9HQpBPJ/SJbN+sa94eUkTxhCjCGHd1wQUU6I8jl2RS4gT/E
jMeoJ0yD136juHREPUqsDfjZtos2P+Kt8ew/44EaURj5xUVPE6ulj1QmLMFdGoko
jzkptdNAYVLL8+ON+94OH1spjK1LKm67ze8d0Ve821lTdU1xkGDpeTSUeDSUIWK0
FVs1ZbNb5cx/MMcrcdCd19r33VX16NggudlRkqJiHh07MODyNelwECIujeH2GoSL
zk1jYmHVhyjSRFcRMzrPAceBVB6gg+DAfvOCLoKqXXNTD8m/ZWE1j17mHKiSkGSn
e+G+hYdPxVi/BuFz/xv1Eu2RxZiVu3jM7UtMSoroLbhGsolnXdehZ/MyiR2jYMc4
mFAe6vtlOEN7YvIemsTIfTqLYkCNdQQ1gzI6/fpgJGLqKYfufpYGbzjPqGERTRE8
oIytbHHOJHcH6xut10+fetndXYqbpKPauhDOjG6rgCJOiNKE0rFrukBx4UxvlZXV
34qp5A4mnU/UpfsYjBEqoetVfTOjfRa1951WxifnaUMtIR/cE3Pu4Kv0oBp8P2kW
50ca0PRF131zUiDyACYDplZ3oHT/uedfpg3Z55IGubd6OlmUaR5ERXEaDPS5cq20
q4ijBt60RiYWBkfPaVvCMUaqOhTC4lMd0CHQyXElqDquT1C1xLM2YLCGI2tM5LR2
3OEgG1txd1GNDfrNlpHsk5ITzRNZuz2OPGccQspVwKNilodXld4nyaKKXvZwxzX6
isrCIhQZ+zuKVncj5vFLEgrlhmWzlweCegGk7sEsZid6xwKbC1LJZbiwDxWNW26W
WG94ekhlBb9pGlWD//Cz3LBIq34V7u/mNdtd9BLZLdjs/twaE+sShd+CR81Hg+JD
1p0xfsbKgpnHCQsxwti3/upV/j/9cCW7Y1E6UlG4yg9iBbhpy0OiDKnvApngQi66
QTjN7iAjCJGyj/6D+gKUpZNnOJnkF2zzB1SZD8lMBkvsBc6MKeY6PNFF1S0UNx79
CfdHRW73s0rq9nHN2FOxDTXRXWJKCBwZDOIAxVRI8IMjN7tgcjtGHKYas+mOYptO
mgxl3tVcIC0qXRb7/0J4XBJDiPjvh8UVxqvUt2RsJMQW2tWGVT0YDWuwwr8AkZ6u
WSmVMTvjpkfPAlsbn+LVB4fRokmrG15Zx5+JJ35HbwcL03Cp1r60PrEBf9apqbB9
0kSCHLOf1K91LW0XWEPgSlZBFXDUF3RJDNBy/WLsnymTMDIezHozpNOXsAz0VUXd
X5JOb975+uSMG9iBmu4b9a9vDEg2rkfZ/ucpwv3J8ATveHdb9TvB+plsFGlq/Ajj
H5wJTuLrfIOfXtlHRM79OK9+TpfwNWD27jRsFVRl5QBw2aWGqrR10Oq4i0UdOnEY
AOGSO6UWMQaLnSp8paHA+ytUz5/HlVT7Z1fZF/JjiItRBCR5C5tgJDfCQGp4mAUH
w33734chsi0F0g5XD5856YqbHjMReQyipjdylLAwTJKo2QmULnNOwU4+xHeA2mY8
K7YHXX+DNAJj+jLUYUJgzT9x95bFSYUml2YPemER2Oo9TihUtXThnw2vJE18TafG
3bxqvLoR7xRPWe08ZSDyzbtF8voZ4xE4u1XbmuB1gz93jAByJwkxvaBOgbFOokYz
0xBxTSXAMXx8uWOypV4AKQ5Qm4pkdApHvMUXzmq0YMS2vWBK/kmSm86wE5pAq87L
S1z4N12diHh1IHQcDz7ikTdQIoxVSR59S0Ci4x2pW5Tm1oSrrST9TzXy511SGv9P
olmMZ6W7Au1ffv3yZzvg7q1Dvmt2C8O/9FNx6YXyunTQGvHwIr/Qjw07bGTvPFnu
2NRS2mYKMGK43f7l2XlcODEqTOTyk+fzhXg2uoC0fAQNrbRleX/mid3cmbKtAyJ7
ENBBJNbynwHA4sQqsLd4fHfvMmTX5DmAssh9OjmMA1DDTdsW9v9jFtLIyV9wAmfE
vnFQfN/NJFDvvahuku+TfJVhAd+Ge4uK9UZOPQnA674xBlBiwjG4UutQv1z7ULRk
ny4N12DKsnljNWyU+v2paNWU6pfV/9NZV+qwjFLVryZcHawNK8sf3nsxSQH+jR0y
QcnMKN8TrS71xS1wu5MMtAgDq3c5V52pnKktQb34EUIRS5RP2T5Xl0Xdz8ODiyZS
fafxlQfURRQIMLO5gPYQi3h7JoVI4LOebZnLNdZrlA/ie/ejFxWYGh5OVjbEbCO7
seeuCzkkI3CJro2ie1Vu1U7nNeX/cqrU2XeI/0mcD+FMvophXyiJLdWenLtDiUM5
idRuVRXjCmwVQnuBtovNRj9v45BQ/6CyDCw2H9H716PpkAmZp+kve9DfkWK9Bm04
qwwUBYEgvPG2a9z8mSMZiuxLQagiiHhqfm9savbaA3OQwjtaV3Rf3CMdpgtFy5te
DgitrZg6WYh+vZA59A1O5MB4Uwt925ccHRLSC9WUbNB2um1UD6+yLijPwzOcMMsG
7JE8HdOCBvh55lka6SU+S7/Lf4036YZjyT1yhqBUulDMisf2q8+QrGGrkGR5xzwA
jMN8ZsxYBaZhuiQZNxm2FF4UzJuPvj80xRUfpnWzB975eec1NnUDYwSwsJK6/dE4
GxHRwDjhVSQRm5dw1UV9Eb1UBdsm8qatLFHjzI/TuJMPoe+EteSVqrjfnKnHpuSn
K8eo/VQyVEscq4eFPWuyFNXz25nrm6bwsQzOIJpt7VwShORsLKhIktx+ZsZTMyKc
f/j64NbvG/+Mj+eycb9s4nF6Svueg82GZu6RPVpT9cxw14KS4GwVzQNSoFPeBo8+
DFiYRvakzaIGMYUZB7zJn+pNPPFNJkQrIUMmBK6pJh1wVhPjtDfb7yNQ9dC11BNE
j5hwYZTAnwyXCNLrTElGSQwFL8qBL43JrFF1/NZKINyzFims0wiO9Xn18tXUFnfy
VL9PmFOPixBlbg4Vj76ggGd82bhmIVjCovFcIy8ut1Hz8AqreMrRgSsRjdzzT+hl
wubIYXdIXR45JhZmkw938KEjzNHNVWSrHH5gOWaq8BauRd1q/zuGKZrwvRQLCuzP
3QZ0xIP+fcIwDQbYTv9l+oKoBWROFsR3IbXyb0b5BGdRNLu/0mjACK3rLsu1+hOe
Et/OgtRT1/cufAztrOIHKQZN8W++3tpd6XgEwRzmdYivKK29qPqZS5u18jppJDgo
6WSbyuI7qksrg7+tYn8mcEX3+J+U2UBHZoXBm33ugN0MhrfQRW1sQ/Gomjq7VHbc
u5bPt66sBdTbmYYO5U9/Ctmf47azlhYybpdwvwwC0LjGG1+2endiWuDeG+dS1kNs
rLVQs6yfmIfA9fAWC6ZYujkcWHqEatqeX/lRywO/M7OrtyHKZTfuq7NG1QgeN0cd
z88avakAPDDd+oPbp8BmEpfd5hae7fQgAdBFWGwQOjZN4M/kZhOYNLCLyyMMaflM
I8DZtkY2b74d8YOw01E7gk9xXalGF8DqZ/UYTnqGGOPX3XJP5b0o6ouO75y2DGZ9
lomxn5lBtaY/JckZnA7W84nklf0XrTz86EDQ6HRRZSVWPgKkGGwEHHT+pbqlGMr6
cRUtWuEwXFl8q+cfya85zTYfRj5MDTRmYFsbNd8jaQSCdpax3/V+peDeaecUokPH
j8c9B1AkuSx3eUD+W4kXurizooY7Xp3dm9WUUV9vIaYWTxWc292flObTjYtkBWZ1
+BeSOU1ShvxZLJtRafU8kpaVIbUC23+FisjRJwixwrm2tAezIrwyl14eP3vTd+BU
ghmkvwdedC4UqG8FgJfTyAYHqwH8aCdY63nDUSFiUqfPb4t1yePSuml5xlPa7Idl
cBiWrg3BNlvu9eIsguR2152i0m13j4ueqU+JK8IPEAKWwpSmuJOPzMLV+PmQUcTE
mTN1epy5SItNvZujBc6nNyrLQ4CqLRRjscA/KjEj9mK0iWDzjPTBldWV3ylIzjoJ
di/bv6G+BZx5hH0p5TNZT/u04voLaLhzB94ktshuYDPIOyoAUouLZId/QQr2/I25
R8/hQ766W2i7oAvNV54MgnKSlRvaTe3XLJiRXQUW0jTBbmU5xd5Pc99xcVq6mpce
B2bpQE1Ln7kSGKw17+MN4bAi0JgWyzHT1w+SXIAoQ7L34Nq+d+C7TuHSe3l9aZ1h
tAGQ6tqzszWMyN9iV5nkAyEabqRNazoiJLKBPH/wBHlQrJze9b6+snaQjQBLnZ/B
VzU9mtQP/R8o2FM6InrvoUaoj/1bTh3dx+EX2IAh8lKyu8GB63xoBZsSUvrrVd8W
YvDVsOxzMjpe+KmqTziTiIXfjEr9xbaDlfVXlmW0kvXLyGcW/pBYu5UUZNA4+YjW
EAfehXdUhxX/DVdUBvE/emCXfwg/FvbINg1gfXx0/om8td2+G5VF8BHmPkzCpPJD
XvHCAwxoXl/uKvpJYDkH2WZTGPr/twfnsu9FeSTKrlrWoLZ/y5I3ioDGqn9Y8N/B
ByqzHeXgMo9NWYfM1VLHmVsEmJtjM+tdy3YVadE3Zq+B/67UyBiiNB3hQ4ERhUlN
leUpUe4dvIMyLDFTHWARWc+XF7bkxoTHcxrd6GIjE+vIuLwoq1FPH3jdTsiEgh6i
iigFOBOdRNgfzxXyz9r0jLbg70N2XPKKeydkpHGurYQN1dZQMOn/PB8hSQLLzuc1
xpVzwBZ/177NLbFTH/nePZmHePpUsx3IgFNs9qM2GV/csvd5iTQ8IovCdsi55dNz
x3nBNGg5n9qdB8a1CCxaXfpVQi9x9sgbVlEtxgodu7sLhBzG2KO3pb4QCNnzwVMP
TQ8+1jLoI6tYQ43KBDBFr0pW2TB8cYHtF6Poo07yeYAy5htT0icfZxNjO93CcWKx
IPQ3kC99trAyMv6aCt6pfeXW3NgQPWRj0gIIB/dJ5az1qJoJuoLnd+MNXq/CNIo2
EWjP9NriNxA/8IvHP0gz1SQP9gTwiQiLMktu59mFf5vIGL2sORVy0dEDOduanRxV
lJCs60sDcQxqmaTgA+9nRRQwWHQBfO/foOvxRbeyP3ZKwkkRdR87alf8QaLIvgfw
Y6k1lYFrLokpJ8OVeQI15iiSrYxMO2LrSrC3y7sPSvq1WPcsd/Gm1AxkcQAzHPdB
ALtT22Si9Mq8BJV7E0qBL8Z4p2iQdhiyLnXnIiQjhQEc5fS+n0Eor9VP6vIDz7WX
1stTgJcf/iq8NyHGPfdLSIeewSeWX95FR0CHHjdIByJZFCF/Qk1sKl/9PzLkWoD5
Sd9Vni47yXcYMJj00gbJa489QffkwnqSc8Ilzt56aKDWnhaWhIKzhAt/kVn88cnC
57J/gEH+8Tc94tXdbwViQDEocfiD4e2SHP+WI1fyZmhLzDwM+8JdqUQYRU5CWbW6
n6HJUHgwQ2CE6FvP2ZIgHHEggxFyNI8XywwqTFCw+owD2qe+nRzdlYW9OtF//Mab
xuOwpLrOML2SIrcBDZiBDnt9PMmllUJaZuNAy1jJeKYrgmD8z8ixWzeXDfr/1jA9
JvhLl8LueQTOhlHpRZHPOe8QUlzgCSYB0hZxMpEGfyox616OOi7CHIr5zIlz8yn0
eC9m+ic4hQcMNYxibEhZTkssdtdp0Py8u6NnwMCuJkT4DZ6ue+tqtmPIB34IxKl6
M+AwBhyQi2lkS1/Hx8TRJuy95JHxabNoJ9Ix6AZw8aJoKGaJngYKjJJvqP4GSdlB
FuwHHR/q98/gUMdKv41wtptXe3QUNrgxjNXHEsBHsLWbgvoMo4Ge9E7JAIfn6WMn
3g+0D0AsBNjCJtAtCWibo+0AoOJPAMn4Bi88hDRkwQnmRAmBeZ46/jH0fOV//Juz
VDJftuPFLXIVX/nS38S6cKAEFMSZQ7uEr5bZeNj64q0SgRIvHJ/r4KPfdyqEeS4i
1Q5Bsg9g1XLx9v/2EmC6JQbdpiAtnKMLMAgQ4Vvn2erFGa38G8+fjfMG/LgkmfLf
JErfYROA9NQGc8WaI+zpa1eztMsE/esxEF0HZSxQRVkwvN1WdOEzMcKg9ZWJmCSj
zoqR62doujeCI6T9TgOzetKqIy2Zn8NNHF5u9DSplqM3oUEIdmrIvpwEympL/dzb
p3QYxdAk5lufaSzBjC1EOVkOgl3hs5q5YG3yuZwR18xvqwU/EUtObO5Wxx0Ldj/D
Ygoq0axJVFOZIKq5Z1M9j9lM3OcRQvL8f3H4Hz6X2EdPIuxbOo7O4yhPH0HHnEQP
E9jiETh10IfNa/EZ4rMW7silhS0Npx0LYluKPCzmmEtxs5WIbfwkVmJC+0jJfH79
AtDUcUQtJiua2naIJyQSmLUUr2Im3QqFi4r3xla8oMbPJrnFvpadJpjWPyuzLLUI
I222xb4FWCZIc4eqQC7jGpVXzfm5sOC0YoN90q0cwDe65dEmMkh1bwzjHhp0firN
px0HCKPRKssANkjJOe/ZzUjNAq1mfZhRDUSBmyJv9YM08NaYl3NqlsHzVV9gRwdh
IT7mTyGtb2aCZb7q5XzCyX+LwlD+N0HlgZlKfukBao77kVZqYt9liebV9D8H2g1T
TkZjpPAgwN1glb2X1uYxF0/DGHSrO5uCs2UTz5hXEYtGi6v10kgsiEJcohyEU26n
UrJwidqUM7TVf5q9SQ5TSp4WBW69mKqXpiGws4mxcb15Nlxkv/l3+UrS55ZXt2Va
cZenlO6vFIvdY7dJZRIipqXqhgYR+QPNjNdqNSTs0yQ5DVrnBtoDtQZJWsGFojN1
JJphidRxTaStQT6k0j5ab8FMaDHpTxlFmG0kKbOCRFywGZ7W0x7js4LssIr+Mo5H
jET4o6xOT6F1xlV8BVO4CvHaNW8KoAEgsPWtC8XvLVNY9fTw5bDVivEs9ewQEHLC
MmMdBzgthj1TFuiqy5eGeIdfsz5PeE4PQJ9xovNuC3Qs/yb8YrM5CT1XWpCtCgzK
HYi7MwcrBYejq5afQU/hObnim2pBQObSWLzATkuH+hsc6dn1+jHW4NCGoXwoOlpY
qyhvPIKpssnzaZatqnvczVXat0owMxOKE+u55aEXMwgQJP0MjRK+dDteH7MUhgho
rV9z7HcDLpcn0B2eVm/LpuCpjaJ5beqjqELYk9SHJySlx9YLhoZ1c7h2XuhAy26o
aGmRVrmgjgaVB8EaJ1oPPuxJG8nNpAs7HsWH8EK8nf5XL28jIBeB+GPyby4V08Y6
upFj+DaAP+323IUlZye1d/oNV5FjjPEhklNOCJezr2hahkllpc7vItw4bKxpYZDx
EpR6n9Dbb01B0mIZHDESlU1ebMcRZX6QUMf+li7hDNnMsDJ8tZaby8NF9WvshMXX
3vy/z0yvq/SRJuJgbKh/gn7G5DnGO9UXx+DOcC4rYM2XhIBTCGEVsE4CvkUOF334
c49K61NalRfvxslC6fKDPivFcP13lj1ooYvftUjw3tSqnXtJrfjHjSLfif21FUba
c4Vv61KdCXflaNg1zKECS12yKCyvkuOlaO0FYgIQyK9g+bqddoJ4lY/q0seZeiGL
WbsqBs4QaWWskj8ATlHgez+2QoYh3oLTKG9UVJ9naM/f7Jk5uS6xQUG5ngKNUMnV
cUtnR/Mv4iXLxrceuLqsWLPpfgVj8W3DzTlYp7KpzNVKlrOy/G2/r1LG599BRb4S
ChAmVwse2My+J49W6onDTQ8PbzZ/QSWaa0eQ0dZSeUA4McmIT4BzyINOj+sgsinW
d5ppyXk+Z4/C8CJrscUhdqsQvssLjclyPVxWxuZOGi/qCwNBAQjXLHUaBh4nTUtu
xvL/BH/cnJ4EKo+xMS6Jo+fttqzq0+fNwZNUHrbNC1KJwp0ZVIaT1WOMqd4wkgyO
7uOvS0pVeogg9ELdEXRl++D9msPpMU7kEgH0TVKsxOBeYnpbRLB8pFT0Q31VTFR9
FekR7xFx6Wi2l8a1WvkN0BopDufsvPnnuvMrsO/VgEDof+B+v/i2brSqWPSZxkqV
UCvO3/IUX2TB492vmxVPNiGhkuxBvt/8xqj+d8rquHentUuw/OF2ggqEjEPVc7I/
R7miNN3bp1MZO/gkUJKBR0T6j9uEUSvo5X1T/Mx6GUHNlJq01pLULLtEoXNVQgsi
yf46NYg0DRBuybybw+/1Hbprv60NAy+iNm4d8NVgQUtI00FCsuPSkydho6hm9s4M
/SjzBpGCASoZJ2mNZ/McMjWd3pEyke2h4tqrv4/YyTAZDq6m9msoW0RpVx3aiFu0
1DjUW7NeO/7uQBr8IXEMAUNh8o9WZ2qFgxWJpmAAXT7lGaaJgSsuehqDuF1xFPiQ
nMVe6pBuHBewtOx/IYLhdMdRG81uI3oWPByLOG691CZrcm2iHKmg/PiAU3ZhIDj/
THLEP9xZUCTKkxv741mzUP+F4CqgN/GXKlaGXahXCGVJ4iLnaRSYzkcwAM0qt892
sc+kLDE8qJKZrwLZH+fQMbCN50NFJf76VNFLsHks+xb2cfJJjlA9zUh1xjyShSz4
vbI7pS96PKnV/qJ38yVLampz47kGDBool3W98WwLp1QM/wu2WkGKsu6ySUk5bJe9
smNes5xKWi/ZIwF2vGnpYr1rI8BIE9w601fnzk3a4We97ma3FgqQVixX8pSURSVC
1R77pb68k+/K1H1HXurh7MQegP371+pYsRByh2ro+j5uuRhw2Mkqfnh/mD0cU92e
v+1veW0aR4tOK5oRCHdegAwReq1bV5x9mcEy0A7oek6YAmBtWNf3r7SqRcTtu+vu
AKUAqV0+TewNe62mhxoaL3TbQfD4iixucPoHgueRTVuF9SmoiBj5rsGNgX3ZP3lV
h4AeXtetaVXG2qrOwS/S3bfMAVjz34tEODgrsI3x80RIF+XmifauP+BEwtowqt2P
gs5zJlaLs0eZVmM79/mTZ2bATxHoJudHa7zFu2yRfDRJbO4ILADs+NSoIb5Lp2E7
QwGl3azEllgijm3tDvcHzi6bjIOgYLT2cWThKQMNImbWRBLAJw59wkDei4KY9/GT
fSZRN6NwKv7C9sjwOk6uzsb3Cofg8MN1hlLo99z/m/J5FhtDBJcqgnk8JNt7l6jm
HO90nDj4MG7KotCjpbFyuIsJ84g2BeClZDYlE1AT2mHihO3qnp2LxLeFLUW6cq/K
k3khcQDcI9p2pBOf4c0hwNDqCntVFJdJ6T8aG5yBsQJoM9yWOYUS/YljDU3WBsjz
rDK3mIPLURIYrDVxZjgzS7OpZPmEUx7NldDhf3VEA1qkXr8tKtogThxOxp4+GbGv
cK6rHE2hdnumZtWp5F5I3Ndmoz57NCPbaWbp+HxaW2EBKq4+9K1iw5a5i0PiD5OF
H+8g9eI8A2ea3elb2n131NGSnz1LmdeDqF/xoYnc2IZqmupsJEuh2dU20SDvhiCG
/STAjk54oa1w3vFQ16BtYRR/EIFI+LCrFKcjdGp0R7tApIf2hkpjW6mHFNOpyGTE
7TtzZbcSdtqj9HY8A+m5HYYmbEV7Z/iSsa7pjbarfnfBB2tqcVkjQEfIilGopkA1
z4UmQmgc5KhcL8r8YQq3K+2kOBbxzu/jPudN05JxaAvri13GN0s8d+LvE1CJKnXx
3SCtOrpCinXbMrr8fEOy9ciDxE0cIgyhOG9XmAvbEG/83dYTjXPywNNA8GMru1sr
s4QCmIwoFYSiI+r3NfjVj7uCypCojrb0k2kJVwoApURrWD5nO03n4DWbcEFcQpXz
weNacKht1L8PuhDNyFjZc1mtBUTZTzwT9mbLGzEdmDH34JohsAx8ix+iiVBr3aMc
syDuJfUkHm1Y2OmN5qUuKCYgI2hwyLGFVav4Gc9l9/QmtAXUWr3oU2BTxxG+qhye
SSA7GnXHYSycN+sXmv48mkhHNkaw3kakTKzGevFuVwS7cjxuLFtm9yX0uPsWxTha
P12aaQAUrCAc+Da4RiNjRjzlEQXX+jmnLv/RoFzMLTvd+CgVehpp2NEedoKbD/u9
UkkcrpxkRgsxpsjScQ5o9vNErrVzYEesqsrZuk/sBRiqAMPVD7V/SqpF+qWTQnMo
19utNDpMfgLRwm6FOEG9+es/y3b5xBMJgSjaLORNkU0T8VKmOLO7sfY9+23tw5xA
pH+df8ZH+dDrykegNqlz13icpnV/ha43qQHdv93gqEOfpNDGdzcqWJCfxvDbUxi6
oB42wznR3yvtfsYNbbozzGFoJ67F2TgcRag2cHR9sKDJCsC7kC532xbAvHEY5sOp
s/sjQLFg4UWbTWJZW2a/3Bro9+cShS9cbZ8F1hQ9aaEvx3NktK0bAtQL+sxw/yhn
S/jI7Gu9TCP6WsNfxkNUs3Q2Tr1WCW/r0j0Rx1vJ+ZPSQVYqChoi2X6dW4tMpwat
6N2KiIwlqibNDC0OTfrSUkp8c7NVUedYjab5ZByUZzZv3B4WPwHiZI3HIldQBAMh
1muL/P1rFSafd8VGtjOzBSh4rQZ4Ip6jT+DMD2+mAwW/dYNO40LdjTA7JUzMuMOm
3F5V+u1CJtfuhhBcaw4iKtsSpgV86alrVKpDH+28/c1ps3LEl/3c868VSKBgRf8t
Dw5SEopjnwSTfStq9FjUCJV6dtXiYSTBQK05mYwChbm0w1XQWiArlhODZw6oREcW
lhRk/F/h0IxEW4fzAOscQqm8qCkBu2xnE7rArEtP6zs1h35aHOFPAY42ZKnoZFg4
x6cLkPg7RJs/yuXyot+lSK9GB5GvaCRSnDpaEPz0mzUAho8E/9EZd0bfWgGRMznX
NcJoFZx8uCYhzFuW7RMb10T0PVwgDrwyeKRXZKWkwzYZ+oSCAK6lk/rdf4jfE1r/
GutFXBS/HAWd7+o/+/y22+KCCqlTbLM71/TP2OeSt4fHLmgeLPyTTdSvvxNsWtQX
ABoPU9A4+dloGKwHdBV2bcKh5KtgoB5F/r9FGtiJq2SKpmTbqkjGCMe7RTlHf99N
Rbm0u7eTVQDmsOuihpyZ+0fxuzcsfKSD6+zxDgwrDSoI9eSXJeM/oVmRaIAbnl9Q
x0gZWdunfsoLR8a2MRa5w7EuRh8+sLWMcGuKgk/7bXZwgaTORgQ3DdAN6SY15e1n
JPKiFn/s4k7oyjDT87rqBWbVP8lC2BYBd+PjX4k7UvQ9rxARL+fZn2BgCguhlkBb
SAnml62D2GZ+p7d1mApQnhr7zqNfCUM5l8p8YlyY9+pYU+QzRhRriP1r6CYOl3RV
WIVd6P8PCHpkK/7K/BfOk0jpYMhbw8jV1c5aezZFB3fKuht6O1ETM5btTXGGv4Fr
m7mXuOi1oFtszNnhC6SX/M1ZyeL1zk+4aj4l5mypdGdnBvDaY2q9eFg73et+Zr0z
ACQQVgw5O9/M/hVD1is0yyyy1GG4DroSEe5FMZhnapcYnWBuWd8rwNJ08eIy9FWE
w16jMemN4HOqmKr2PFTDP3fRtc0jLDKqmWf3VoyHUzJSWjxYYuHt1wZmd1C/YPOn
w2NHGJ1QYBjr4hZpbp9F0opydfQzishHn0a3O94rxFqH6fMhkC1zMcvt/kDWFcnY
q3DAMOQMbPD6DFrB6pku+myBuSMEm/sSkxDmHOUNsWdJ2Xs4j5uy0UZAVRbiO4PS
AcNpwhbLUq7l9S92dnuUh+jUWokDBkpgPrJuwnRFjLyI27d+4CF4rgjTm5grKJSy
zCinCidSMh1BnJeUfl/bioH4XM1uCOmm7dr/nGfqMKMOYdlgpCmGa8CBggBQJ82o
mvZj1YoM8m1VCLdZPhQkyqD8yPHeHGr6V9Nku7YYDQ/SYeyk6LRbr/ZA331CNc2t
u6NofuQYV4DmmurBREpH1AZMn7e1+Apk/osHU77EHvNJveBBnILyBVWgK9xysOXO
wQa6q2FHaaLt5K4hJmG1X1yTzqkbIAFsHOeg6kISXU/7E0FhusbYcHNHW19r77SG
UmN5D0ruOYRrmb37X2BMncjxKerEvTirx/6hozcxj8bUMlim7KX4dYxYrOXI693k
r8IzZ2DN89q9NnxGQkbzM11cocPWwBl38gFOPeXuHlgjKcqEbxbJuQktmD/FlaI3
kXbMoBpSgj0inSc+fB6QRmrH21UeufWfWiJUVpSkWjkS8DZ2kB8AZOYCIuczjRTY
4FUoIPwy7/MXPL5TYU6rv5U+2LbA3qYUyjRZ9mJQathB0fqsX1eJMDUtAdLMHpXQ
gTw+tDYivtifOPzoZn3eBuGayqJRH5Eg98lHD2mTQXGxtoHLwriUx+q1PcsRkVMx
BJiTe1orRJ3PgK7JyMeR8k2cFjbFY5yk8XYGQ8O5pWF9Sd807FSNNlUim0axJFhC
U6qwGeG40YLFN0TTLyjPYvQVMgZbGsTu0zKykpcGaaOwgyDknYEQpUvVqxGbEg+P
RTtkrVMGRb7YqtSSXgTTjxfzDaqEcsic2GsskZ5yjxx6Po5aXB25SaL5obtBBqwQ
rYIr4KdWeXv8S0NGkel1yCnNq4L0ZA+IiGeTpz5LmE7dML2GgA0mMC70ptpxGdpN
3USftaxXYum4hgbhC17W50K2jbwyKHagm8XUR1OVZtZJ0t6MmNFBhEkU/1TR/qea
WUSfe1KHsSS7hucL6+c0Ld0qOZhx7FNvi1K/IP9+h1bLo3avsNhlWUoYN/AHoKnF
nA5uyuRwx5mpIIYBeWjIU4DUPZ5G4NKkRjBrtX8JoSEiusXBuUyRseBl/0CVy0bd
HE7aB6alHlgzOoqrhp8BL0bIgccHeulxcHwovt9lRzdA14pv0e3pmIB0J8+Vnoj0
Lev6A4gnPazURXi5bnwNuXTIjn4mxxgdSt8OzHEavC7rJ+5MRnvK414ffQNeVSY9
6Zs13y4/7rzGb8jE2vwn7ZPpECbWtMTprIQmv+2Pb+2btq1DoCycc/ckL7ONDQ+Y
NoQQgCEzERnvzDKTU8uJrxVAe2lXZCkY4H7/uw+XzTn726P1oD/1S9QzZCtzgl7a
vrcIHuksytEuVbe87sgPvqReZkWTq8wsp17vL0JSiL2YiFzPl1jzkJLriQlSYTaF
6jHpmK/+mrRuTl86OEAa4qr6NDBmaNJ+Oh7icpN6g7YvNdnzfFkS6o9BT/5KkLvE
GLaSlHFy2dp+GXgaR7HAQ6rMdV4QQCTu8MGio9DxcyiVNZziOqqZKTwuP9Q+VC8O
UqiNhagYuyFaoMBHz1GbGCQRd1gM+MJ3BbeEnU96+G+ABVsZjij5Xqd5iugIb9y+
vd0UWPc1IoE4d2tBzz9s4s0icG+WDU40QR1LNvq4NJdDpJxWLto7VPYXS/4tizGx
05YwqKYuyH1dqIRfdsapydNwYY1/aMCYp8PeVeK4JZUkkFN65RhMv98MAHAE8wN4
kF5vVp5RUefabV7tf+snnruv8otodJEXZR7hTAQUxthPUAfO7cI6D433C3GfDVpj
M2T1qXXOihTjFS5VPCdHiAwY++TlDy+RYbqkLaKjdrB4misJEKRt65vQeulWoYa1
xjH3Ql6jvelb8tBQlZTmbC05zfdODVluGWnPm+c1rkMi6EReUhzi8ia41R7v4snV
Gj/DYkEppeCvurKR8IOjcZRpDTQ5vcpM9mIKKqW9ueY7+nr5TFV6VbrbsOfatm+G
NKpnbz8B9irnZYvBRh4BG8937UGvJChwTB2MqwivFmFpN0JnuqKbbNmGSxiGLfhX
1q3Hf1HEx5VzBfssvURwfY9CNrP8Zq6NN/7SRbsqW/zkGOO13FrV/DrFoRlAmyrb
WjMljaSzLhIqU3qOxCt2WeU47jdzS9OGq0GCohLEi5RGOHv970ANt3yQ6f0y0sG4
pLTL8mZFhNfeYVjb6hAJNcRNzH+TVZrJ1JnysHGwqrlnIlF4KD4HSUNSU6wkzuih
1+GUfHpX4D+bsQ8X+3C5YoxgawkNndBUD8DQFbbWv3y4aviPtGyySUho217OWI9Q
zh75kur9/nxhhx7AcFX+REkfqt73OCqZuseMDUZ9s2dfknR80gxJdvR0TJtFiEAO
JXHWX1JPrvQY3NEz3UVOwIMaCLqfJ30Qv2LddYrOHm6ZXdnUKFoGPI5wZ9u8lxfF
mi3LBLF+W3fjzoySPmyLLayDyVBlN/JyQ8K4BsWp64qm9j6MEJG8P0aHXiZaF9C8
c/AWHO7g2vLHtV0F4nvXPE3ExWYf7UcJjOLE4xRbRL5OxKSfPMbxw9GIiZ3v1StG
SU1WGSQWo3nZrtyZdAKMt2tVoFCkP/uAdS1tQUonmcV9Lc9cLG6FP+lYT1WBzPnr
eJw6p4SzKIMZ1oNyQyKoyJqYSzWekmitgsW0sXJ8pVQkOoP0RaPd4hfcEKCuNETc
kYk3wazewDgbEkxZq3z7DkmTlA0cUaGSdZf/mJmde/txgU3H5975LnEVSH5AxpB3
jUzETVUXxot5wrNNf241W/fFXFLrRUMnSNOuNpJVgSRwJg85T8uAJZn9kL2hvzE0
gxnqoqMW/9TnGx/zYSWTIedt5CEGrXQK3k1tHyE46eYliyagqATF3QmdyY+KLMlq
0g109JqMsDjWpKy9GjbA8ne8wIoy95JkXKBKKJeJaGLgV2DxeEGW4Tie1e4lCLf/
P0uvk1lOTQ6oCZfbV4t/pW1J7XX+LrOVqW03NnmFPRa9Yv0rIVVvFM+T8L6SVdrN
eM/6i9LtbppF1dTOZNkP4Bwnr1Wis1se8Nb6aNS8anN5ewBbh2NGoZNBm5VTZT/h
JfSMGBBtFobx7geO2/AUYVMCXG0HlAPWIdIAkVodZzeHlRLiJMec5P1JiCcwwNoW
IXQxZcktMDfvHXCog9BGxXXOkDHW2JXSuxLXw3nKTbgwtwnyCh0rc+v2wUnuFlGd
8gh4tMM/XPhz2rfv5gQu1iwX9DSlBbVt+9Z2ay+BTqdtuenKdqh/aWJOt7SvIhob
mSSpBILQUDOlN8b0UwEVsv0tSUIOy23mYfK/t6IxtOg0JMC7UBp3vIQwOWbPQRPK
+Xa6WqyNAhBWQ/Cb2zifiYaudR6qpdKRqPNNXuDXkLcM/4vqHhxW5XZ5rtbEsZNA
mo4hYixal6BGlgygf5bcqolDvFhS7sQkiNmLFWMuHfHkUigWQ+TyWjFhDQj8hUly
FmmHwwVmjfZSquq0NnTv1jg60qzyOtH7PXVQ7h6HGM30JXmfitdfPgiW4maLQvGu
JSg2x5bQJMLtFKMn88ZdpMNYQQ9jpqd0v718mYVSXJnGfyf6fQ8oCuEbLoVaxGz/
1ZDbSJyc0s2+HhVo0XRKjWL5gmIax1mKkNHT/Y2/h4N3lgRiHQLsN0SgT2pN2TKv
6PcbPKpHzndfBxYvwx+8AzSCcb3c6LQDFnfhUwg7xD/faekP1TairE4KcLLW+2fi
z2aFmN3ZXdB1THM+xeEl2vVUXw+tBGLTFvIstwaY+pNja2aBx5Pi1x5twl1VYwIN
TWAKYtTuf/g7dyZveS/aMKflDIz1iKWPqKGEP7eV5O+q/uXXGzbouhCpLfzOI4Cb
SdNVen4SXE8XcsVgafaG6ZieDzV+rMv2EGDrhznxT4qY2IcpcmR6P1E2FDOkBM8i
ZsipDVulwJPUCSb9Dk6N08NkJ9iMVLZqHp7f5Yx6rrUkRQTJzUJC5DZoFQHSyWLm
APmBsOvjhEI8QE7dCHpfL859cdYqGieahenN6FTMz+DF8wrri6GpiLBnF/wFIg92
8fVrWzpj3cAcbpKLsXvxiCrZ4ZlZHGWEQKxQ/HvjWWNAkDUzgQu7uuSUyRJZ+z9c
DuOditYdi9T3dpAciK4qWjTBSfiUTDaLNuL7xBPPqsJGa4sI5VKF9tWD1uRQlhtx
W5oLszDp5nVIlIAOycW472NNuWNbrvpw49NdV0hfXZEHKCNGIYqxMGNJJB/MLgH9
gQD65ybeLXNEvEMMKk9szLJ75fRUUhdYrMvTufUkZzr5S8kiWQ2sQwLpKnbpxoP0
iaZkKOw3LSsKw+uApuXUMiJyBAjfS+bN73eDqvOcqW1Ade9dhO20PiERKLxEovHm
EVssYAzjxju4uF4bU455oFvAb7B2TsHEnCTN+Vwi3DMjFVJUHrr6loLiQ7JdLfCv
RrFD1ExmJINGpQHpc0bUk808JOqNcOAXWsr1vlw1Z3JFAXLV4kSosJ317I5Q18j7
otI6JIcX1iRn8snvDg8FghjnJJHuEgV+DVLCC29YPlYl4vMjPCxtdQAYU9BTqhzb
OrdwYV23GeoxBJs5NFqOrpp6Qi/8u1f/IPEGDpgCYyeXSNdg7aWS8/lG2xFAS99N
6eIgl/pm5oFe+7qE5nV2ggQc2N5rqJa/4A7K4fFO9qTFtUggY0n3FZwZ/r4YgToj
csZ8tyNcBBQx9d99HBFJuBDl6WIstWc60KmHBYrf8bQG/MyTKxuhu2GamZWuzlpr
Eo5PVHr9H9fLcW/FP32SYT0SqZ/f2UX8D5UtQPqguROcAr6/bvO6AtK+klSOvTRv
JlNH517lzqACyDojiZ+oaS48hVRLUAQ5FGmoshKoVNjY7ylUVj77DCI0PN0Pf1Er
o+wKVyhiyPhHjDVKKQgn7G0tmTu1HxNWRKONVCb5AruUudrEsVyF3Z/M4gpBT7hq
H0/1+m+b+NZd+Y9AsQ0WzbmGD/PqqIoBk12LZelPiWTtLSk11TnAyCCfmOHoj/ER
GrpkowVT/IXQXN/xYBsVdj7+DgKFNOJs1/AjjRAgL8xF1xgPiAwTTcsTtMdc0FS3
khTIz1CPsqwLupw0SRSblH6SGyV/MHVkRNxqtyH+I+wESC4/1OvPLZa/VYq33rUi
uRhFy72jgkCWcDyfjysfDEYQ/2dqgvPM3w2RwMPK3Cbh0+74pgeqhJ03kNGwMD0m
nvyK45cnl+rUEowFDOkCEKysnGBsnYWFmLAkdozKzjzqc2hh8S5Ox/W9P81qxXsh
JmVmI7BK3CZ2B2ge5A6XQjKZzAIp9wPvx0BNaoLbWNSD2hSsT2lyhm1tFCiS87mV
kbMA0uz5xeCpimyWXGt7M/f5PXMRypvy2SWZpIS7sDpNKrCEf+A/xA6vNQ6fSozb
WCRQQrGFW+LYv2rRyikrbiIRaB1hW7qGUvdAapEbKqv6LvbBLduIh7+UyLgn5BR+
opTWG9EEpplIe30gqO9bKodXBum3N9CFQ7O9pYwPh4aVHBY0KeGK8lWMNAK8u6LI
3jt4H5S3Wo0VvoGMzF03vvogBgu/udp3FYHsqDWfERAG2tAlRmK7OpGZcW61nOPt
wF2h3+jMDUGBwL1pGc5kGbIRfnxdX2VxohrVNNCaxmV8RSYj4ZhEutKnN4zyn4tA
jSUysp2O0+TMF+BmmMuO4F7uISGIwUCTJIRTg1F9na5eUPqtLzvfFCKMcXOhjrzi
PJuQM/1/kAUUMSfXNb88ZMd7tTLpFB3EfGdMtHWlJneX4m66Pxn/aLyWN8keqjlT
/2OdxDJbdCCt3MG/6PPUqUOgB1Zfe5P98nKMplw3SQ/DENVp4aGwUTBet+KF01Ot
LalrNJfdJkfMHBhaclsj5IwhG+w38dxIz4sEmmVhmdDdpki0LFVdfsDV72Vzjq9J
UUTRc0fOG3bCyjRZzxLOZZNXlag6o2OOeGpFZoPnb/7tsSoSpUglpP8bpWT7f3g+
LSvL6tt2O5lgceopVKZvAf+6n8qtFLCIDBzMediyBDkiJeRXkcqehj98xalYZ3r/
QXfEQ+0ACVi8MRjG7aw3aqonXs75FhzQgVzHidwFwDiF3C39UhoB7C/ePAbTmXBL
XL8y1HeE67Vf+HVQ2nMbtl/Nlvn7RwnuwRT+aOYZxY7SddobfXVJ4nvUUkD3ftyP
ojA6hCq0igLXPJzQXlGEiGF5uopnmK5sujCWEmyKJp6rL8GplRviTJ++oFAgdV6u
7R5CsugX0O+Y/uivIRinqGRnyVoZDPayi5mlN5T5Xd5wERblXXLwQzIe1fjIERlv
rRGHorCqM/wFGYGdod4nabsMCJntm6d9OZaGVDuvf9VcwjW3K8q7iT7fzAYY+I+p
sAwqnGeYmTZomGgD33tyye4cBVDp7KxxFBT1xvBFa9AmegM3MTsjHmS/kRK2eDNQ
28V/XDFJ1g1vsi60KMG0BN+CRxSF2hYNp5qfGOEjGfgqtl1DtOJCRerizYsYJASe
9IhwegQCC9OCzAvoWewC6cL1nhJtXvtxuyFhtdGCP8JjW49xDGQLmdcY2ffG/U/9
FXCaNU0w0nqwRSMqjha79H0LLMCrpTyWyy4xvxw+VhMQPFIApQQtwC+rCR8wle01
xo3j1Wus6YPnrLiwgCkLQuElWikDnwsseNIo+VcODnA/OdeNGvCQSr/If+HRTjPV
RHSjBbC/FEPeN+45fEotIxeMzAJNThFjxTIrAsYBPrQSK+QbOFUhL1qrl+JSMgAK
gw6ZiWv+U4TRkA6hjxo72CJmxD0hAVGrZO/QUloks1+4yks+7rvG7cJmMOfPTIU4
hfd27jIT+Tp0Sz07nJ7C42MFNxattbLbNmOLnqQtv4t19OtA+9gDeoc0XftGwLns
86D9jd2DyUjcH0yPPdVLAAX+fUHqgYWBFBzKua6LRqtYPbOqZIz9ODxTUmuv1TgJ
QzjYbzbhUe4/ikClyhC834K4yGfaKJ1maFBHQFHVtJs4rCgU1JkWHLJ3K5AcZsNt
Congfy0QexFSWXwRDLHk1IMeHPjacDSkE4SkXdvwO4P0E5M7isjtKrp5LEbscmWx
+4+yt0zKGrg80XVAPkoWhXC4k29LBQOIDG/b/9ruQn0TFKBXxVmWyEotGx3xtJE8
fPcWaFLIro9a5TwgWslEUDNEJ7V5Q5XT6LEMp+gF4XR7P16xIHbIO6TVrxyWJpzh
x6K0Bgqf9/kpWQrLmZbcQrcahjyWU2YNao+Z134QIyLIPZ8vYQMqjK0hAlufRdT3
7GBzizLZkMXm4HMyAZR8TWvSAdKRKf9tG9N6wMxrULqsXIzRuzyKpxkSIaQp+/gq
73NA3UZjgCiR4txAUX02IDS4ogJH7jsanaWlLnX7YaVqoq3/zShree4LwQag/0Jz
g1YFigIyv78IkeIzFUdumab752ar5vFpyU91Mpi6Xef+BiE+XyXQ0euB5g/6KBXX
HH7Re3O1/rGNXtGMurPSOIJmfeyos9jUeX/FUI089HXCf6cDZu8BgKH3msuv+uxk
XfMYcBIiKidWCje/rVmLFqqiUQ3zyj2DY6qIa9YBEXElOi+0ktIk04lIzJuxF+4n
2NEcWyOdjzOn3kzlrMcN6SU3LuIlAZlN0IZb1wHAEpmabowxIL70dELy25dV3Kdp
yaQxwQg5Lilq8AcQovulDInHTrfCwRnR2etXo5bExp3QkMIPu2kKYydoVlQ/dveu
Kz/GgMRcUmFyhS1pj0U0x6KVryCTuZNXMPIoPViyBA5w7clujQ7txndu92ksQEu2
NHL8xzORzAQfEQn/U/N7rPPdAhEA9hNxs/G03S9m+oXuxcYVUFRMP4vqN4KKVffc
nwoRzkq/hrpe18XPLmHGqa3HNYJw+w6dQcst3FE/3IM/wzzpJZ4isYkzwBd9ytxs
cqBX831ZMhI6p1bX2oFuEkKXZlPaKzPcDeL4YcDOmraKErHWV1wuVhpgYdLCeRlm
G94sNixXc3cEOY3XjA3BuJDoa0zx/n/1DkjR2RLfTpFMiJK64iJ0+cUEhHQ06x0P
8VR5hqXSxPZzVrchw3sRURFXtxMGpXWSqLyn4FyqVw2dXxlAjeVRXbpIxEcrYNMN
jmbwvP5hyE/EuAUXupEWMbGpRxi3NgIcZlPVSTe+7KJwcbt+acbwwOMr09sDbm6a
5XEPEFDnPTwGAXSHBSbbzSmUv9pgnUtj4awQVYEIpMnXca56Hb24uJtZZupIfAYV
dE2n3uDrlOHUJJsaGe6mSvC/HJ736/eg738pk1o/6V5FFfJMqeO+1NZ1ORUuDFc+
55DbsH3gr7jbEKJY5cOMpGFUF06nbC+GtNyU8aiHPWDAmfIcooBI95UbI0OzQfKv
9uFrBEiu83zr2WVV08e8M1WAqJrZkCgunJm9t/0vyJ6LRAYWjQ/Gj3MgFO8QZU1+
RK3E9oExs6Oo8LHugtmAMrKNxsA9lMEFO+Yrt6HtnENmcgZHmT1tK3tQh4moxnuW
Tsj6UgWnsI0t2QADxoGr0o+RilN1rujoWiIB+AqwkhxrYDDWGYs65cwKSMOYqnSF
pK14D3PyROGR4qSpDxCq3TloFx8lWkhLtBoGr+zJaDaXRT6fYS8u4RbtNQF2l+6z
8RLGPmI+t18ec5uOgBXAiD5rbgmzUq0S0TRALS3kAI+zHEaZArZywzA1PtynR/5P
hR+4xHW/h4lq7p8wXY7qA1XRwfbWIJ8kfr9SL3PIpANiZPVTzhvspkz+KacyPHhR
O6mCZD4suMnMUOA55kzmT1yGiXgbM4/elF3IpaCM4wwMEeRD1WuiJCKiQBc8v4w2
nG4LnH7PMNCdce73ofThNsCeV4NT+r6dO38cc28aSu6OOUNPlWAdoA8sBb7wHTYi
So4bm2ge5obd3JYpGH908As/78Ktr+WKn1QOIz8KZFvylE/St5oQsG9wQsBLe4r3
cC65oDYH3n7Vud8DP3XTncGD/1U3d326hEZ8uHSw2Y+5ixGd8ANtzfAw6tVIAMPf
4jZvf8snLdTO4SnuD0yr9XPil6VEvD0b4q3trlRHbILuOj/WXRZ2GOmAcyk9Qwcp
pUbG0nBMkm5dkxAyYPLldqVhF+9xVWBG3H4PxUxeEW/FacdCtkY3EtdWovvnIiKz
hIJJYfHHzlW+C7PkXR2CDL0KerhM/gFA6pYtx4hRCtK6Ujr89indka3BkxJ93nVC
qkVx0IRgEbjjWmEpSlHvrZ3OCgGUTyqXTzhqJXvH9MFBbOIdg1FeT7bNmWKEuLUD
XYhDnb6n0jatm/dpC+WDEmOFPJa6i7a7CbZN92RxqdK0/+B8fuQQC2TsZ0xr4stE
c6kylzz8qOfeXn9lxyAlsKg5wV7ZhuQAzpugwoKe6Nh9myJbrJid9zzz5jbIKWEM
ck09IBvyIxnz5iJk18YTPyslIH5JVzH1ByCelfVDN5LouotFAIB7SuAbDxk+h27G
008eMl8khDCVAco8z72pOx+RVX41ziTxudtXsx5jM/Skoc88E2pUHZbn37zeOmkm
0p6ldWkQXJh+CIdejvQKSP2gZ4civCbOEmAjNLzaGW1aY/9UCJkXL4ZvwjWc23gR
p19e8BflOGPND8Fiiy16fsW4DrhIT3qxvYv3W9+N1EJC29G8CXGTfW6hGttXYye2
6sYtTYMkGR72S4sZv3G88QNdmJPLOazLD2YITdIAtsIavkZVLL2K6TVL3SzJUobR
DeegyQG/3wU4+oJ9EtsDxEYwqd/A0WOtyBy2i9Ev5fzM/10xMQdIjO/rz1uVyH4o
89mM0h896Om6P6JRo07vXSo8nVEUCmt0fkk263kj8k4sd2C1HEThokrSrmazeDUj
cHHjBlw5CG+nJWahee4FMd0ltNPNBQWJMgnJT/6nnOgPh/HKraRgKJFNw9apn64V
2CCAMMtPoGwFfTvsC7VKiTjWG2BTr5EOEq/KSGXXHTssg7LldwKk0m8/zXFj3Qvn
RrKlLgBlrzVXATQa//P/le2k8mQvg/wpjxgChV0GOfmADdT63p8hGoDk4sUIpxRF
NotVk/SgReptG5gqeLic2mu8HVk+Ju+RCGwoeE3V1aDeY6klKPniovF5e4uiradn
ZwWNT1GXBdJ7KHFEo0yexG7m9rdatcrh8hxvtkQeRLMrE6QoHVdOQgPYOihrom1D
l9H7C3wKMjQNnvesinz0NKaffq27VyWnYZpn2FPXw5SJ55+toehbgl4XXf9Lik4s
uuSD0wXbyQYMWcCAqqzEMm+nmEbtDreU9QnR59m2xKQ4ySd5AT0twaEn785aJXcJ
p0vdmMDaVyA9Wh5d7AvqJxi8vLnQbetyrOaZDBZn3VR4MohuBSgZ4MSHOe3OHpXZ
YSt9ZRSHx78hcJ1HhsraoXuBo+em0H9TbfRFSJ+2jNxCxMly/OOA1l7s5MImhMVg
ZBmfJuyoRq8cRxYBnBo0xXhXKvPEJjXwoXEbnOYvQ4Wh4tx33RHqNCCa3muIxVek
oSClRGa+sMhSwFJLcJN02+9Pq7aqtCqvkJm+OnJLuQJ0RHmDGnhjgS36EwG6/Do9
ndzmBMjZKHnmiKmIO83Jjc7ql8tahtL3lnaCe3Y2VvVfWzCIY5biHSBDTPom1Tbo
W3LBqc5NP3QFmbssUy9uXz7xTakEmO9yYkMmcJ+5Ev4g3mpevsbOC6BTXgP42PsV
LXMT23pVzd03rJAcv9JR0qfpBgacWtFNIClIZrjfJizIr9+VuEznwEMd6mY1mFsj
M8Npd92B/KheIumLlCXpaMwuyl79qEW8+8oAXPZtWeTAdljoyzzZjvG89/1DqyUr
vn8R9FZZSVaETsBp3Vu0BLkdvTBSGC9jU1wCkFr2yqXO7+0YMmXBZ2AhIMTgEYgz
hDZ4NbC1sIzAKWzd1fL7VU1sXr7kN74DzrvI3Yv2QLyDZ0mtYSKF/Gssn4h1SY9V
bmmtflbRjWRcTXrjOZl9kD+bj84lvw2AwRoZJta8ZN463qVJtklkJ1CdRJa5kb5B
w0NfHS1j5Yucz2dumvwMLzaoMLkitkYfvlZdIirbTJ8bcUktW9ETbT8NfNMP8Yf8
Oe21r7iL4Hg3uIS1E6PabevsrfWgk4dxgRY78rnEPccMHHQ7uNe7+CuqAyuHXGga
5mPmaTXN6CTCWJz4IqOMFn1LALaEQHMYSMBI0UztKGB0OOAPBcPy5aF8VqemtqAY
mBzyOwjjkPb/9UVsTL1HiAONNC+BckVSlGcBSbvN10G8+iR2GEzn6GsPsMJUT9YS
wLmG5JN5r3o75Iv6a7d08W5h1GPTZ1Jj/Bx1FYPWDJVNV1o+S56BjMo0Esqhy5b+
02NHwXwY3W8ZwUgfyoTE6JbnWkSXb1P8T06i2Sc+S/NtGVk8Wd1Sivos2OIRI4L9
b16ffhqAa+rVSHjbKfcqdjNX44vqKAvapfhRcnxZYpkRs36+Ev1nNRKwwQcH376f
YX2RqNMM97w5e5DAXdJjC8RYvAk24XCHtmPjYnE4IvFvuH+65VJaCHUYd6wwMUmR
jvNvjPabumtW0VI76ge1i5BcSRWPJOFtuTr+Z2fWwVuqA3nGikixThStOF2hH63c
iZhjTpkqKL86QpCaaDiv6qjVtTRSDisLO42SMNXfYc9xf519xnFO16DUi15+Pxcu
1WrUGETFty+AjOQcVHPkECusq2txwPx1vEiLco1Ep/oJWzPuX4Oi4RUixPXk3/fc
E79QjuHZvjQ5k7053Y5rRmhA3JKqyc+U9LaeV6j9V51PrphtejFMGA7K3RiSZNUU
ZkA5xwz9dgugP6/exLOJF1PKomwhUSvZS8JgdeWQPLic/+KzUGOtXKmO24Z7Pjso
PWXqRFyI7EglP1P8MtLhxPLbgJgecU9eln2aP0t4r3TXAJpGNpxS6p5oXMEgAp2K
3pRmNBMmcFGRzXVhNoBSmPFyhPprh7yXig02ulDMwYF0IOKzcZR1C35ZqrYObFbs
pa1KFTZ3sA1H/G84P/q6knbbyI1hnl3I2gk4NQ4LFKnTkUDb90/OCpySbCcMyxFC
gZk/EGsmpUF37iROosfHADzxXe+QNMT+EKPUg9+F9bG4H2MUZ8mZaZfxoNmZhFJ1
EYhrlu131Xc3ig29mb6eAY7qEcpWa8SVP6frvVdMTtZzS+E34DcAbeGlyxfBoMhW
yYuTL1nEySgZCdinNQGFi5Elo2bJzfI7f8oiYYgMfkWaC7zCdoR7mjAls9Sw6ywQ
MdS5H2sJC74evJmgXvMOMs+FyzHJoATjCAkJ+NS7PG8rIWUe4Ng0VRR4C06stmyK
xJLk0tPzUA048irDVviWYPN91Ma54LZH+UklFkbI2/fYb7KM0VD2simSy8XGa+6B
pff5TfW5SyINXj6hIHNsur2T2j1ydmTWgKQxMCYXXQwWBhbNzvEGOIam3lmCl2QC
3IjQJY91H0LY7gUR04+Vphp7KUfubjSZMShFA8jRGbTTDKwWCyoHTZgNRCLaigyG
ZddHKJtS3/SSHEbM4141j7DA3j0/SsTFFUNeQ6rr4K2EH0mJmQxzz2xAhO24mP2D
dbNz8007saO0QuWNsstnUqbH4YSv8WV5/Pf0mD8vr2k/4Goo2OmtcsOqB/Il1I1/
Cd4zCTCgJvY/BoRE5Wpn26aWoEBZee96OTZ6aVrOXrK5+ZsdiltNxtlXb9FwI99w
ssvsYJU/cFxo9mjuKObH+/K9wRZ5dpdaoI4SiTqM31AS32P1mFYerC1Y3K3S2UXA
58Y5+wLZfUmiBxP0WF3dsE6YZinUwb4JviEvq98RhXMeklMI8wX9LpuYOgd5zgEJ
7iUiL8drqt0lj710Knn+SsbpjP1vBPa+qxXWbHYFptT7YTXW8WrLLySn92i7QJcE
ivoG9OSe51uE/89gVc/Idqabwf3P6IIyPpURfSV4aRV/b82s6qp5BXVrtBWoTCvr
iPyyrO4I8q91xSP0l2TvWz61C0NEEAfMNer89Plas2Zkf9/0CVk0SO9u9tJOl37f
c4ihtXTrLcvbSycAz6oXxxFsoVl/UMeM0krrFiVcI2Lo+QVPhCtGVQIx0c/3ellB
VvVJDpPMDQDzxvHtFNjLrnKpllF6Y4O5RL+IVhkyECt9KA7Fervhxep4fXq2uAv6
5hPhf8F0e83eJvtcp0lgI+5wcDA0MymrC0+bAAuTP4uMONUiNggMsbSb1sXucTfJ
vNp58vTbquGNbKVMA2LnzHLSC0+lncdOpPvBw/r5n8Ilqu+mnQyN+KSI0dT4yL/c
FsyW1Lke76aiNzd6Ajp5fAMmfXaURnfk3ftJJnJJ8Qihrkq+J3cPwDQL/IQc+NvL
Q7DR/eszMUmMzifpSO/e2VJJYOn4WXHRLzB2CTxMIdcTcwlds+tDIN/nmc+x0WNe
3VZG8aW658pD28v9xZh6/EgBYcXj+WcRZ+UhOEzSgxSf+L3gFaRYikGqG+y2tsba
5Dx8eCe/DUR9wMgTFeP35Rz/uApID4TnQzZg2wqjoBz+dWl0bxw+jA3aKLCuLZvN
oNBXMVzLfLodIr9fY/w6hG/cli1qmlFHW0wkolsUKG7IbEI2jfy0cDnjBAJN7zUP
z7K5LyeIVU0w1umRWPncPU1EDRw0R0zolPuBMw2neizFPY2ETPkovsrrC+MaI1dN
seaZvH/R83d2TPbOSjFHNNJz6XyU0LS3EUyLXZr98NHnMrXaAGRuRnBakeNL1a55
x+0Owq3fqYTyld1P3LPdquR8klNR43aOOpMoecdQkFnZRpAHxJa0oROPeHJtxvM0
NK7Jh8x38n3mhE7fUKQQ2PingDnOPYTTlPFCwry9mZ54OWoLYC0GzdOxIJejw0ub
4eiwff3HekCWt3XsjWDVgqYKvBP0s1Ak82NbGWDt3y+ITA6SO+E5bbGzUGNYgw2A
RtgQIIxK3rqtzJDjzxuYm8i8zy8M06xngmoRZ2AW54L8dJfD4JocqjSYazMF9Naj
oB3OKodGALFlxExqGa4Z/IA9P6yjNsUdwy6U5f3KCY+rJTYNk6iRCQxICJ2TS0qz
JEiX5QrSY7yeFEM24t8INln9LOLNNUBJinMQywMoqmcbWRkCvxLVkdP3Y8/Ozwi8
LzrI4caDxOPFQZH4qy/pkEO+WEYw3uPZ1o0d4Mq/em3s9b9Yhol7OiTMbv1S8szQ
UrTsCJFi+Hl2A382POFF7L8gL9gQ/wQi+H3lWeQauZlPFmBCWJLeVa6jY0g5nkPw
1B9rQqeeLZq4LAFhnMF2eHGL30a6QFjVoS2wmspHNTTnlvCS1M8/Fd7171v3eUsF
O1nHqNewDdieScTRWmojQwN3szeHlBZaTG142DtBexhEkw8h63t/qqclTn/IxxO6
tlUz19lsJA6kpBLaaY9yonIxS89eDgU1FO8T5AAzHJ34bcffYYSesBpf8UDgFlgS
7d7tdSUOo6fGmyVHGjeV8k2ZTwZqWPjlmXF18sa9Qf1gzlMQNK3P8Ji8+DPttfJ3
A6S2mvmvLaP8fwauu455s/4xLmah57PMBdeaz7wfT5QrPmiEt+PCDC81BemXV1Va
f4jUm4bYJhdpHLnpmKwOlucGQUTfLgba4O8GiCvSZAoV3RI9++2O4U9bAVPBKihg
E0zehtdyXo7HfXoN6mHFV+ywGHimOw4WtosvMaG+lMDypaPttB4rGVBweraxLO7N
6F6i9rKUYDg1GjWqBER63FYdfS/nKOSDLxCrCLZm+5zgGbDJbf+WmJyuARiWGEAD
igMQwWY3t9IGX9E1JiFPNAcsWhiQEweocfFCFKyxOHpiZOStK7cSnDicAGD3wLyu
xCowKh+oLvCsC1q1z3iW79+f60D8DON+aDKpAmL7wIsjSZ7gxYBpwFEUcPxIxi1K
dd3+ORqKDww5PxfBRH/AtQLJdXYXSjX5CxJFwCW4jr4240OxAgBfdrvnWMZMFdK5
c0LWmlXk58alXhI1BbxrwqjsKVLjiJ4xrv2AyJJZ4/404+HnNwF+ICXzJ/iH/Flr
k+ZeloBMlCUABds8Vn7Y0Rt7ynivSnzRuDNGLn98+qNi9TjTCPa1WHUJPjxF5o1y
4dAFZoNuaOu51x0nCEYoTK9M61J3YzlrZlnDOOEjfDI9K/WPLkpp71IwpbYQrRlO
jmtKK72PSpWFGgZTSdDE/w0LTN9vJGbHXE5D1mhixCUWSohO2bL9GenjMpTIYhLA
x077uUMJvLjKf8qezXs6+AmLs86uNF1KkMWuhRziKafjAD+cH+UcG1bz27A4P7+P
tymaHJa2kX0uT8Dyx9FiuhHqXlnednISOuHIZTws+WLyxsx9pDbbv1RUnD90CH4L
YqgkDNvNZYWKgbnGA+3AkO+ne3n6WrUxelnibfrNx/zjU5ayoGtuamECohfUGagZ
gnmdG2emhnoyalJkLJGy+gQV6t7bCZ7vPsIVQAfiiphjJIvDs2SO229AMgjmyx/Z
SUFwMn/f1zcNETebTvY8r+lubd8n17jEyiUCMyXoyyKbrEf2sJNTNfNpy3SDqvfo
jgM7O+8T+jyUWK6QOmcI0f/1rQdwsXXikn/jaEDV6OmevSUpCwV7Lms0lLWtLPg9
II18U3+aLihZYp7ZWYsAw0sSQlEM6WO7BdvLi4ya6eZIKqe8aSKgsxN7glly0Pur
xZeAxT5toMvBdmDMRQ56Vy5rP9doFMTmTFlMWeMbr3gC0QW/RNBMzf7aFlY2WYKC
dh9lJsDcOXkgvPmcnct64VW2tkqgcz2K0voPVi8QkUAKXZY4qLcskX+tCcsFBDme
L2UZWzed/AZR0BQbvrDA5igLQuB5GECkRTdpsBzz6wDOJXD49K3xkyB7LA+k/nXg
QibCskWyymkep9YJWble87E1KjKCXtKAJstGvyJuJvHVFFv/uz6L3o7cwqTdjAAM
whf5pGpaFeKLiFfJco5/hsjur8Afxmt2oJ7tTK0Zkqu9pq1uWXHzPg3uxpvNHaCY
nn4zsWqAJ2OPzjEWIPF6jVXShJWyBuczCiqOVo3B3EkRM2xTx4uAMVjziipP5uRh
9wzJmjpEd3KToLSj6qe4z+zIIw13RDVqvvFn85yw5evloUh5eAm18+hUlI1ay0oA
G6+wK5PH9zKEmRKzxG2/vZMLsQVOO6yRTCBr3i2L2QHLF06MSJl9wMk04mdRAE7i
+hOyRcymu6pOKVZ0lg1sWHMiZbdx8sekAMp0FJVdPFB3MDN84R9b0r9DItRzg8gU
h7w2ruK/JiD5Cw+TIW3GCcqsk/WgesnYxogWbMGdqVkfZTAbrmx4JcOl8cOV0Wpk
e+BZLKhO0AtV3IRMKeboI6FR2Um7rgCcyAwsAfCqX5oh2o/aZJYK9yWySe+y22ow
9d5QlG2Kjy1R3GiANLP8iMUh2clHx9ICEDTN1u8fV6drfZA8HFxZLsah3etgxJWp
v8KqxbfEzkClWKuEVCEF6ZhAcYok0uBN3sQLZ6TqwVQvl9jt6s51D1fIYhhxBY5O
2emKd4BqzrO5HinmqsQedjewkk9kPdz8hXG0BRRV7dNvHY47Il7MJY1Jrn5dflTa
pKjhcVxy/PThplcr8cuM585AlbQBvO3tf48v9NuNY6fqEnzJfQoromI1yb/lBs30
yvXFvmeY8rhUWjjiTJU9McwC2eBq37vvR8KSHs8Q4HiJIPJc8XIWY2Vo3YGEtUgX
ArmSlS3wtoCSVOz5FNf2gJC4kYIJmMx7htyt6LXz8Wja7s2zCqNbQh1kGBSimQ0/
Pv6M5j2zCRf0bq9zYRBhZ/3QwkXH7EqLnFrqDbFCencuuYBEJABp8CkXAM79+DKY
+DHCTENhSrzoH3oRZJywaJM/y9GjeW0iIo2/sk28jGNwE/hcJ+gjtXRUwrEOHrJV
7GFBDEJP9zQDNZK8brS8Ln9WnU3tLWiylWV72+VOW5U6PoQSOcB29LvgIJi7Xgvs
tLO4qgrL6MYWejeSA+MRKfZghrIYR3FZSgHtX24LUHvMwG2NZWZYDYlLq+3wOEg5
+YFdwRseTHtMAZ6zVu8ONdtHzIxY2R8Jmgu+0jYKVfqY1pGAi7vqs/j4vdcVyvsl
n6lTwMfVsS125e4Lv0eDF1/QfA0OP7bMK1XME20hIX6Ltx+CboJ9876WU1FdKs7V
Wz+jNPXJqqByK+2ftYy/0xvkxvFEdCCbZy5SqTN65sTW2TuiXauJFhNH9BujNYJx
9gmHCJa5uBX7wroBOq+uleKen8ZBAWWNr8Hceti3RAdzY43Cg2xSb//KCZkiadWG
QRfeYbfm9x80QRXKokrvbpdaNCGV+uS7a6TLs33PaQHDWn2M77KIMWPBxQvCSodV
VmyIR3ROCYMrKe9Ei0uujnbHXei+GTp7GXty4/EztXOVeCNjJFmiPEQb9BoEHr0t
DuOwqasmztnUfIXi8/wjsV1BoSQYXdCGjuviXehWyFVtYxBNqtq9npfVJ43OL3Fs
qPdbpszftr7mU3Dk1QhLFVI1EDf2VurqWRaA1Z2zZM/EO4yL6EcLS22YeOiVdBxz
mJsY96qtQudjbneyXBBVYZ5bZSao8kcAXqiCv4ooEVrm+/6LMTFYIxGluWyP4h43
RrlK3A+9hxV6HntG9nOJPWF1ZS7dJyUK2v6faSQ5NVcX5kBj0ymap0FvRkecVk2f
EBuWVUe8eu92ZyDIL7+5xRvjTIHGK3Bv1jJUUhRQlYomKXuB8zzzK11kzNmsG7zq
wCC+YnIfOS1E7Zhf9f9oC+xeSIYMe/PPj3fZtoEF0IwwxzqRPzApAvnKttLd6SpO
ik7ejRa1ygS/1ETiqhjch6aNuLDNaiughQwvdDWO5RhkgUBvJkl2vVGzNVekghTg
jFGtaFu5xJdC7bjzHzi6ok4JkLBwYT/GdamIeM7AfHAKurRERpS79sIfQOsynUnZ
LFLVdtt/74uBLQ7rtzWWoZyuJ66siWPTpLARQpadqsGOm7reA+QWCSFCJX3u6IJU
IQ55T73RFxtRRGXj/Al9/PWSXXZ17AAicRYPSVSPKz59swyuZY2Yr4Sq2mJ6NLAV
NrPawKfRyCrkpApCDCFPIERxKcP6TKJ5mdudn4cNNBx1uv9bIRsT8wjMhL3CInyT
AGU2FDJbUsErWu1FXRcxbs3PvqojS1KAt0FujJWbomTQNNuZMN8McgAgNGABmSkC
LIwVmuHWiL7yrP0HUApwJM2F4DcH/6J2GOP8bxzc8a3H3B3+4MFJHrsFvWLEYGQT
nH2czHXW54W7oIHWdzQ2M4DRIeSztxFTku0jnqwh7gryAKsAkmpqXG5sbXU8pAyZ
VqAhS75qb9l6Llfq5Bg8Y26lgPMFHAiAlijp6Wqk0vvMTA1WVoXF4y3eqDZTm2WG
8D7lokv8KPeMtnRN5yLNNEfGkO/32iQmfG3RyM73cyLS0XO8M2LUT0JlsC1UyO2C
mkm4WP3RVQ3ZlZ6/tp+9n9I1JUFo3+WBcXhKoaasT/KA/3CnYxleHlG5pVb7s7KF
+sixu2K9RUFAu6i95VwGi/FDzqsoDBC1knsg5Erfk1jnHShL/rACYJ7+U+/SFcbB
/gYXNIQsZCK8siQLt02/ZLD2XAT2/R0L+naUFUDJWMmMmD9wwk7kQQ/2CfRxTBA/
6wCKBw85Lk8UC9y8GIbQXViadsxCXapSvel4YMvAjwbKJNVdp+78BpVILlZm28/n
uOF3aCD8CxAmvu6JYmnTDBOrd/0wu0Rzl7d16L0LPBQFnq83/BXDKGKJ5jyUlUZX
YNHEEPxGf/ghKPWi8BRnL9M8a+CuKYp6hZg8mZsqqO1f7XpsPbaAA/mMWanJiddy
J49Y8uqeAXsjSrGfqAOsgGnBccTgQOwjQ0IwwnWGfM61hNCVCepJI7k+6tb3aXSu
Q6PQCLoJHKXcHfR79kvKVSURb9nd6wLW7Cki7ZuZiHfyNCcVQEb7Gktx/x+uB7Jz
JmcBQIU4CC9DWfN06a5o+29lFlm+9ZLUj2cWDKXlC6FOTvAaxvqEMXe15fWjE1YC
zT9tsqk6FpgLjDXk4TA2CMdeLNWyOqX7USRsxzmIzEHDx+sVdGtXUNutMEGxbl/k
rf8BXObsJtkeCNvX76qsD9UQxAbB/2YkBAJQQyppoQMWZZgyre7qDAYK37Ni/0kk
ztd5dZJcJiYwyr5TsCpVN/tSiUSozg0MeFgZ4dkgkeB7oXf8iErynLvvQA3ZgfJY
NNfhmsUeszJaQ9XGOLFkszGtUYxhmuKN2oVhtN5xwMrkiBO1hZh3saxQk+f5cHpX
mIW9Bqrx8nzY0iIccWZ+iEsDThqsx/MvcbeZj+PYhhALXNEh+npJ/W5rn3rozcZ8
acH6XqF1Ahn8cMyIJqf6AIxdpaOEXpxMjJmlBjTDAYUCxHiJu98aaxSewtsnSAQT
Rj4vPiazY6YBoXfYPXj/KyWUNKtNKOSo0jRSGBmIKVugl8P7EFzNpl1B9kb1j7Ju
7hu6IwlMisBdXJiscCS+UMWDEpXsMegUmEd54vAHyrbt4IPdeiVO+FfiLMoGzMZ1
xQMx402JoARLRYt+Ny9y702Vu4Yy1mnWSYmEqUpHBClnVGzuETG7286vrYuF6QlO
mWpZ+ppr7EKLjxZHapk0aVyZYQr3zuXaIOxcxQb6IptAjcwgN8i+mX6ruelgXn+g
CEPFUaCCDtuCnXqBePqq+C9NVuweAKPfx6zBFTKPJHEez7/Apv9ePAu3Ve6O/wRT
GDTA4OXfckk+KMPijR81AYurYQ10MYREl2meBl8+JQ/L2FkMpcQiJDI38eMURIeV
xbtiWdCSv2lCAl8xx2rhnueesVjuHy3iXsmSdWbNNdvOIZIPAok9YxzARzWi3Wjs
gnaaZvWH1MGR0Yt7x4X4eaFoDsEXnYv2irrfbeZVwEKUIddF6VBmVAYYz2WAFLtB
2L/ZL85KeX/mbkLjn9CSPCrlxqs9dAWWJj4or1BHCN2CIAwBXyKyUiXSZyxSU0Ol
3jOfmJ/k4wcTZ1Xere6bNu7ABYYofzoeYq+IYHEiz8nj2Zdw7UJtSGzpPOiQ41GC
YMC6C+CnFcsOUywG9k4a+JSq8I+76ns8e3hoJjiQO9inE3wXFKdyR3CfW4IMOT8A
jNgDiYq0/qm15PGGUb7SPM4OqxfDkc+13o/cfXwLYC0DW7Mo91/lOA56V/fi0WYY
qqOASjB31WTTkc36NcpyNvFykBnWDFYxumVs05usEDt2tuvWhADowt++ecaFGvMv
rYVPT85Vbn7sT+zlkPJ0bUMMWQ2VxDQ1f/+DlDMNU4fnCoY1gzu8LTdQn51aRxJK
/fDsmE4vx17C1GgxiqNIxQ1LxkUniHE/1EpiWvl7PWHTaxEy/v1s2rVcmyj7c1oN
/sUMqdfqhfcjqwHNQ90q6+XCZ9Ra0OEXrYQLQ5bHPiETrsqh6raZaatABUtLGRd2
cNN29TmE2e+7SKAw3FiGhnuhp5gr0PN9nK3esnfqoADVaPHhxN3OnsaF0+50W5ew
0OpiuxoguUl88Dsw10KuGedvBD+80IzbYnToHDNkTxYm5Diw+RHEV2NYswUE6qQo
B1Uh7YLSCUkDVu6w5/s3OEe2kZBplOks/se/XRDpr8qdCjteVUJwB8eFkrP/ictN
YKpPNIQwvElbHHftXFgJd/Oiq795fUC49y0/2x3bkPvx568fCVEQ058XBFGO+7hE
lImtStibhGl21sJDJ7JNrjxy9MsHQ0VJbYn8ICkAJE6e6uvOa2qiiHb0+kXMbhv8
fYnLv+1IpFBuMuw6oQrn1G/HmOKmDWDChc/Dnx1YKu3gb2u17ST91rSpIl/qURZz
ZIDzA6x7JnUPz0SU7JAbN1xVT+Qs1ElE2G5woZAwsMEywnonGyELEgr4rsunbzEa
CyjYK1FPp5fd/tuaQ6tHt1W8bSW2bbFP2R+BBnqnQYVvTjvE48x/76cbcJ3JkZub
Ybh8WwUz+I8QFRafzguOOTTxhaP0YpjW8+yG2Ul0MZJDzJ5IXHst+XW9ohiK8L9l
DnAObTGMGNcYrekfAl6uBRAphke9jRLFMHDVgR+kOE0nsDRCmcG0ShapI6f4YxBV
XoffIZACO2iOAWxeifNCqNaSutWI9b7akBRfgVZ3kXOEffcIU4O4U4WZ2LhfvNj/
Clw/Srs8y6eGmle2loQ7I2RBiLdV+Jp7pWwK8jY4Z1WcHpzg2TP0Zi9CpA2aMdDF
dzKjnZhgcfGzyS7OvhNFc6cn4d2D92XsrKTu6rwiv97XFxd1nJsQ+27pttW5ScnL
T0cn4q3UCj62E5iApyESQ32Rjnn8TqqGmBsdXXJKWzNQkokVuNvHG+9xfCgJYxZ/
VipNI2py3OpQmkY5LS9dy88YejenRgRf0ECCQf1RumjXmzHPuXiIC8mdGxdpyCZ1
tcT/xJj1mOy8S0RJoO5Q/ps+f7PKlEw4EZhmVN2XPiSLJ3xRl8Nn2Y/mPLt0DZ9f
EL9JYMjiD51uewtO8IPJ9bDDV/tLy4CXNNDu1ZiR8LWx2ZI3Upj3LgmwJuV2I7gH
VBrUeq8fgrlDVbMrVe6JWdmNWmVbtftg9QsSFuCZqDHPOdk5BGR2K979fYYb91s/
vm/Vraf4RdI/0k1fjySMWcS0ep+4vy7R6ZRxu2a3IMoG0+/ZEas/A6UGRHpS69/c
fwLUOix0+lYByVqVd4BE6PoGren0u3/C90FhA5OKMJCE3W7Ph+UUBbqgTjBnVjWt
IkS5lKOssq0mZ659Y09vJ17zMtVJQk+oLLjzYdaoxxgtch4RllEVGkmsmpL7iyDE
3PI0cLX0oOBS80uJoE9ZXAaK/xbeMgflLvdJCXqr2pFf99M272MMyM50SR0h2vrJ
Y0SigLcGjjaqM7jlawrneWlC9ha5MfKKUSNlQ7mN/TK8Vuo3UgV8IOZGqSC80BhK
5N0nSyARLLQyC71yH9rThXPf68+d5bR3fJT1VACn8yueu1g0gsIDJdBTPesaAH+T
Ln4l0bBONbivdV4aYcdClYUcpIJEsAggiQu/jwO3MLGfpOA3saQHiBPY08a4YjRS
rDy9nWoCSCg+8TO618LYj4/ER8tGaUFIJu7j0/ysFqImcjlgl7aMgCY1bOfbwqcl
+65gmb71qVZaNozgkBhZgVqSvrOlryV5r63aosi1hlK1ccblFyrSdbgRkil4Apv/
PAGaTT0uvoCBIE515OMVt3WX8QteiF8rsREBT/38+PVrOJ5EOhan8xtQB9T9hj8T
gEbQPcSzlrlolYiTu36pI677iJ6AXxaV52bvcAa9zuVNycz/droUrfOswGRr71if
ji7G9a09hon9SFgy7Ni3HFBW0rAdOPq8xFXw4NENuRHwFmcef4hRzdtj2A9mwJVN
1YDKM1L77eAUNclYRveEzSBMmNDkaLJxTBFzCpKrcZRH1tXdd6DBmLl+8NBxMzne
o71mDz7WFTEewzUJXvscnOafJgvaPYm8IcvH6MuWLYXdCDUC4uPjSUy3qCe9/YOH
zVh+muPP62PN7FQlAO1HtA0Cq/at8lVEc/+pOtp/nugfPSWk9VHP5jEenx/weQVc
KBNMCd3D0DMt6ihPgxmGmDsaBIgW3oJRSVOws2vndsPFNkVOUC9lWLeodV3vE3AH
AKwASxz6EhtxBuJNRoxxSlss6etnvBSXicgfzTlaQJMXuiCo5TGbpksShX621LEj
kJPDDVW1+wwAe5guDiUOnwhkPBOGvucwbq9UA3QpC6ZqMvRS4vwmXgzxS6uG+YHI
yUwCw9TfKClaFjzikfmqDFKP01Hop7NTlDGdWGBGhirBC7VLVHcaJqpTy0gAlLZK
ANQWTS37upSqDIZqXp/KJ0SEnAoLXJW3xBYEVGDoUS2Y3yQItefycl08zQKH1I7a
AeR+NUZDUFu8r29iFQNhutG9GoLgEsvzwQ4QCuABldbytOmXlrncVMMKWJYj+SaQ
yrdiVaR+EZ4GGR6dwVWTIo7X/UDuXQaL1/3IvedS/1+GFvuowBf09GK5nePnsySB
ogSP+CTf3kX5p/B+7MWgy8jwltUi9lF9WgB/WEENWvsG5GcGXt0PZ/ynzrmIsx6R
dNd8lSdt6yPK8/KJ8a38g7RoGj+1U6Eg79xC1LwLSY7E95ujPltdQ0Ibo9piWRuT
aqjKVfpeTJNrFA1mcW9Qg3qlIQho7EZw3kyZzR4BgGwFm4TAewzvjwVf2ph7d7U2
cBxAR+m9dXt+6QLR3tJRwdJ+S5HZ+ONs6DlOihCVrJqqP7nADaQiMyNSbcg/JI6e
J+m6ZvhjLcuAv41K1mkMmB38r7+UerpSZzXIBeECiriXWS9WnZS4NFnKHIfPM+ln
Lct4GCheCFpOF/jiXWS/PnQumku5lWRYPlvvNkNvH0I84PITuZkEHEYEHDSJtFMc
rUA/zq0r/fzFWKa8iAgsewVcnM5X4FeeHNDST018Q35+otzE51X+M3FcrYcn6U+C
DFAZwpVdIcAOg+xSFybc+t0/m3GEVAkwvb5eqwyGMw3GniskBMoAZCBtcH8MWOjv
b8avUEnDLxKbU+l6CjJiwrbzUx+QR9H9+82wZ1n1wZ29sizaDiNpjXgLQNSn/A0D
HaP18YOrFjv/9eiZGxZ+HXkVEzSD9VSLBvENm25q4eSYZOEdojzFXurGxzTEyhb8
69YqDo6lfOM7dcdi9J0T3y8Ef0l4m8+5FmQjUP23JiRyu1N3KHfVu8oH7BOjyQWN
CQNWF5tI1WGKjo5o2Wm4CEaBS16Lku8VU6hmjicZqR8dQhDWwETdkOIlJHBVeKGm
smumVu5EgUVMhfG2gj1YOWP5JgDWyVqUGTQ/zGJZsV+zBego/ziXjtkOx3UnHIic
DNZzPjMYUa+fmUxAxP+V9CzMnVvTMGXmJcARlkwjsbrDD9dRfxMpW7hBG6DjjnoV
c6+z33FHd1FOga/RfaxwijFAQLK5PP4RwBzscmey96nNXeDw63pp7kM2JBT/VgVL
dWxkl9EbgXkWcj8A1tj+mkkp8daFDwZl0Gma/pl+m2sACs3tiV6z4looaIc1ArKC
/xsl24WgTQ2sfX2oochRPzRRED4Oz2dA567DHLiIJeZo+iCBjEHz89xIiFik5Nxb
hx6Ua6IcPavqpPItShrXBCfUwCeP4jJ73PgM+dKeHXelS1AvwQ+tmDfcVQcVaKFZ
0/vQsNoNL0q3vSAM1YurWEXz2ZNdtyeuLW8s6ZFkvFND2X6qkh0xVbKfj3AjGE19
w7knetYlPKr/hb7hypq3Z7XQcclNB097N6jlyUwT+EUf5KBHljmjHJ1NPgJ49sCO
6ltvVI5zTPIQiCH/Q2thVuSNYseH6okcE9xsbh3kiO1aPJ3NtqrYnjURnOT8o9dx
s9H0nsBWwCIS9m55i4FOWuLJezl5wzwAhPyOnEHkAiafm5lFvCb/dNVsZfJOoaY3
WL23wjOXW4WjW8EeJU8nKzkHrRKLYhlbdqKoXNhbIz0o5x20ZgnDAqPnYvryYPsq
69WopkfyrMh9NJndOaMhEM4XLH0XWNoSvfRs/tAa4fe5VUtopLHrQlQfP3IpqXJi
IQOG7o0Gm4hili7qAcTKrBGkXcx+hOFrn8JfZ84IFs8LXP4t2IB5284dNDypmzxf
ScY5I2NoyyDUa73xQEQ2eZPbBb4dL+d1upbcxrGuxrLa8q0k6ImKOCXcRXrbzQgJ
JAlkXuT7+FElczuOTJDt8zSKR+jLS1Loce7EP9240z72j0pS7G78qT8+yRRfBDPu
rsfPOsTSKQIo6zEcG4BYBPq9GhJVUC1T0qoKJCt5Preye0GxbFcvlGz+v9lEtPSB
+wH8pHWOGp6OBdfo7JzA+qhaHn7GYDRPjyG4fBP92gYiCNiQqGM6bezyRtlBGAf0
TEaf8G532fH380+DfAzMkCOo9HrSA7kRMkAp2ZgLP+CSBNJMcAs4NguSym3fqq9Z
jVM0vtMTCFBMMs5irJ0V+3OGK1WyFnFwPFcQOnGvfeIj9UICNXXZEsXZQsq5c8P3
vmtnIf6Fh7uAk/YOCm9NE4l+VN2sBSUwZ8IzEI0FD3E/7ZsHP4FEyIkvyTuETlmy
Bg1mWf5RwC9bfV3T8kCoo88U5S0SaRtWLQ0B4yw+/bSdtgwExh5n7zR2S1OozcyA
1QkImoVa2sURbbXMdnNyJBq63vD4tfoi0OwZ3zw8H3QjngQaVdeRwBog2JSPQSRr
q0FkWp2cbDx3h8PbFDZJWHDZiTp+UGsUUhgEC2FubonBf7Xmxr2lsH49PV2InUaG
z29P1fS9cXJ1Ulh3RWpt/U3QSE9y+PNiNQ6T7nMCa0U08x+l/oruW8Y0T0Vjf3jV
+cdNrQMOIw6PHWgxwhOrtH4jG4qiYJoyNGLoR6n36mIpexuWubUoDSAZmXIyEhSc
YrY8V16QXvfJ/M2bbvEJbjerAgD0iUh7rqiUN7zFyzsATeGtWHfysu0JU4+qvWXD
BrRE2GV3yTzIcKWgp3BVc39VKxDAafyPYhGNFl31095Q0Tz3gvRdCJOngASBt8nJ
m+YIDajAjXnRX++jAfL+H+YLdluX9pAzbllQN/s8mllzzrLFoctrLEH7u/LNHtfP
Q4istyaihrgx+bRnVfiUwGc+Gt960Bd8p5DNvG1bY+J63HJadMurOmStva/9G2AH
E8QOPG1IuUVaham8uP2SOrXyus970yvP+PJEWaDW6eeSjP8dN/pjPWEtw8Utqrpa
Hepa0zy++QrQTAeT+B3Gl9Ug24Kn0mEsv5KyhG7qaPYp/MjCynOvzkk4m2iCHwTR
+Y//ygERgFrMjeOL+t4hqku8SdxZlLJ71DF7BxCer2lV8F6prt4j36At5lKJgnSf
Mhlcl1RRuPYHVvL+fDkULRtdrMRMMsrR2qpXoOhm2o0BGsTktMYyQ0kxNSQkmcXT
WsOnDMwGKA4y7o/lREEgQAOnrnsO3gBDpcbt0y7cjGQ0fJlCMtHO2/f2j9W9XzfZ
Y2bIcIu2WZV1b4VzbJOMJwP126Akvx5t7UzXu/U/b+QnZ/VY9tDCHgjG3drlMDWE
X5qB169CnbV94IHv7XOc3W/gCIeK8UDGZI/95SmTnS6pCoXCUr4ROhm9udNBZVlz
yJLc9CL5bQw86oxDy2aN6e205eN02RIORm5btied0BZWGvYroEx//pXd2/k4dqyX
99sg8TiUDqsMv3W2B5aOSSKGnuc8tqsDAllrnMy2howaWERCwYcO8DgmyoDgMGRc
JA13f2HM58LpUe9FmNHc86f2MhH4UXd5DKd7BTEfyXNe7BxXa54mqPNk31bwFYDQ
LyvholU9D5WIeXPMcdhcQyRr5+0pCX4s1UmSAtcRg2gp/15Csf5xWyLKvwpjr5RN
VPWx9O4IekJ4+Rs6vbzItnHB3KksM/CXKo1QupIhuI7CdJtZud3CINDmpn8pZZ59
Y8I+WOwtNju8zw4n6gsL5QX9gSUbm0icJXgtMQczIjpKcOZUGxy2augltvwZeKz5
gCLJ4CCpl/2U6jCm3gpEGWrSHwYmQl94zYIWL+MAqqqt0a4eWobTTwbOlhr1Vwac
1UIE+Wfn4gEjcCGBR1s3vsw8J2ak8OXbxaFwZ8bA7uCCR4gIEMLGK3IrO8BWSMTw
C5ZmBk0V9IpR/AbQiL1zHwMKng3qEt1IotjM6N/i7LDKkOxJmh28cNo+Y63FJgeQ
enBcep+4H50D875S/5fESvN6K8CgAfikJBQhtrIg8LzzC7N1cSn9B3Zj4QWlOEmB
GbfD/vs74dvh8UgmD7g0Q6a6xvtFR1zLC1NFHVEKDzdtQIYbXscHNv0MwdO8y+J8
rZwrBXDd20rHGL/e3O+BTdzthEhkEI+fOlafvURjaNkRBD/F8ep/gvO3XrpxJ97Y
9oTPiQfzjlTf8VL1g8VOHxYT814bYSoxSkiq72mQbWT77qvrD5nUmzzpVQzSECIb
i/Bld6GBSAi1WuM8YvZahckFpbkCbhxo0CCBd3z8Cf5lGO57zuttglYwYQLdY9hN
gZUZ14qSkjhTsCcTKDg1senSqlm2dDHlvSy3OLLcO0RFMSAMQ7Yiw/zUedryZwC5
Z8T6ehfKgUKlYHZJ96avzezjPGST/5mH2smkiHq5LSPzBL/hO3UzZiCoCUqz/nDH
Tw8y8HuNieylWlCbHS2bzLAQFLTsez+6xYBA1Bxgt3xL9U7/SRgJnPrGGpbKFFpP
g+MecLmCWFqqwZYQMM9CiiwQpjNu2/NOpxZwrZ41F9hJ1WWmf2MPiBDJd6/MIVBo
bIsQyQTG/Grew1oXuCZR7QZME8efMZUZrXU9OgoI0n1Q2aB+r2PQEEFpAEs8eU93
VZbFxPX5O4VUyN02Zw9pQhaI8Cd4InMYp7NGvTa1UVt2DXDeNjujQ592HzJd9YJ1
ruVsmclG6Ycnvl0S2fpO7qkaXjIZGUl3DtW1zRn4Q0gsHQnBozAXwWT5ac5NT2jj
si36RVU1E3JshLw97Z93VRP0bX6D/dZpfOURZpO1wx0pHDLqBIhGuFB2egcuYE4s
XqUbDfWX+U+0CYSthIlGYYtc34jyiKADNP0BVgoeLGNUiReBCAbZXdgfzb9xcOx7
Oev/1V9ZNuzUSL8o5IeIOTnQb+Gm9EesZYRVEqm0XMgWBB/bXKlqnF4EjwKCVdkp
d/5RJK/uKHKi5/Z0EYU+9bJxj9fWgaJPwVZyfIUNO5RWCl0DKv6Bsda2pCAbrbQJ
n3x7+/5LfaCdxuiA0nAXrcqFkAkObd+w3pdDa/Q/whw6bbT7Fek5jUq1iL1PL51A
kHx8qmhuAJ7C7R+khrSKn8943lavVGNIrw6H9iAAQmrSA/oNmeEs/oNvBnpD3AlI
ITyYFExzxdMUq72dblhhbEeVBhu+NcxiBFVn8CQWsAtexcbKAyWddsMXQFLsvVIG
BtILO3LOHCRE5SKN85+bxf+ZUF/j7uipHmxe0fO9f9tmIRk4a34JZDkEcIW3Z41S
jFTJqRV0urekPCoPuaWXWKXHdw4L6RrogDOt59lhVsE9yx0Xp9dg+RLy02wR/G5O
d7O/C3i0eG/GMmsoFQGct9LlJBB2M0EwCVWAMwXHStrfdzzAn6NGraProGBzFFwK
04PZBhl8r9dSuPNzTqN4inxZYO/m7E9wMjaBxwLhvrW2QOh7uw8VUbceAt4vosJ9
taNOLDYIJHYrY3sW3FGFYPXlBJm7bGeSIvsgRXALMYoVm+QGKEiWZle1ggcht4FG
S9LszZ+Fhsigcx547G1qDgWx7KyVpICty2JQI02FDr7nZM2eTNhaLmvcgtPyu8jM
93jUZtxdjVSD77XY2U9PrmLAjzY9Tl6z40Qi8PFr81gvFCYeu7YXFidOijZrYhmD
KWgp5rsYAEOmgzQLDnBO/q1ZTXt+fWVo3tF5CJCzPEE5mrXYlMF+pm8vYGpkApNT
DfE43+28enVJOB57YJtbmJDInc01hjRUWZ+Sp2liB3HttQBajvGHyhhYA6y8X7wI
ei3JgzkZF6DJRh3OQ8EDflBUTzZS60FpaThuvQr+BvmWo7g6h5y7FjWUEZabkVi/
9Js5fxNjV6JAniipYx4fZ90gM/zikwruzVjKSoNMf9ZAxrqGspcZEswqCQpm6gM7
UJVs/ERqQDXHI3juvQRe7zYa16kpByStYKv9OTTgVW/8qP1d1LYQ/XWF2jITtZ+T
Xn1PfTfbz60ivMNxISbEy0utsWYESBHoCDtHwmfvnQjxU3X5sSnfD1tpQQWjgu+A
jwuPmLWboJ+EiuHiTLwOYubYwTCtO1VFeviFmb4j8OWSDUukHIfLGxYB+nD5N4Ne
yi5N8I0zNHW4mxjanyKn0q5bOzu0Bqc6T55LYsp8LJ1yaQZ7E15HHWK0NQFK9r/s
tPDYXrAZHwGF1kLJt4+AVJ6q2lMjCC1VXylY6uo+JFeM7HpVLkfHOWM5qRqCJnts
grw6YdXncZdhVwg62j0PpOIeYPRUrg/rtsEyrqGKH+FH1Vfr/PDGz8y8k21Gw78v
C9cJ5KxxTKz7E3rTc/RvAwMOuFXO3qgXs+rz3YvsBXaRTEdskb2ZGe/Y07wNwc+4
8jTk9mjkkznndUpNu1ADDfQxGAbEBQZ4c3msCvSiBiMPf/L3ab2n/B9khqhBw+hn
Gx17z0s9bqmd3fbnVk8fQhqg5qmp+3G2Q1DwymMpoRw2MPnw2C2P5CGskooWaxKa
6DnMvIyNlsCtbYoP5LRqmZ5bjfZv2riIeVnq2f5ZjoyQKniXUSOlh68wJOlhATwH
Sbjo08tvHkI+zrkJiBzg8q6+1SU1AClqKR1mcwO5UKsuR9dTXk1AyHctKS/BcixU
veYQXwmfxk3m2IgmgRLvJcj0LJseFpHBMLKUe03a/0meFzcJasTGrLBcjzg28xdp
itMiaC2KyAuw/PlIu1Yexrob5tuKRLTvqMjYxGpctjSmwlR8+KbHQgVbP4GYfLfg
ut7JkH6R9a3RjGuNAmRCYS21fQ09NXUoDTljQOz/aRTlU8YNHPgJEm9yTLhGPvog
uC3E0CxqGfa7NDyNT9H3SCdxYWOcGpD0vBSk7G/FV3nEpUeiPL8cwgXQ/axy6mLw
bcB7sMwSvmz8QgEbtSJx4jpaGRIY2/gxB0QADauGl6VwQUxqZHtNIvkJGy1a4RzD
8v9ikGNyeo5iWhGPq1frhaM8pp0wZHxiIvtyjCiFm06/zwMF1dyGzxqnNemirguO
jCR35qYxITsfZ1Wf1RvcA2HHXzFA+0PFHzNWv4xjGuLMI4eS/WFAtgl4lRxoiXOS
DLyrcWemhT3GrUhfWsDzQgi34oASP/7WMKq/czqKJdhEiECskraAm/9EUY7M/BI7
el56b7F7NelXzl5ubiZPXSEa5una5B0MDW/xfNSt1IRo2dwJpnYQYO02pt1GzWq7
H9otDxHMDWop0q42/Q7c6OR4ZV/or3O7kNE0uYlUq6DvnHfr/QGcuDnPP+oMoG2E
QYac2Gbe13m0TZ2UiIdsjhovUJwXJQgGZLVydGouvkcTBv7EKZ6JYMYfoErn3XIV
IP06qnxS5pDRejo7B6SHek3pdvSjr3eXVsXtiTDEqw/LSD47/QYjJZupOzEq1KvP
YDNCijwL4Cm9T9JZ3ax5/yN3a40EMTQqq0cgucYt3hcNlFu+Nm+R50nmG6vmY9qx
68Sjrh28x3AI2/LpkNqVNNOSkGh+MxtC/tUJ4C0nJtkc3RXQkaivXA5UVzzLKF3x
kcuv120SDfY9tr5qG7WbG5xL1TvTRo7EsNiyuKuFRHY7Fzx/FfJp4ivZHSNz791Q
f597HqZ9ycmZU9QCw7diRNQKrVspcQW7FXZ5irgdrUi40xZMO/3T0nmcuZB6KxPH
uyWa+7sAJsQgtJFyAia7Z2JAhSjXuJql/fvycw4+oQgyL3Hjto/Yhtqui4KkPi3w
LPJzGWimDBmho4E3PNjkmJi84wT6xZrLUME8QY+7AaJLcfokSIy+K0vbhDiX/ZPE
FAUdXxkYTkXPjE1ub0RK1nOiFRxt67XKodia2PZa+PM7mrsBcFrINAYJ5hYHVh7y
Dn5V/Owa4nkv2f1+VjY0rm9FNufN2aRZxp2yzyOBXNutkjP8zSJrrOgXIPBa3D2a
B4XJtnFxv7pHVhbp4f+pn3mUDAsHZevxoW+7SJWl0Qfp0TSVjR57EVf1Oc/9N+TL
Jfl+Qj/5PBbMFHMmFtGdluqZeuGbJRdx2IHwnOmDGV3rgbHt9q7W0t2BGL4eFU93
MBdYP8Z+/gBji9bVEdjnvY5h6SfuK1EU9uOl1iFWqNK45oGSFy42Mlcp+zOoCYcQ
X6OGBVUxgBJCFMoplaHVXWIwRFxlK2UPEg1MPrmSd5BfyosKNyishOQDxFK5GOwb
rlosrS/xzr6l43DQwum7VVATbZM5dyW5TH4SXtzOlF0zHUMCY1ov2J9NwqkQMK5/
GNgEKV+0h1KI82DBRf9NHEZwcy5VkR1jvf7AtQuAZTjcLBYHMx6doQ6PUJXX0abk
719Yvh20ZqZz4N/LPgdUE9TnnSM8xMb6BkUvf7zEpY92wuqBSn1dLm580oxthy2D
EdrmXkadkRdGlHCFsjjftv3gQYFVjZDkclz0b0KRzMEH1EBx5ikTgboRl5kGWrFq
YvxbG3KRnsucucNSdaC5XE/narBk/YHadgmq7hP81G9ZUC6CjaJ2rvoGzNVLo3B8
UUtrNPmZ1cL3ZxLwX+nlYunKi8cjxm6tgyySLdDI47f5qrO86ISb0Whd7r7tQiaM
92DqaxYRMy3LXVSRSIexdGfatVb2Dw7qyVeY4TAQyAEgNlkYDUFqHd2eVhCyWgR6
DF07+oMCzYgJ92bBKKSDfl+roaAH4Db8htxo8dEPp4OLNMe4eNmfQJlrPkHP95NW
Goh7lG9t1ZQ599VLmyd7Fh81/TnHiHPmgnoecJTwZfB+EoIoVhgWhYHXBsqw+YDm
ZCwRi664lqxqB3MnLnqGeyM7IdFn9qO2IBfBycQR/vjQBzEPdkRHhMKYmwWTXA1q
8aPFy2cJ6rpeIp8bOa1Xa54cliEvmSziF+P2+bvPw0n5AP80j1dzaKASwAQ4vB05
5+0YXeFnOhtHoLL7FfxmvDZ38L2MXNF8hYX0r/lur17JzqVGvYq/PHCVMny9QIiV
daljxUZyZ/Rzz7PdnnuVZhAAcMdMpi37Ep5YtkTiic6EPM8ldbbw+Qf5B+MohKCF
QnudUihKq950SL3xRL5MjF7U+m/X7ZglpwV1sGGl95vj8agIwcqPArJ5mFd3X8/W
E8ialurixq3yAeF2gN9lUFo7/d+3f9+i/nKbaowdr1wmmYQzSkUjscKLXkVoj/yf
zeUzd0Dgu5pYxn0hqPiDRDRVgaujXNyUFntnkzNES2EFh/J1beEUGEmg4GuWkyKf
sxWUuHKD9fyiOZdhURfQd0vqpie3wXGuSXaflZJUBuyNscRR8nD7mj62LVcKC4D9
IumIQib0P/ruFWlk11fcwqJwe+LLxXxccQ+RRREsvJ999a04IF1kROSvpaBdMsPC
cAS8CTHMSuwlLxQ+c+6THSzQtC6XnNccSlFoFfVEEofT9hQgqHN2WjEfolEuYa8T
EciTx8rQyF1IRmAeAAPFjZvlde+Y1bfBK01v/KIjfAp9xoBBgiTdJYv24oY/BazD
f9j3d1WQbhNrGZ3pEXuvhnxPK6uD3YcPYAoQODx9NYLomYfJ1RbvrHZ47CiqAc8C
H8awe2AEHW6aD2gYWqLvOVOu8jTwiMxYNyk0Z+kxa6q1sPqNmg7JEi+GIsh25rXq
0bF2RNa9ks4wy+w20Rhb/wT76oqk+XraasZWHd8wR7FgyY/VRloLmfuO61w6zHGR
kSSezD7H5wWFEjaaBKOpbpPqPEPaNzOPM5PxXfjR2JefQ4X1V6JCq5rMRfW0RRpV
lRwvNllSlYfnlkf5pE65qKFbIjfZclyiAa/ysKqNRH8mhMB3vy6coclW2ccSx0AY
JSlS+vW2rNwuYPRbscAnm5xX9tFku2a6m7UtNxwxLNQEpVEf2DPGyKpyaE9ElZPS
zfv/BwFBuK+aJkoZlWlvsX8y+R2+4F8w8yZexklfgVcZ/eEFYDHAyfFP1YSp0jmb
TlrEhSCOW2985/fYnCecwqX1u8BMLl+XjxVMUpFAlf+HurcLQWiM+D7Y+WU92IXp
rJfkCLyV+RXRhwT8SdORtqKbK/eOH7wfEO+SiIW/OzQqbT/BQhhufCccF6OFd99n
MpkG2P8vAYO+MxXivTDp0DaOaUNn/uycnGgM6o3aN/mCg+YMuxJBtkBJBwX+3MiP
MCS9ZIq3PWRMuyt2ABEAt+isMgI6Xpx7h4XErEDFXk9UP2bt/STq4EtE8qtlBMox
AUrQUt7u36fmR+WpGS5Ds9JCOa4Q1SjB7dl+C0r3NFU8AE6NyvkpwuOY2ejkp38B
uJMs1zn3C+DZMEND1v73DtFAw1xrXdZlH6rPZVkAI/u5fGMld74d2KXX5hrDrqsr
KCVVjd6ZEM4epvqPXRfCzpua9cOZ4GsUWz/l4/wptXn0t0+ijJorrDyFm7euPQDj
7/hPMtYoLZSeACk+z0kvKAMpc4S2qLX2llZBDNkIJN5nIv+QibMDwDn2ZsuW8Ox1
KuKqM12IkUyb0M+PKGgaSj+7Tt+FVjTXTmTk+RHrgVEFkZi1KubIe1X8vFFqtrz+
lrpg8U/E6AeCUWCJyYqpbdbUxVIrVUsRrxs4aDsAeuq/iPwJopaCkTsEqsyjaBoP
eIIWn9knSEERHxArZ7fcAJSn46Dh9bUVV/DfxYFIgdvJ0a/3IvgdhPgn6tt7vmfp
dMi67N2rBkHM9cZgB0atXLw8cN2r4uaxyg1qsjlLNX2bEzs/ZIswYfRv2z561/yd
sT+OUTxd7NPx54upSb4wNRzh8fpZo5Kua4YN1dxFqWB9pN8cqnlh+x/wXFyfhrjd
Z7ZG4Lx4fDULJG0w+l21I9LLj92TKNlWBfl4xKsPF/8wuUG+q0mnJNyxsQLAqhn4
D4MDwZX/1iP48/XQPcHi1+8/Hao/5oklDo8ZN7Vm6PtDK+T+pgsB35qQZvhwjZmS
HRdEZoKjuMd1zrDrUaoC1VmTqVQBVWqjMaU9VwepNzLlmChKORGjCIq4Sert1NiB
pXjHN4b5dbtqkC6sAWRfJkyzkad6QjxqnGZVq7j338Bo6llHsoCDh8YicWuwp6ri
SnUhiuVDzEujYDTwlvQXuCEsCx/+WfjD3oBWxoW2hw+VAgNdcfyny7lXfltgZjVG
a0hd9i4uZ/viA04/gsrKUjfJ7wupfEk36xWfWxkaPk5x5HUqt36o77PYqHiZ86AB
a7czhR5uLbALsJCOLhbwHH3+0lEjXaRtXIlj/ReIYMRxgHDDf7nSD557IyniOfKd
MkPmhpdqMZ8rWqYUlKpjnrnueJ5jJhwgHewp6XXvuxp5nb9nR/NTYUUqACv/FGH8
T78wX8E8xqpYn4lpfFcGEbpWFjFwY7jw+BO63meoC6CdEBhorFGWDntCPzL9F2Pe
D2cpVqRKzNslpjNF0iRAE2B4FT/wfJQvVHyiI0yIxSmgdBFFAl8rflQBr8Yntu+z
mPZaNhgyPCiqp2L20YM109H1TQZq7KYpUmkM8wlAGSzbdcu7pnpoMr05VuJ9A+ci
w0ih6fi/XY42j7FrGyhgRpKBktlPZgFnsMEWsVaQztHCSDFBOTQz36troa49iFcx
cBcVXWCgG5W+ga1vBSJH5u01sxLMoloDC3z4VeR2heHtC9GViuqbGXFQNQru3xbx
LM4nN3Y+SfDBErpgd2QtkWAqP2bMLj1zZT06qf7O1mvwdg01ffRJl9EwsEa2MRVu
m2wbXTpR2gwivQHgimZSK5KbeJ12G++SNdEU2uMjzrBGHRYuCTWNVaqJ9fJrImq2
iq5R8KqllOoPNLGpyoeH1AECIP311oXQHPKLf9oJlIntheEq4pNjKy1gmUdqx+25
Mrol5aBgAdi9CkQTH3LuvLc8FUD3C37U7iLOgXdbPLDrV4f2uWfzhGJdhtHO/6ia
Q2WxRUB46x2uUfSWf14v3Mj58TnV07M3uYBvB4+Lvkv1a7fO4RhbsCZQsPbjEURR
p26WpiR1GhySxq7JJHCRY+vbKYN8VoLwE+ajzTabZyrgsgxkquRcFBeKozQzPdIH
AubEjwunMPVecqMsCRHfcTNYTDBXv1VfISIQJiNEqROb/6QzyupwVVMd1BqsRLuK
XbeCYmxWApIyQ6b8iGOccuVKPqQ/WWEByIsJQpwLjunZN/5r7kMPvmlrdI4drIoH
6jKEsk52sw+8RhZgwQnM5HRLUbTAGlHQlYOmV0ZPL2bcnS6PlJL2/d7H1XZsXpEi
ZxsEbSuI8dx2EVOQI1uBe5baTBBs5AXaOtKgsJejVQmsQaP4vbudCDo6LNOtBadb
o2Nx4zUaT9XU4mFTDC0DZodMEGxXg0QKQ4FZNcta6JFoHNEK8rUy0Gh5e43d4aw9
6ZBvNPDHUWUpCjnw5cIjc5eB37Qwd7OZwfFbq8EXPeVVTidmZszTG8pIQUhx1CmO
dOFz88NMA1Oky2+KyoMHyyf9oFpdJla5/1eaSckfu8/V04kjRFlNo1Ku0lwVoxqK
ye7e0fAq474yHzjmEgAaclO5hsdkLp9ymb1q5MshJZ5gw4nYXc/GdoVXBJnzBv/W
8/m+vhERFDTbpVmXYAFlSxInycOeaXNPBbBxcOwCkD4RwtEPt8CJKpurIA/p/4CK
TjiUINeF5gY+cCnShrAupRM1mzuMzllHcHXKUSMPlYiAgsErQDxcnh/UxQ7Eia9r
eD0zMTrUYCsHIRhiZiYnOiPZUOdNaRyRH4dK3Sgx0bESi7nt6rK73SRs9zF8ZiwI
YAYeEFGwpFdFTeyf17xNGAugOttcpVPvAGTbKjTmISmSzeEaZnYxT/WtByrf6N1n
Oiil9qD2Y0Bk1nvdafCHFOXDHN3BHsg4hgEg+Q4W+kzAlhxlPik9cTQM/ipwTJ1I
+ITm8H9cF6MoHuK5OItddf6uOk6C63PjEA6jUyGpasDwf3JFYPRGCc1FgoATswoP
7Hk34Ii+zzVCBsgwd2NrcO2Min/Fgx3KwwKPCoAtMLd0K/lo17BZTWfnPHbMeCsx
18dK51+YnnzMt9xwmu23YQGZDtMHsn0faSL3+L0lqJ2+ULBd6VnV4gRHg8u96B1w
v5vvV6GZoXOvNdwJ+vZY38WnVY9jO6W3wz5VYIe31GJ7Su0WxCdXTUF8sj6lWCLg
y+vxZbxEjXUBdZ0D/tD7/cBttfeuiko2RXEDa0BZvNuhu05wsEDxhzSBEoctu8As
pTJF4AdO2pvmd17Lo77Jo2AqkLZJ8oJgKTeR2nfQImFeGL8+8gd14hDCnJ0TF9oQ
Xrndc2Y8i/m72b0yxIhvo6T5EVsZK1tLJX8kfmqkkdC9YKsl0GUZFqLwseGT+oys
Q7A+bl/cPKqnR7J5KizIIhYXEfI7qF3dAnUPjKcIyWm55p4DMFxzemr0TJEh7Xu3
4DxsWrXH01IKTjKawVT6Stb7PdKf6efYQiHdige8UI4B2dQWciuxJPlDLYlVkkTV
KLzgueYREIKVj/14VqXnr+YoWF3nImD7F4fLkeUvBmi35QnItQu3vRW9QLm7d5rk
XDMeCfDBFF98/cl8Oml6rJFIe2QOoOckFJofS6r50Pfmn1M97Ozeldunsyz9CQO7
7We4ix0T/t4AU3hy4A5L7PA8I++rn2lxQy/hqW9o4c8lg5MSHu/E57CkcDCNRjHe
4mc0XZ0GI215uMe/dYSgffECIJ/yVPMblmyB6Zl5qs1uFPafwQD6U7zFHjljwq/K
yjq6/C2iQooudwFJqbOJso3gyVUch94N8CKQyuPt3fydl9+MhqpdJprI88ib3mx5
p3JwN7gzYRFbDxYmOBNGygrbmRy+gH4oWHEH3q47Xi/h14HAsA3JXhunKxy2z2GB
yNS62dCH8gjDl4RbwHBw5oofld/bePNDiq2FGXZG/LtdV+ek5FW2zl+CUbqUAQVa
WLnLnNythA0mMI29Pl5jKSXPDeuDMbIPSUC7jkXMbjaAGdLtiLqzWZKca2Czoz4M
VToEgrLEP0fB/JHmoMI4nPIyvNkttnIBkQ0fxbeHypxZtebKud9hujXacOb2LTlk
De4tDlP6tnHMFzNq87FmFg9hQBPX+KluyzSVwHaAtRw0jPfWh/iW5zPGjj/T6ZPf
tg6qi+x4uONjF6/LbGyHd6BzN8+B8dqeYAocOyZ3A5o+9TxZSG2uZMqDIMv9aAqA
r33QAWzqj2nfynEGIU0H6Q5iB4Wv4k++9da2gpcAupLwLtaUZ0u9/jeDJOc/HGnK
wWBZx6EtrpSprl6DzZNtckYw+kyeP5Rt3o3APIxYplB9A5bxoQ9CAr6p8RWw1DcL
ztC6cUfGnL3KKS0uV1ciUmkRherolO+2se5RWSWiSS2ZGoFTE2nB2CjesAJuNtYO
ExMM2z93z66Kkad7w0yoCKYiAasF0giVW+/cPgM1tIN1FN6ctPGYBcrpPQZ2jaMY
VVPvH8vDUr/t+JLg6I7GzSV2TFObeqMfjIig71UgdvH+G2rQoVApOOK4i6tA9XQg
vIJJqMpJeQZH/Kr/5VAIHbekpqwZxkFKVfgOX2zkyO2eVWfiIdCM/9RDdPD/tami
3Of9z5TZAxYoZoHJB+ZzLajIajsqAZ0QrGlNZUTxlwYKr3vaC+OK6hjRJ+9XXycg
etqqaD1kHP1Q3Vizvi3f4/6iziytOduYRvJFjALqnWyzAqBFo1Yg9SsXmEvs+JeY
HziDmk/opFr7Wk91EYzlaVaqW1hrIhzY0bJIYYeCOg6PL97zOySUdsZw24DyBtR0
a0pcFNb9alqd1BiCYO/XaSilLttIcOPDTdJWnuDqXSTReFSzGwfa92LfWEWTQJ/6
jcFMq4OScb1BBbIhiJ8LRBihARgCcJg86LVeyBjCAXuRmL5bP02F5H2kUPZ5G20Q
y+eGrbuo9uxDrO+rOtMNMCMgtVJUpNwFM6BPbfNvbRvRIyZ7JbSX8WtiFtubQyP4
0fDcLGf7r7lRaRTCOL14qOs2nrcFSQb4cnwlmD3CMIagJS28DVIOZIE/p5kA3fig
95sEGxTHJrv6VpkJlKLRrRdMTwWIDIGKrfcVdWfxlWHSVLOQ30wuQPGv2Erg/6IF
Q2JukOrbP+ZQsLvpjgJfbLtfNsTbpLlKV2UKXH3caRrH1zmHxr+vgkX4lmtAdmMU
eoz32SphJ3/LK+YKJJxG9zCSiluMP6Oq1e1UOEFWA5MmKBuFUuk4N7KkfWzSq8Mb
qIlBYsGznGF1NSkfiRUeaLb/oRE9Xh2+1UXATemsHxCig60o+Gw9FqzFNyzAXBis
Yj6raTIwxwo4MPU0OX3ItcnxOZq3Gbs4cTVuwu7DbYMyWfrhwrPXpt+MEwCM4P1H
Skw1MVmXMzsteEDz5xps6QxxGHSROT6Zmxp9k77Timgt9k4iBfLhzdFo5kIuOI12
HaNMJOdgtq7ssiyJOhjZpLy8Le6ym0LrEevrLGg3+StZpwGG1A6NjX/77ewZDhLH
06G0k7Oa4i415s83KcTZQ+MgkUgTX+OLW/vaQPNp35lCuz+PE8wao2Wg4UVYDEVz
kgvZn80vPnEC7aOZvDxBiauciid7k2QGucJbCUPBszEQrUCfeAoSC8HBdKo2Zo4M
b9YAE1XfaY1Wqq4qwhGElzGVCHezOHBTmn0ajUyTHVi8hMb2sCYBmzsEfq3yg8GS
DSrQ8DMNVE+eNSUknsFsL3da+tZcDb7pwGGNsjD5hqVI/rF1XO0vX41TJXPyvf3Z
gPWzt77lN2hGkXsUKYyofp1wE9J+1YwmxR2qf8xquOio212FkL242rusJFg1h7WV
gsgNr1n9omhgYAbkZKahIj7yuSHaUljklaQEBkkR2kxazaQtq20GXuOCvzi4UzrS
ry+D+PclL2C8ZSz1irP4prOMb8kgWFwmb/YB+WHczOjWQ66vwBpcFCgDZtHvEM5j
X1+ToWuCwqOuZpmMMQj4kd4l8N7Dihi3d2S/ohPOgsxilx2hl6kONpXhFLW8O6tl
zqPHph4zrnbzhiLL4i/ChW8a5fVk0NjhVZHfO4Bc6yXMe/WmR/Qfh/2hDoIF5kz4
u9RG6eLpue6XrF543jCjZFLHhd0KtynAvyvomwLy34edobeXgnjPg0PX7fqbzXCP
SGoHqXsA9WQxOJndWU+Pi/BE61n199gqQ0yj6SO9snpjvoEo4SCc77OXcybrWHU0
ZtYOibI79p+KlJSTKhgktLAYtkdsARz28L9ki4BkEtRBNxkfimKSlH/hUlloi3bk
aMCOCaYNB1m5UTCrs45/E9wnegExptOEKPPMauyU8OA7oPQVim3BeO2HpV+ukuGU
mq6nGi+BXIQ98qo/M61vXKMPUTGs1lzUq7d1z7EwlkjPTCaOzSuAYw3aa9ZP6WiA
qLrotWtCUeOaUfYZRqiFeb626DkFBLI3zhHO76BW7zIPrKE2nexHI6cWJBI4ULYI
iwnDvJ/GoD6VSpiHlzcqcFv5rKsNDHouEkgGXG56xeGWip8YKqZ/fHKmROs3vL70
e3FqbGP+5gz2KcXDJaXJEAeDb+RwFpkyxYZ8KMmrb+fVShac7tsbo34J/TxHOzcb
SDWwMOJEzym4Eg6nd4xVs1bgoZ4tvpWS2G6UVS3oNudPYGAvbG4V6QzEtEuX2OoO
nzAyCnVF6Xl9ETedRF+DQc4tEj/S5184I2jhy4mWXskmDF8WrkTlP0ATJoPLI0Hi
83Ljt1/hYsgxUrW2B7lFgFUwETtE/u6jI5+gZiVAr3fPBCQhAKZIEunv5QIdYlaX
mCAOZJY7JP6RgUqAWzIqjXatrfDcwpkK5RDhFt5gjzSiH+iatZav0BqKoIZMYo58
0Bz3JZDW5iWMI33YaWqD8KuX6HVb+rpa/m+sH1ZZHT1ph9dntTCf+YMW99cY9shn
EKcYEoOu0bz+ctbP7RcPs2p6qn7Zlq0uUtjIaps2SlqNRbqZeYZwIkNsF/jzmXCc
BZ8mtJrm0lZ+kYur8fW7vHBCQfkwwF5V83QZPtuqvi79rVn3ClSmsSjC/qymGhPt
/Okgsv2+Vbf9K90CQkqWJ/PBCBBYhLz8XYAR+5+Ui3Ymmx3iETd67i4ewSytGa/Y
cMq6U8aZhXRG2nErb6NPuqGVBcE1sdSQ6ISmN4mxKWHg3tJvxGeYfpdD5LlPjAiv
Um3uutL0DNVB5SiDKJ6ACONdmNVMY7+A8CJFWymsv5LnXLqSQwk5HOPBLvHqa3ay
kzgeAID2mxWfFSKlp2pjdoc2zn7ICVUZlqePldMqNChBZO+u9LwtalHms1B6v2pM
PdEMOl3uSe+p4O2rIYKnECWs50UjQ0LooWBVY9JweiDutEpBKaSNIiRKq2TWwb2C
hafG9gfna2zum1FVKQtd/jGOTJoXqvwtAPeuwQbc6UBQztpunYN8UxSNMQTVH4u2
hYm3NQaTyuS4Fd33MV2j7ZJ8dAcm0PZbIJxUG7DDQIiC0S5sUflgC81/I9fUlwpr
ZJ2ZAAXLm4OT2+9oaykVKsdUwGOahDWZpvCQADJ0ZBPQMp1KZVW7+uZjmNOp12b6
aY5Cr9lf5cG+eVWETQ5NwCQ8rJQq0l/Zn6pBWLrbsbaI4ErfM2Vdw9z7itPZkQGs
4Z4XvegvWMzaRR9ssSxkJrzR/EAA9XdRzxfYl08Thw8D1hAPw+Wyv+iKspBFtDW3
vYt7zi0FSCH8TpUhOJkDTq5D472ztOSYV0fwjTQeBW/Wewss514lpGDU9rsNlhsY
e97GDA/DE35HgTdccItjewgGcmNp4oHBm0sRVsf8HA/uaPWWPT8gGduVoY4HCKu+
WqhB0vnXWJ1NCPBik5HgesiFjoqXq4ZEBu6tI7vJwfuR8XDOeaJnIiChoQ98XJUX
lXbfEvbvqeUZZs8EsiZpCKkMioMS/9GRqIi2y3spO/IrmWGQY6rHKnc3poyWynx3
Wk4v92o3RYl+9QKRGEQZCmrXwb2VedFfqlsBMBlKp8KT4UVY4CTC/aYjwAhCBfst
li9VyPG4AUagYqmk4i+i1sDbp99egVUUSef/GlE3Sf4EtILSiDaDTRmGdEIROrn7
d0Me3r58T4dWG8XPqRff9JglXk79Jc29/zlCnDis9puMAOYES/M55hBVF33oLEtc
+pL7gA2K71c6Jvr1RzQ4Z15j27A7Z979jXAAVyB6utStC5lJm78idFdIv064zhaR
Jt2upNjV3G1tNNDCWPcagyagIJSZqi1Kt7atYgk/Lq5LQnP5lvreMdIZ8qx7TaR0
gSIzIEV5MjHcE/h1sjO1GMLblNeNuXAQ3wqwUVCMslYhFh0M8MADUS1P1WyGiPgb
RhBnMfKaiU4PlF2icc48Wpikce9AMr37HohfS0IoyxQhCmIrEToi9Lt/3dDVESuJ
qvVtZ3m5ygJiSHCPYbIStkdeMkC+cFMQdyJiz7f0Xxj6YFT7RFfhXqao0WqYL0lm
5UTz2rs6mPtdYelzkGBqWg8XiHdu7Y/hswU06D9dMiR+v/J8+hPbcfeaVH9pYZ3t
KcQw/SAoJDH+1KbMAgxeGDfJ9NkxT4QDU2pE/XkF+KLa3a/aQppO2S78q5M9fgMo
uZKFgOTBhVtRuEpmeJWzswfEJztaScxfkkH1sLRjVKlJvpG0zVCHR3M9OBPzoWP1
nYSdB28PPugkDXW1K11apUHK7k9a3Fl0lJOTOMOUl8spo6xcHBQWfOugh9Wc+3gk
dykhGv0V6pwE87pKovVsLlzoBbrwwFuN/HKxhV+r852DyfxlNPa0HYa5t+KKVaHA
BXCzGEG6kR9cpwWjuhBlnE3iyA2a3RvJgD+g1FizQFGUHuwcJqRwIN9oxDdZHZOb
TOE2qjPQBlW94TYksQ69Ue26LyUXdlOZDsQVs0zo+9eOc9KXYPDL8NmsI+UjtFzM
rks9B6nMgyuy9d2T+bNwm9PadsTKxugTpVIj5tEuE85T3jbHt0HL4c75R1ELNsQ+
gBnIm7X1t69b8Bf6G6XheXr/HHDYE12auQ4Up6r+4Ztaw7XTTBg3AjM5iKFDD8lk
u2G+5d3atrs5zahy1qn/z6cUMGqIs3BTwz/uI/BHxYa3IQQXOfhZZF7kdleG4We+
YLPeqzauWNT1YEgUfoGUZK+E2k/4rcEg4PRsLbkEzRPaKxzFxVjMR+8lIEff59ia
lBujcEF+/M+JVw225DYNZeE5om609uw3mV+MFbxs/AjmdyMyzx91zBF7AQ7m2VHG
nsftmWisap3ohy6Jm7JN6m+yZSSEchH8JOfOt7zk1fukKPnUTT+g0sU1ZPPnlVCy
kDYn7CwUwy2uDRieHEfmpxn/pwKaav8+Yd/sIpPHNI0yUhrUtLR2yEICttnnCz4V
gUCHB2QRQ8xIewNAB4zRL9nM6/t84YWHhaZDukPq2rIXyBJG+Z74wrWGSlIvYlrC
/gvp4p5yxbOGF5o6aQGSYcLzEkQ+HSFf/VKVpZ2SvzAqwAd4hXwtSr5PUbXeXaV/
yKV1RHYT8oncvZ+ksqbc/ml/UDC/SvsEz8YrOcyRr9CvnsYjHVkK+xsmI5mDaKnC
1Cx1/CSNUZ7cTyEOtBLTWdu7EjgXbR77r/vUG8ByvFMQNwzgRsHl02BMXujwM06a
ZGetJO7vE/uJfuw7agOKlBNfPykhKn1z7liyvLkhXmX0h5OCpG/Sqb7HEqgOJSOT
XLO7R7K7jjFbjp9KzWmJ62iRFN+bB9uroRiXMBwsL242c7W9fi1nivfDDGGC4xWY
fbNwD0of/RiNAQFvrBDCXRQZ0wkwe/DAluFUtWH6CbgT8lIPbdmHTomzUwzPubll
zusgQ09xRaIb9F/Cb/DybO7+ThIg9GJqoaQkycnXft5IFdYTZazDT6LR7fxDM9wc
sY+G6nLv4wHUIssFBWkc5TMYJsFy6JSlwEDp6fb2OSDOyIl4J950G9fWGKpj12cm
WLsscNfwdyUqH81pAgBZuAC97J+1hzJZmX8oL6HquMaZL2966CP5kaWFRpuXF9zP
NOt/af6FeOKOWhTplHB2vpqHGHi9Bphrb8dststseF27/10t6oO8Z++5YWdZ2Vs3
S9DHdiM9UsE6JAlnYO1Uc82OJe+Bg3GyNE5D3Af1vMhGEdI+nlIXNeyj6x0omDDL
3TDM1RLbwt17kyMOPGXyfxeGGvNsLohBxu9LFigScB4Lfn+9kQy4EABdtVx7H4Jw
Jsgr/2fhP9w5CypUSlrt+4EHxZvFFrnzR5yzcvNxXF+6dzrM0ujufQtISsc440la
xniaFEUHnyXPZxSVsg/EDG3xD7hnH/moy4NqFE72sMappMiO+RdYWHavzwQbW1WI
rq+rQdR0oiGsKOVfYQpj+aJfrxToP1iExaA4Xt8ZXy0Kum6WI/c4U8ZVxv6WX0Ww
kJjvRxmeKld7Rdb9oE5y3offWUbOjoWPj3cR4Ln4VabuYqYxvHFOeHgIkLKZDpt4
9YLes6bnMP2pIk9zvR8vUluRnEn3730ZUEvKOVUtfIe8oCOLd/aPEeqJS4nkYKW9
8Sf17D5A7LlfAYV3i72MJnm2ypgm3HeD73IWmRT3iNIX61pah0vvOUF2ONdrfqJj
LQWukqIrZaKGQX1sbw1FqT3AlC5AChR0qjsvl+ncqQ6Ycj9ntU59s46oBsu592Pb
7txQYxNQhLIoxjXpCz6WRYrjkUZ+5h0/R/Kb/v3zzdMw5hjYkwtjaLON6fa7v+mW
C4y6xSzxcpNJqDMr/oPtR3oAIciWz4nvd6+gBEKDr82TiEM0RqkmfUp9jEkN0PS7
BvIzfod+CUWYYmuEIcINJnESZ9T/MufPv0+IE7DZagF9htkb0wqtH4DqvdFX4HEj
e7s6Y8JDvtFkxN8VTJRRe/C0x+JehcIt05qQ97/EIpOJDcWLf2c5AnV6ZRpDp6nT
w+6mptlB6vjeWxU9HLqH6lZ46tD2PdrZzXL1zvQaO5HHJ4nBPO1YlMyzrctdx00k
rN1KYgg21Cl54UR1T9WPylG19FvPeayxxz5K+CzUSIcFTR2W2CRhmTkRonfvujNI
Jh4n9iZyd0WqDsJRDwtSE5kRgOT6KjvxKK2vpfIqidh3y+uY9l0Wsz9Yz9W/vgsK
+nqQGTbuR1CHDuWiBKXPPZNnfGRO1z703aIczaK2IG9GsMLNkvXShvEzpqUvvFsx
fmS2ed+5QEdnEu0NpkTMGhSeuO6hjyJKful8vgBZ6vGqzGzLj0F7mRKefOeI3yre
m5bZ9YscYZekYkK6ZYIp6nDfeLF+gaKYzgjc3hsmz7Jdrpw75Oda/uuLlrXAbdHu
o2OxaE62e4H09gQ5mAOJ9d8rPfZXqDzy9agfZnYPwxG88H3q2j5OUQPXBnOCofGR
FbggXJLfVR4cevh7DVqDp6YkHVr0bZgs+KoHRAlowzJvHVlt6S36WJtSSreqRH7j
NP/Xcz20n/nnhMre00KGh7uk89pEvi0STc9vrKYa/DC++NJ/PYW2Y4BsWTMYzQoM
XGIEstW4JJLQmn81H0F7rDao109kJRDeSoEzst02z9E9P99NMkMawmuhPJhd3Esq
em8xTTPJYwX8ML7SJn9s13iaiG95cvpD8CIDEYfAFgmDaXXVhXTkqpsYmIMUfgNg
A35/hhc3lsTaDNDgdWj5p9TZiIyCHOICylicynuyMR7rqlY1zaVsm8CMAkT8n+QO
V+PXjRAh2T0ny+q/BRW6617px31lH3t6nTowKVj17VHJ2ElR4QliiskPk6NHsHs8
TaXbWGg4xVLEM78I/0vR+Us8wlmxeiSccPv24FSousAnrbFHXMlmWDR26OM9qDCW
cSNAoyP3yFfH8v9k1BUtYNilYDDU3Vet+fMylZPApKavx6UCZX9OX1Bj7uySIFMk
lKU1HsixIHSAV+JwOGbAsP5L7gwOqSI8xQORiqaRCEOvILPrBPI4l4RnNWuGqdal
WnuhceJ9hoT8JSTHTm6GABBUNXGukGceHce04wFdeQiUhUE+Dmao3eEqDmI61Xmk
xXQLzeo4vaIQK+OaYqa0AIlzaHinPoQWnVYB+hPhGUNbQygCAXU+vxOIqmI4v9Ae
ZvJiLBi2cpjOJGdgY4G/uKlYXogdWmHe0COjwPfE6egSYPAsLJcEdZH1983NycZw
6HA0nQ2OV/ujOx/QVuH3i+XTJ6D35CxSZVkby9zjPJwvGD/ojrcBIDwY7J2Mjkp4
AlX6oO4EgXk4OP+rFQT4m/nKWP0ZmivwhcCIgtMg7SiVlHQlUJJ8rhNsOYd5gWs0
spTTJ2S0KaOWL9Bc1Mai744NRfUrTkLG8fd0roaus7QpFGu7KJMQsjo/q+3QQtjL
ZvhLLL4ufq7q/8XV/V7dOQNhSFVbjxJ3LFGTM4IaF0zI+k+w2wGDUI/iN7hmVP46
OHzOYEx8KGJhtiN89CJhBdlzvRN8mlt/yn6IIqhh80DohSIuzLHjZ6XEp3zNi6nU
n8FmK8ynh6K2l0HAbFG8UoRTYaTiOm83+0Ae/hAaA+UBIYK5CpWXUMGtryXzH97g
m6j9TgFEJmo+3HdPVWN2Gi9143uw0C97jUc9m3Dq4ROJUeobxgX9OhKPnfFO7LNA
kY21jyfcj6x28r3E4kW+SnYWhxHC0U8vChmWQDdsddxi6ZKYPMeEZZBn62PeFYFh
wN9/Ypa4uQN4HfgLwqSrrEdGKvEOylRKLVD5SZ/4OYDxv8Gg5lJkrVATT/w/HKdM
fOtsE2ayzUfmDoEnpA74SEUEXB4jhK25US2Zrg8BYjcCKc0dpr/Y0sfaQ3ZwmwnW
j//QAgKD7x8iigBOIIeFYEZH4mZ/5p8dKwrXKJyllHn6Uad2Zve7k/SVkSHizsPm
F+8TauKCMXLqovfQC+5E58gfOy4t2T9DgxUJuaMcWSjusZsK21HTfjYK6FQULAH+
DrOK0ZRgoLw+neEOMS+KtISu7DxjSOuZcfw/KrFGVf1RCrCfjH7AC+dfaeJhAoZQ
Z0TDHRM4EOHkn/6F/HcTnREuBzWWKKOlkWOfOSg68emxU34XpBnhXWgp5yBCKWnT
HT29DEDZDmprtXi2uB3Z7A5mO7b5kS6D+0oL+2eZAWODTG8lt6glOQrqTeBhqet8
oqBEVM87B0+J5lzNcjB6+DygmtrFfq1097hzABtYh4R0ucL3IxAgqDerRFfBe1RK
fNvfVUf+hJO5m7z2Vj0lAlIgVr2pgThHW8zrh2vEtPGTTfW3OMaNNpRp75+kvZc0
qq1NkYKF5zvDPOzPp5oIqyGYeGqxdf9LLID+gdZY3FvANl7n4rZQG+Wt9VJH8itf
EVQOZY5wKTzn0xvacbMjvqDSuhxeK9mk5MiOTp8uYROSqbfDBX5QohyQTzet4F5i
/RYiO24dTlVIcD0rjHXsqt5WEkpnoaXhPdeF78/peTjDSZghYWbFoG0XmdGZRj6y
M+i6z+tYI79YLHzsO8YWbGGlI9YdseCYBV7BHFHmznZlU5MFdkOqmLuTSaIdjvb0
fqmGpvJM3D9GzDQ4fThPXQCD71Lg7r9eYxke+8USyv6fPWVY0LIzeZYae6ciYKzU
PULbXBD5kHAUS+0U8Tr2eziJ7OnsL/JeySoFucsJGuM/ZJ0yA9kCYl5jTukotw4F
0BqSdN6jLJoCYcztpBOBn08TpjfDt9fpVggOezr0cZK+L2ucR3wxjG9HwDqiXjoH
KVOm6XHYfbHm3uAwLBeOiCRmMCBpVjRJeJiHG50QQGUgPIySJpuch2IlWyVZuVL6
bKZJDKXKJIcm7VIU457j5gnYae69MMpun9QEYxiCKEGw1Z1+xf8gwhnJ6vuPZtIJ
cq0ziSPK+jpx+4sS/3Xuj5MosCmX97iYJB9l2CH9lzeN0MBNXUny+AJoc1ituf88
UefFWa5KOp87cgzPkavjOILQ81PZkRxNShdT1BWm5St4Sq8/YMuMa3DsIpNnhLV8
VQB8WzZoAARfHlGtEnJ1XJbiteUSk2IH5XhspuzEd+PkW16nfyIe/o9YSIMMsd1Y
325KM8tR1RJBdZ60MO9IkcJ2s95wEXmtGdyCnh7bSh8EbubwOsYB68gyOijcroAI
05LnxFIxe7BQtdiYMBCQEDH24cF+NrOKNLJ3xj8MIc9Qau8fGN1udp9/arIK7DAa
6ZP+Iv2w1EBJB4IUAN7vN/D/uCWnZsi0Gy0l1ZALU48NXXa6nLILXKwqrXJyQ9RX
NmZ37u+f9jK/2YOyNVlsfPS3GnFsD+pbujjyQqZnaRdsfiy5cxySteQBose477Si
+0j4SKCfzsziHjJzG37XOzblMGmTUCboxAegJkZSO4VtrF4zSIFPrBmPfHOG9xk+
sJvwzEASM3mRPN8nv/qMBGZp/3F0YzKQr0cgdZkr5wmIcZH+rrOhQy5IIyC7vjDE
O9YQsIDDbZexQygCxiuaLUyCAKQ5PZfcPCs4yljJ2JNJODVWvFqJdxpNLVINrB34
9rjkKaFCuwjQZLQlR/wXGp/mLJRB8hegQi8hSa+iMgxSL4Jizk4CgUos8Z47Lq5I
Lt4LYQP8XXlkO2A4BL/0E2Bglj4sHTfW+xpegZ4tm4JcdMeyS9ZlkJfO3BEXdfpd
4nFyBQm4XxaIXM7/MGvMQutmpq3HTpvEA0i74u2bAo9nQrM9cNtdiy+g5rpZsSjR
1cPZ1VlZe05BYAAOL5fjmgw4prCr2yIhXeBhsRiTMTzxHR9QyYd6JN4QRCZ27r4C
pK+h0bAqG8ZI4oMnOuc5f2JVV7qxlJRoRYIPHHgUkbu7iDqcO4aD/iYN12h35Hue
UJJP5XmSCCT4aKbk5LXwTpbW8KZ2l/PO1rbhB9ezwjzee2zE5RqV7NkoA03JwMcZ
5eFRoNOudbjNFJ0CIC5ql9Z4HqjiFGhTEPvttMJ4X05UF4CjzK0gtMB5oZF85VEy
5B+EWm80ddKsEI8WLRez7ZsEWy5GOoJsYwQEMdPxYCYwoIb0M1iV6WMDlt4Gq+nP
IIu1a3YaWiFl22giZB8+Ec78BmSK980sakx8p9d6Dyr2JF3XkIedYGU6eEngQvkz
I4TNDWdRpAGqCnhe22ruClC8HoE859pUGGwRUJwHYsTccwWNJlkt4BlQoJBov2xI
LlihantqggsPxP6ZEv32URJ/VETPyd3RGdx77TtnTfYDdSujF6aeySdcsEJzzrZF
dSYWGdFVsLqRgIN/iZtgfmkzF4StxCFPRinvlLupGID4IkSDj6Pv+TlScmUe+HfP
3alzvGD8wSVPZZVROzS7ZtqfIOOcu0YVWioLwK+ZwIbqkSbNtAAKlxzqD57uLXvb
IpWmbw1byfjz94BLKSHApnZId5yFwZCq1BS+14Rgu45h1xV79k9PyzTbdXwRnexm
pwj064TejPKRNaaBCVDwK4+og5HFYy1Fth/xCK1J0jjktIk4WYQJIHaIchdVFcpl
loYu1h/WSumldiGPOUKrZNwbU6kvhpwahlGnB3jTWg97sjyhTJWsk8HSweyhoLf+
B9dcrsgTITNn0lmlWyzj1fgFZOtJ6Pzb5PghJEarm19qHiioHFKGLqGwp9d9DBsf
ENKyZ4wArvANnn5treCAjS9R6L6c8SOPRaQjeJoGOduplQ/VGb916hlW3BGDFioO
sNvjwXNPmpL6Uq9qmU6dyrTdHrcpiMZl42J1UYqXrTHASKuYM5PljNPF1lFzWhd5
ZsqOpadlHwCtNXBpZxGXMG+5DBtJ84ljrlDlkY+QqfouKeKsj3NqeJwK/c3lLvJe
J9HodSDi3CekqaFjUChSm5zBsvHQRByY6Cdr09kYDxoOQu4inIftX0/7hsI/+nj+
DhgStPHAZ+lYJrasOGndfccX3/DuzQQXOFaC/Q7O53zsqknYYwk0xLlsgEphpU1O
4Oh+WeWW0RJO9mKzXOw05Qk62BgERy99zOiWc4puapOqg4TGHucCAmUtFgD+ALSR
NYpfg25yoOnrPS1tvqlQdGdxw/hR2orPbQSVbqPn2vKIk61XLgPXT8sxAdmcWwYT
8KF/wazU8+waVyL53KegBRZJCTFpv9Q+lcXuLQAIrKnoHtxgmIVZrgnW4bEdhcnp
NWS8uUDHyV3aVtso1T0rvCQ1aR2GMmaHbz9zbZXYwqcNvOscFVdxHsaMJ5wRBT3K
ymBnkvwby69mNX/gR9DHlumg1mtm0mDPeVjjgvEh/vyaajCyLLo849BYxQ/fWa6s
7pKKFrHlniMwX2zQcx5T3ICTxUk+w+9yeB54UWrwFhBY8rFA+hnUX1FOmt1VRIdm
luk9pgpIMqebtgXlQpKUnLhUkOTnBOxtFEaUH7d+cM0Tu7OMvhfBCXvRRDeAlBGf
w+04alAkniTUB+AiLTCWzjPmmxRv9/OPrDZAv//HfWzbq89qvbgpjWRBcD/FRLEF
QG/MmBTK+fsRJCvzAvfL57cVIP444Nfvu1o/mNgzoVymvXR3eg8YiwXW4wfpDSMv
5zxY5e9DjpCy2svk3TgDrw7wctUaDQRCjDkOcW6MjcMzcOHZBEyBJMO3axhX/eh9
PM25eEF7Y4Qf+qC4IpjkpOVjGUjqIrEFmDPvUsYRfwsyXe7734YWjsLRnNZsr3I7
2Ljq811Atf7kHo9lcUp/ENQvYqgzYvriIPl0HuPHYupnqsAl0UIPvlTJyoxdzZ/Z
mePSDgFfFMnT+BkCAhBnUAyCvNBxK1ecmCJgg7jZLV1J6mpHRkJFDUPe8qfEJn8Z
zqzHASsciEZOpPbCp/l3sEmryHYESU7KNpMxAetrq6vZ4a4ncqOYRkOIaYfbwDCO
Y9bwV9MnL+U43gPGWobOgZI/eZSu5aJMZbjTPN1dkv8ygX33Nizdcr2FpPRhPGDd
eYwz1JS6ICuYJQwr/j3TZAiSaouwS/XHQyMzsNGB6cTzaip/skCK72GIDofLmaKD
54l4dfGr3Rb37m8OwAO4sguqstKVbyZJN0cbreXZbQ4qZl+FwWBf0eVptBsNP4aT
rhnXzveacPrpBrp1oSmgA4gu4G7HMsU7eRSelLYIz8gqBdiC9UOmFRbeSr7kBPIl
zp9MSWE9r182GDxdWvYd1fNbsnJ9rPvktfTzoV5/PWGE+PZIDgEzydzcm7dhR7J5
Ea7LdtKuxVk3oyp2D/6kCbtbda/Bwc+ggv8iE4v+1+ojcdk1k5dKxpdlSXnYRswW
aeAs5iQjbyBiMp20Ebb16S+Y8GiT20SLtULBcZquXyMk7jGhb7VegoUzERpQYuDS
MkzkeoUWhUj5ebSq7cgTb1pguLrIiGHzxoljzXsDz9pqvrJ2PhcFkYHK+vTgJ2g+
Vl6xo2lbA4fnebUat/r/f2M2vJ7VYxgmyc5s2R4OGO56NZkVT8K4/yXJdJlf3owP
Uoxc6tQOlBgSB51uvFWZZ8DheMSIvvrZioMZh+6ioyNqJwK3flj1Vm51YndhYfeq
V9qIwMHIQfotR40/Wk6Tqam6qMaQYP6UK1jcKqcJTjQD4o5q2CouclUhvI5VxAhR
aAzC53YzI0jmFaq8pRTQGjdtagtF3MP7FyQQJTrdKKrgbfRUlNJZFC06PFMm5lM5
pWpCDr2MPhqgSv0rXXHUpNsPfaW+Ppiz1I4U7x6wHVf8FHJxhdIuLWGnVyQABdki
ZaRWGaLEtqlEk8aHuQreVWradSwOR5mMnATRy1PBRx+lPjIddgU6kMWz21paxVxS
2jmCHpUxs1NxAEyaqO543owL3QmEdlFPHUEt4lWwk+lYXCwAU0Q8iiCZP6ILE4Ho
Kul/04TSiUhCpNIUV1wtofrPBsQ1iyWqklDgPFU+G1zhtCXc9DJRwd1/q1MrRMwL
2ShvecuO15qhtqbeIHHqCWm5EbqpoeXMkSphK5eSufKj6+eJow+Lq0wAqpPVVJ/h
Ud4X2D4W8n/YrAvsZFB2LldfASOEQLqyOHNm9PglJ31qSmdUqZ0nWLh/ADmI9/6V
IlVedSZ4Ukx0pXArawm3HoCV2I6LhbPcwnwB/R3PaCZxI5ywImAwY1QnYTcd+3Ay
X3laxHkYSS0woPis2QNkYmHAua9gHn83RgUpVguIHyL/FYN3hx8s9d4QgrWPuAhD
p3VXXfi9WTs088z0Qp3trK+pJMfqAEr1Sa2VOp4AgZa3Vq0THdTcb0YV/XJ3t/TN
J7mA+pgiPXz6TNuWk9suhFJt4aYF7GZS7hVbg5DrxOHEvNIaGDqvbSUpYGiuFdD/
GjiLy8PuIQv8cWIdcwlUzSIPQfPjIm8lze1CHDjvew+orCzmi/FT10dQaX8QGIyg
8DZpK851GHdWD7xd4cTrTUiAvdHCb5qH/lL9mlttSTvfLxZOTR5D0lGNT/tzyizO
WT1fInFDQ+vYMSrPKW42lZY0ITaWReHoeNyO9VDanI+t3P6zgBekojY1yAm6DxZ8
PWkNeBn2R88uvjsruFey9kFTYiuvAJ6SQCBNk8rt460pT1WL5vCN1y3PJTxynDsS
KltEcSwLG+h24IuY6KjlFhhUFnkLlL/ME0JwKiAIzrhNtI3LUxn6t6E1b95AJnXd
i+BU77IPdUW43YDEXa1ZMAd71/p5JFhjOae1wK8wY0msw+yjt4FDBnnyDMBmQH8r
pPYpR9O0MIQb+qyLh2Rv49aBW2/WAEJhtLmMQ9Xu5PzFm9pwU3WDkS27YpcYi8Kf
6/mpaFzHUe0/2w7cptc2aJMobJ9B0fy6FvAif6eF7DkUwL2bU2zvt+Btv2B5TOum
/NsRQghbOJjtGp94llHSvnh2TyrMLe3H7GZAmT66YMDsLbo+HkA9Wc+QD3EwY2Vl
F9ZUhgbg2IMlzSHsF1zXWuTAMaI3yAmQwEIi/6o4PNa08RqLeypS6PpTsVw3nCz/
nkQv3ijVkDbvjTo6Po/0/x4aCAPQmDFMYo4OL8d8hGWbKDq/DB9E9co7oBnbT5aG
vfKtypODzoTm8WbyYfy85idcDfpfdkrEIFyf90iU24P+/5gwvhUj/W54RGtJpzMt
/InroaLEmXLAvPKXPrSv0iFgNgV72R8xcGU5GbWtAWgAY8YONsysFWrT6teOjT+M
nIO/l56vDOzdrXQnwk+s6BX5F+uxGAg1erX8iHaF4OK/8SHNdMuIwCz0JLw6pV6T
dqU0wNdKOR95Lebpzigp+tordbjKMZXE3TK0sTMilYuJKJKLKdIqqatdAoeY5U7c
IzL4jdUQ8S0aJ+e/4DWKp8e+OqPeomaMs7fxNh7S98bUuceRMrmeyErgJCbfcqy1
keRd5Ssiyr8xk/8P7O1J4wiPX+HRUGn0haeRuMN7WmWuJ+dPozKG02rchkDEXget
K9P9KPFrywoCLB8kvxDq2eBeZSp0Ck3ZRlTMK3PVVDbNTGp2Kr+oJFycLf/BghU6
/HRejTL00lrnTlB7v99rdubKnyZkgGM3lu3tAc1L24Za33F6Z62POUA2Ps27mwIu
NFb4zcLo7Ajykfc446iSARvqEtupGh138W2NAnQ7bszPSxqQX67CMBsnedhmBDSS
0AlDAxWwUiVDOv1Z+sEmUuzzQHf3+e8wwc27iknF0ItDkIa9qjad8h8A5WcdAJ+j
mj+V6Fb5b4ld1MX2F/zD725y49IO4hdEvOXExS0Cx0QCFCcA7GCwd2TUhtQ3bIsn
h3eDPm2kNVmJbWCHV492mgxPyDsGo/KM568lf700jn25X9uyA9gmCHoSD5s7qmnv
q06BzWMaHuAM3Xjss/hOopw7lm7WKyIjJJvbJUtH37zWv+dDse44owgYf4iWPD7h
COPPR3a2rSAUqmO8r8kI0yiCyRLMUc8dt+GXi3ReZbBSNf7FAxmrrMBy6OWpcFHw
j4a12aVm9xPQdVZ5aVolW41+odk/HRMAezBF1JLuFSNTa3sc5R1IoJ0g/pyP4pSe
E1Nyau0khGdr1TnUOFiztzHOfCrclQZlQumJ+R0iGx8JCVkdG+P6/PEcHa0xAqrz
q43zKEl4gCooHflNWp3yVJIJo7CVXqj8HFzUP1Nx6ax4dCExWF+7flmiiH4Aah1a
d9+KFfN5qf7fgR500DxiGZNYW+sOao2woL0dSWk2mpQ02Wjzi/Kp82PQlhzV9v7M
S4LoY8mQOhx3FWApbDgw9YJCQ70zYZOt4pQDYsRi2Oz2EUlC3ukgEh3/vh8+sLFi
ILCAIG6vL/PkD2XLIe9SlNxKwCmhc6zzw4ocBBUx4IB1fEtHyvTLWRO2tTudPSnj
F7o6/zoq7nlFNNTTUTxVHLBrxj5IQIOjwUmbjLJTdAjkcfb0ZH/HQDSvkP3ENwp1
nKNyZz0gmCPy/tprfErZhiMmcqu+iNT+36zeaCFRff1mgjNSWaXU6DCw10X5y9Bv
0zR4sUaoqekevoLrg2PYcIou5jlVzmeWjXpGlBfJctMAlh9AZDPu+XheGqc+crE6
g3aPPmI7fuE2dM8qazctXrBkfawmRQD32AgdHvRskV9a9N+k8O9GevviWA8LH48r
sQuBA1c3sHYK+kuH1Um9DbZ5mSw1FXHu46vI6oDqvaEzeBFIsSCvUrFO1DdX5en0
HcKMUtuXxIUeByDdy1BOD9eekLjlV7CnmtuGAQkT4CQn6bu4pjZm/4gXA9KCM21J
7YsfDh3d85Pr5Y7IaDwMRmLgxafoGbdJYtrUfG/ddq4PSGXeFUQqIsG30xNAoXxL
2yCcguWHDSONtMMxKVLTNGaHMIy6d4bhMjFlM5+tWf1t2u+fbC1quo9B4doD7JN5
UR7A0PNS4O28bf11uhhOkufLLxUD27k/KGT6cdqLSX72xTw+j1sDl4od4qQsn3Q6
Lwejes0N3/1JzPxMSngiWsUbHvFFwOxzb/C4Oefb2bUKjXwjSCfJTgn0i3QfEe85
DJR9HOD3Uk8mWy8UmjINF7Vn3tI6uCgI6A79alrjZuKPElZ6elyKObMxXoo9gvFh
eZYW+wuyktEdRA5TgZ/pM0rgKsqeV91kUvthVMiW2tfz3WZvY1EwBKA9gFqnHWYE
pSvu9nZMraqiv+DPasQMXYc5++l0C2wr5ErM30qRpkgGuhdM0OeFzCeOkHOZY/cS
GVbfepKqEVDsHJ9C3cPMp1A12EO4RrL2Ot5/lsINH8iITnc0qao0Syp9vzOYCAle
q2awdzaKZXEUgWZsaZv5CFYINp4ObCvy2b5apZFBmdhEDlMFwD9WPWl4ZbeGYcXo
jm/wY7HR6dEUwj9a6RGtWZAYj3Y9xGuuf0Iwi4aM11f/JsqYJZ63QBU6VuKXstTa
ydrBw4PGJwywe/NpPmAoaAdEykcCyaqBNoThsMRv4jwRH/uLDDcTQNhTJICj3JTi
uEj4rF3D7nAW/ltd5lgjgjBcwGGTnI5n+I6o8BEF4h4MgW8pCsc9/Oyrp2HJYnlI
Iv4cSZ1ddQ0960APmNCQjC7zu0r0mcB/ZaXV7IcWGxHMV72h+E9xDPwIz5I40IWO
ddd9U7T/o5cAh1dWPLvLmWfwozR6ctrELBtwHkUCd3/AhCwSJe1WN9ikJvfDHNgj
pO2itJ2v8KOHEjsVALjKKKxmyH0hIVIfcv8hC+sFxs9+ud5uMcvWrT7ZQDpDuyml
NLmiYyaHSTEGoaQ29Soklm7tYp+QF+e5uv7E5/4v8x+YWrzntCZ47YfAo79FGG9x
gYESyUr/wx4Ykesz0nrGiXakm0oIO2q6jBOq4CiY1mvkSV+gDJ75Dvn0skMjEvGI
EhBq6wGwwoVopSrYq1j4uRPkbGHwRoOjo8oI89KjcQ8v1RuatRfGh0Gx5Ing/yb4
EAn9Q3vG5Gie9y+748mD3MsCuJV03OXZb1VK1u9DVxjO4AsxmJ9a7yTqYs25GMfo
cUs+eNyS+mZ5JXVulffoXiDS0cfBvYQrKBahm07Nang/Wdyj1Tv/O8SqY9il1YJ8
70xu8xD4Xt9Ze+B0wFiRvk4YXKNkhYw/uAeyacgQRPWTBtXUaRhXyUKYRBuGJ4PA
+tpNnVH+8/oZcS0h+pXkIBgsKjm8ZWJAd+0wLyogYL8z0kPs3+Kxtl7zGLIpEKW3
qQQoYCa7YoRuUQrl42Yp4OIcJd/M5Tw+AaqvZ/CBvY8K96W7+TFVpNXYdidgtYOJ
EsbObmTx0KEF65fCRmqWB/bfhQFHN7bzjm5X3sU61byVXNz7mWU8oGGyyWyIpK3c
LqdoL72YxrM1FV+kHQfMIOD/CTxR3DPzAO2jxNVy7j+2GAV7kVAvAM+uqHoIBgGF
su3hwePgaqF7t/kL3KngaILrGDHkIzRZyVLrDoCqG3nBxIWmmR68RX/m2qdVbBgR
rNo2ouBfSEh/AbipqROBQJvUodrHDgr8uKYyrcDc4M0bCNCCjeWy8+9tKsnn475H
wK4UDgWirBNT4CEutrEWDuhAey0PnWEX137cct3W6NgatVcXfVACzj6OYvsmqr1Z
g0Uv4Siwxf1rLgpUHdqBUUulAbXr7Cx8AQFOBpSIiYz0HE5bLjxXiejmz+9Niu7Z
nwukMVr4uBnfzSRAuYXLGVpRYAQIWTygbrv24xBdF2dZOrYc4aex3aKLoCt93P57
Ez8CqiPaPnbWTefF+9rVat33IcyO+zVoAhfLTZ8bTBsb8Xhis4DirjF/YCaB9LaR
PZ5Ndw/kpnyC1qTsEgTz9A3h/Z46Oy84Y7PgKmcCh7RXwTn1wlsyAGGF9NyZAuiG
p2sQtHsLKU+ZzuXPl9HjE+hDwn0lI2OrOBBthBHAOtMYHXHvZ0NRV2C4VT1zoX9s
wt45yIRoYwCgTuCr42609CU7G0qf3QPI6b818ftFjqI75Ez6YpTc93Xw0vh0pl2P
2w0z+B/GqEB5bEEj7YmuavQVrcJyAbfU/mMPAGYhDh8fnIitwXg27ZtkypxDuvsG
axXF/mTBbu2hcewDVt36do2zFZ6sVOaqJJjR5DX1vE1H3MSCX8BWzcg4TJ/LQ9r9
OqL9Vp/lazGKOFIaaj81keBsB2ZZfJvjmankCwILuDqXPQIwdNf1R9COnLhPMdFy
4M5pCb8vnZiTDDcFaIVsSpHPajpeLWhktakHrwi6PJ8ZxOQzVd8npqhdX7amm6IF
VI2dp/+6WPl9XzSb5RSlndxsIzyhSX5AF7eYiGMa659endZqfjACQkdfbFZzsDWq
IwU7soIeK34S6P+a2qzDOyjeZqJbetB17MAT7LNZA9mO2rSbUWYil5BX8d87cF6N
KsXNqpcNkUpTYY/m3MikJJ5iWy6jo/I9e96kweidgPFZZglhD5NsaWWIrEjbV4wZ
+gIaaTRRVVOLQWo3HKuzlc4VTKvxvVvVQRivSmAGzT14O9ZL0M/w6dzQMoTnvUP6
71FxIbqw2n1CGV/soGZL/3NGtz+dO+RC4UcCGShU6f/hlppLhwRCBAKSKK1wt3hO
q42B7PomEE2GCo8LkFiz2r9IOKIuxSBwB17a9d6110kcewUM2yjG7YMbouKKU/TF
cJeezHPHLIySe1VhLm+aa8ucvGOwY4bRBKaI71+3VpjOcsrh6clmFjqpM/OUaouC
gUgqVgMNGaJ8yV3Sfcu8aGD6f+UDQMyg7sUr5hmXJ1ksJt/LTvkp8IY0kvfVfE+H
g+Wx9tgwd56Pp2KDXGW1czQRN7YfBykQikKoazch9KwOCRRdqnIGJPz5cWt6CfAZ
Vb3F5Ft/4nFLNoXXktU2kiZhKeMyp3XInkt5ccuY6A95qm58/su7BXDG35yfeRlJ
GMoF7ScQS01dOC2sL2Y6p6e2ggrQYNZU8ZUekLFmySdjn+f+bj7qJRfauiHPj++q
WPsBav6xlUUgNvgphKKIjM6jMv2L6yZKfQzCW7CrJa1+6kbLzcOntaQqjKSOURhp
pl1PVIbdnhSVtpZ74d+rLSgamJ8JxUE6uaR4XQAbQ4Cjk7JdsC+rh/CiwBXjBHVi
sCXSvJAzvw7HMwV0OMYxyCgvaRLbfgT2MX1lYUX0ZPEZ1iqEBuEh9iNGjylZLc9d
/QdnNqgf1lzEwX4y0XjTr9LrBNxqG3SfSk5NgkD0AtmJRERkwinhblEsXEAL9H/j
YkUn13fj+xTbL6hR4l0SuyJRzjBo8NMKRpFypsvpw0oy4O/zUpmLvwR0DLbEj9CC
M6euwy4Us2TeTL0yUZ7ZfhWJLO10G87tE6GrtNdbu+Wu/a8+4fEsjXKXS4RfVYST
f1FSVwKg8hf+9xXojdv5EVLXosKxETQjputdsyy5KHTGnQjWk580NT8CbWGZHBTS
iNAOL490LbM+uX2W72WIA6gHwN6cIVDyFN4e9w79/YiiwyBbtZ9n1qnJRNz+Z0D/
L5cCNILK+QBeUR54Eyz+LGZT3hSMtRxRJVGFUZLYaS7VFGXyU0+1jnJA+BFR9UGL
YugjopdXQqAricW3d2AN0Ss75/NC64R48io+tgywo2+zuqkuEUGPZNgo0DQZWEea
0o2+Suh5deHGAkcaRq+d55DDKv4FhmxNQsPJhcNNrnk3wjsFVPfRX+8aYveLFUud
A6uDJuK0b0z5mVaym7zu8RUvsvgVtiba6rw8tLnPL/O4sQyE0YdVMIHVoPInY7l6
Zg+9OvyOLTlShEV6Ztd5Y8ny/D3IDpW5zYWkbWAH3vF3Y+3ermCgGYQS6stcCmQK
9BeuU0+HCCsWcYvzrSljBgMBzv/+5v6/S8K/iqisR6ygmTNzBuKdbnsnx+wRrOWn
NpJhiBmJCxpnxvZq2UtwB0Rgy0+G41bWjC7FqDgU6GOVkSvCzcnUdUD06/hAygC5
fgsV56vvASevjih0gCGgHDDH+rR/Vvm/4wHHfxeEtY4p58nx7g/Eg8jxkrUGonhc
TKQUh8E+52ZZw4pl4VgiqXKJ1sLQpTIaB3tFWqMXOMeK3phIhPHlDdrVFJhKh9pF
zr5KElFo2YWUp8PVG9tNnZjOlG8N45Sou5urFPWr9ZIBJU02w8nfAmLaVRTtBvBy
FDbK/m+Ahb6EifpJtSSKpW7cR2GsF0+S7gRuyxbG7+zKptOt4UtOE9gKyXytkvZG
jNTyL8MRGZ5eN9YvrCEWuV5czzj3+AdZ5EmQjMY8gj1lsV63/jO856U/x3dxhCE1
tJoNET3unw7tOarcKDMLV4bQViBIIbaghM+zIKgvO6833OGChUCehf6mR+NSEzrC
m3BLhiqmQTJJBbswnPQd4F5bgq2yToZHbEIgNBgBWkrnIKGyerCHGYsLV2331ZqI
g4o4IvmT7+pWwMccLL31FtPqFMY8rtpLyQNKzl3lh/lpHzuRfnAGqAulTLbPD3TZ
wsLfkgeyZIPiTDbC29YUSE/wHJBv/ihS+kPnKiR9WLRFE2hbDvvbOAVbjJBj1PRx
TUUSpBbJdcmS9/daInLP1TnDfxj7mdCdwDdUI8VcbVJ4ickksCdyCl+i/+dO9xB9
Vo/m5wZxjo9p5szClET+1mX5ly6ig51xNxTzeZJRWlRn1lpnxJFdWOXFiUJlWFHy
0STR2EWjbob55kymSDvcmT4SaEnl9d5OKUdYF0tgL5j4LKR27OKkKvIIwA1A+Zkg
2daRIp4h5vXBUcwAFxWs0IDMn68mWXwOj7reOVScpJ+RyaZuYTpMK513uqxXbKcU
0+aPW1y2k4wz6LYQwpUwgjuGyNUbY0F++6EhmfdG8wBksYmRDkIGr4usjTf5RDpU
HHmVK2WWg5PlcSKCF52inHULY5t+cuStReTAf6TMoxpADQZBRK5yJNusVPf3uhTe
3O52LkWWmeGasmwdt7QilBJeqr9DJmue32GEYJ65ZOTVDbO1JeGHAWfXRNPHVb+/
OMR10oC3FoNhiJrCRIMwgqkVSL3VEoCMvW1In7AnL8LmlgQgFcNgiudMSe5UoN/T
N+8d7O0S/OM07ydlXRyaBy5hg8j8T1Zpr0b6XfdTPnswGQx9In7btLqTxjoPOaX5
8WOF1OjSLxzFBH2prZUsFiEbhsOnUauQfvbc0foKzENGZHqgrhjmKVIRL2LxOBXS
lR6WTYijbWyYbixS0r0eVCGQO8za6HsrZ8k2zptpeA+XPlCaI2tQtnztpyi5Ibbm
olT/mMo0Mvak90pTrg8exktBbEY+5iGYkwr4Y4qgsn2jCYXBSgpjnCbwSLi6mGFC
qcPB6qXRuX/I815zdrX+PQWm4CdYesFdspRanc9S9Eg0PWcvbHxU45UN0mmTXh+Y
XQHqGPcCJ4NEzmqKkE3MxlEh7Cr4RMuDHPOAMZaoW0wC0wgqCrebpbEb3i7+U3wC
REBpUrapZjC3xVBRjQW4DlwbP1QTQotSkolQF03yQOxpzIcoVeMVKvxWYrRxWtqy
EqvlfFoI0hxPEoGS3plUO+q2SClK9SefyWGSjvFXL69AdqtdrIDbHsBNoPHtQksm
WaPhthkE5J51GDaSedvWtoy/G4MnG8CJHYBrGQpK5mX8ZD1feAqIKAuns30+z2T6
8G4ZLFdnmyCCX6AhuR+ltbj2WjKhUp6jiFa9e4F7VyPN0H1DxnLnuxnJYzVKIqwM
X6YpDUrOGKxfkfOUxHDQ/a59yNKvBsD5vH2SWEmqDQrrC6VBtr7NF2ICxrQPSUqF
KCCiOm/2uhVIISKiseknCIfPl16t+d7igi5sxmaLEpCRv6lH1d8YPohi7viwjTWc
eNbVi4SpN+jWOSl04M1msjAmP7jxxkCAYGVKxy+M4JTu9diEgpswtFyz3sFfIrJh
wTtrX3sIZ68dV+1u/ZsnBAA+zXFYbkQoDxSSIoiajhU0fkZTqKLOUpHaGcnbA8y0
yqDHkAoucNT7EJ10Z3JtHY4pe1LdaPhfa8YvLCn5Y6hfXpWYke6u1VsrV/IkMrbm
xNlbJ4eONU4LdzM+D/OHPXan8RgpL9LO1hr03zASDjB8JgFx8q31uqHqcVApoVV4
iIKazBxMzeCKceiGMTWQmAfXuLIFkyNJg/C8miBsazNwVouWKYyQRnRmYt4j8w+h
B3xzghb4D1UT+QT3336SYTlNy1rlwwgnooj8Uw9TRVVT6GRTdsUeYIvQNro9ixIq
Vbj9Magd4SdnURuTu/Jzr/i9NNRqtn9O00Q3eX8ZMs63CVu2t7M+aigWidi4F702
NUrPDYgD3TZR/YBIt2SK8eigV9GR78oIC92xE1xa0F2p4DeDyJJs1bbf4T0mL1RB
+nMt3t4jKkS1idtmNDA4jBalu3Uqrm+opuYw9n8N+dLLXPDT1i/B57Kt1nBF0wQb
fYwOCaj70bB/0a4M+kjqbgucZP0xgRBMIJ6kcwx0dO8AZjitriA79LgIW/4CyFq4
E+ONJq+BHCKVBMnfvG6w4GiMLHLoKe5QI7cWvObT/uipPQSQJzEYFLI/S/f9O2Ax
WSxdgzzwpOauYOoLFIjJ9NVWH3peEktIQWIFSjp2bZjaqyRoB2dNTZA94j2lZMwS
enN53CPZCfJF+zckKU1o5k3HXvOtlsyaP9kxtHnB50+wR1K/R1vAtuC2hnXksZyP
kBsQVxXl0F00uzjU2YuMeefdOf1aA0MyDQIGULR8maF5djVeFNiHe1+dl6FSSPky
+MzBzrvBmH5NDq6m2zI5tEKeXX4ePoM9xrlKC5BNfT6EY4SpSLYNEdaNfAJKNQnZ
A4Zssj/v0NXNj2NoVLgt8MkXhXacWB3B/2jhLqWu9BtPsq9m1qcjCLt9HRcSD19E
OA7Ytnrkr3T/EZTLMicZfAG6j5SSNaFkvPXGRbL40SDWZIjwiStEUtJVvSNopPPZ
J4MdFK6HvY1sQH9bDOapDciRH2M8O8xXUNKlzucdGcl+QStt/jhcoEHlrQb92P4t
SpWomQg/jfV04o0VB+kWmfEF3r2Bk07suxpfRKkfZrjWaBz/VWebuFLYMUurJx+w
0mWGrVDO5/5vbRDaoX5ntEo5aQaK4EOt8+ccpwU89T2IwK4lx6mQNF3Zav2dJ5h0
7ODP64rDmcaHNGUYPxqdezXKfomTp30wM3aC7UjOInuJnFqUyDvGTgmqAL5WQGwi
RmI8U7YCF5MZvECERN+uK1s/Czz0FPtDZ3WMwUZ1qQ9KKpcPAKY2wrhnXM5hgLa+
xF3YyrVZ4OaXcDZLtq3kug/1HKfbaGE5w6n2kXMjLpHx4mtFPkSNIB95WSDQO8yT
rrTYWnZgJJPGaWptxknZ40F8Oms2vY/cUYF+FlIUeBrDOMYtHrm6gtle14pie3HV
99Ep9I1NKGVea0WygvrpQNTXQtT7ogVEHnwnzvmgCh/sqYoU96bbYhNc6lpmh7Ec
H+uXQfU/VWT54VEEaiRvBkg9pW6QlV5gVie440TALSEdfi/g6aXFpdL5rDMfEFxw
jewfcaQdQxGiiZFC4UbVKrHh1sQt2ZlkBcN3xiP83tq0dDuq1Mnk4v/VpP/jfxXk
f5RiSL2PngsD8Hk27M4Bv/iYACu+zXZREs2EBlKQxa7mPSQM1dgDqHnLavuH/8hG
1d2szQwMWlC3BF1e4An2zA5piaafEWQNmCAWjtN3MWCm9bI6KnURPSx7tefQOZ+P
qXlO9QU5KloxUvN3BjJSbZE3BAniStVbGL+/lEYPeC8sQiURE+mBeQOkVHn9yeaa
o6KGK3jBVur35RlIIskT0v9gjfmu3pTn7ri91Pm1+ddmB72UmKDSLv9F/M45HRW3
qAo5Qm2+kMrGqAkEMjpCChbEHGx9kwr9xU1B+1uZodxe6vJEvNaWhbJdaX0HcxFR
E36g+UCa8jatsCi9rc54IOsnsi/1nN50Ayqgq/z0HElUgsR1snQB/dIBXoTF9uee
MorXOVXbU1xxBokEE4R+i9KJZh8VFkGzUYDIJaNFzBQoxDGcw2vFZmtt77AW3snK
48OK197QBE7bMHyDrtXVmzrYKLeiYhJepC0ToOjid/JoMOcWoIESs9hItsKIE2W/
TgwcEZ6W9E75wLIPJYhsPguFOhdmK/8kHNy4bMIZS0lDKwzr8qxDHZqTtZeOb/kD
+BgdW6gN9YA3od72iHPkDlEIFKGirJCI2gSVPSBFdfVTlpTGftP75rly+9qS1FSZ
1UZtkbyk6fnj29oboz2tQaxppklpAzTZ9IWYXXk+LEmh5vKIMHvvYjIeWZTAbVWU
nFWYl+jHmyB6/DTo3z/6dKcDGxukwXv/yh2kj0Z7JEi7xJV06poxXm612hs/DIM+
o5kSRITNTLhrIFm70gLj7f9fd2npbClmPzPUL/6uEcW97wm26NoWsNOynGvm1MUM
1CnWkAVNkVqHAUEJXc6UzHrINIQhazKZjIi8A/ALAfIh8/8P5PFXjdvgDnEC6bPc
g7GBO88bVtcAjHbtQO7DJASTpxKBlfWm37/i0KyT/DxD9toFKbiviYKh2J6lVXsR
ZafPwx76Dm+ZDtCM2tk2lMNjvP0jd/z+dTSv8fQ3eQIramSYyM9JyG0xlzYBGvMW
IYVuPV+6YoQGgjTem5r30MQLNataCQ1kButzkQjmaaGpJzB+xXB83tABGo1x/dJL
8htnv6u4DJgcuOk23xiGvhyIvy8vFmE8s2Kt4yywQeydH5AfHmzuCkDGH+MN+baN
Sv2B+ZH2yeKt/+RVu9FMytavCH5KrFEBKmXv8MBq0sPunBRz8SE7QtKSWsyPZPFB
CWCJUN5hhnhke3fCJoOuqV1Svm3e3K1sObJzVx98eeHMP8B5NR5VTgneif5//+EC
KhUy5iwQrxL7UXbPXkMb//nrLi/6J5OBmQRamgBOXdmYU8Z1uaWK4j5ny3mPa9N6
0BO8IhsHibJxYYyuyW9gdSNoMQSjIBwYSnEaRVh530AOJ/Gs74mmrlbSBPfjt9CU
d0eX4gWCiRci2/gNkKhuF4oRDeE0+L4msnk6Imh/SSGagwXZkrwVvtJ2YQBGHKCm
xtQDW8P8gwdZc9HRdT8rAWMp9OPhPG33B+AzPevPqMxdIh+2DtwKDtnbkyMU0DKH
K4PRM/qshZvqFchttyr0J3OzWZe47U6lT5WZ0zMAyNBxxMwXlYpMZwcMlxX2tt1G
ZCm9IecSERmLJZ06QCEErYp26Io2acNR+RkU1RsyKG3IgPnK1iYldVrcznUg3b9I
13WZqlDOiSRWjscZpyC6xcPnSpzvMoXOOfFMZTfrOh8WgmWOjb4lim4RQWOpyzso
4jAnuqFxOJE6jEMjvXAtk4HIfN5tGxjOLZ+Ssl5xDYMfwWx3oW092LzIyYme4W5M
md0CgfxbIE2dEwmPwLn9q7Eqf1xwsUYTxhiFT7JFVI85nx6/elRC45/VNNyvaNy2
CWKMZk7dSL2cFfnfE1uLLxZDHhTMu/KO3++mUB15IJXDQ9bFp0x9pMgFsXTW3Mn/
PBNS8ykYW3bmbEu+mnMleh9yaXOH6gfNLHhjaZrD8GGt2TvPqM5Wi7Srr11U42ga
AHr6n36ehH3WXN6gHErfJ6+onIXoV5anXYCalDvX596ZNRWrmcR6+sOhDHNKDw2y
ddzK+SR4FytmgYnYluIHCIROJTCMl+1WtB//+G4Wley0hJm8zcbaPkrRw9hNHSyk
gzW3C7Owwf7ep1b9eStwm8Jt5lkM1eJbmRcpx0AmyUYarcW/5mpH3YZQKnvayt2O
72ZSsYNs05e0xOwpZd//oFcA1pGCZzGhO4A1x3z/ktpp8OajRLMTCGLvQAAeDXhK
gkdisqCoBv4JLux2xyC5LjV/Z41awdBzrhkU0w5tLWnhO0+3iD3Z8x2AVX/51jBQ
CrgR4zyDHmBXpnO0f3CWFElqvihB0INtTmsYyq/f93Xmo6sfiydgNNEpYyejfc0S
rgp4fHrQ/rdoV3qZuT0P5dfhbNBcbz7G9Zo9Y3YfuAM63tJA3Rn5C+2ZU/1aqdOw
OvltXPPeAYrHhYDMg8ZdcKH1QMAL/GQ/bczon/VtHtEjZmSnHC42omspfJiXMHEH
u+eNobFK51DDKrNuD0yfEffp4J8CBsjsUwHkCgJ+PVE7gQF8xCare53to+FlMx/2
62fDzfLUsaztI9cV6k70Pi7PllhhA09584yHp/T9vVs5jeNQuhf1GQVLnj+/ckbK
L8azpM5/65gDZiIuplkeBnVV9Xn1JZjBSygG7LC7ifVfoK+ilqBPVw6R+gbY8XC0
Z2nzvuImxQMwe5jyNE6nwsgEMUPfL7P4FfFyR2Mvl5x14iFAI1fN7yIh49AhxpxH
1n/PTr7ohO/pIGoribyjVAl1lj1ddEZX3BwHLk2e0o2/FGMpc6H5CSAZsudAQtYA
1sDx8tAFsyG8269MMobpmXD2Zogb2YnB9ils2+upUUSiuiS4puTJwbIkA89XEeCx
ABKrDxJa2kj/vxumR+kcuzo2A6/hRXR/NXE8Rh886ebCBGAdD4VA9OSreuUrj3EC
sQwPaY3PZRIUfDuWpLw0ZcfxbGFlisCxO+d8kvD/8rxKXkT5dwFjwpskGyjzl1U/
XIwhfwbci6/FEZOrVljOqPwDZgZ14USMLkM9AIu+aOUsKX4rC8x8eVL1IQXv0OVO
4CJblaEmGeSwl9wJVViMN3Y8y6rG5y3wWVXGEoeuKy3sP57clRz3vTCpoKclb0gN
ffCIyczecrPEo4j+ZMMA7xAaSWvQZudAomS/+9h8FDcdSwywkvkUDqmpEVX53e4K
eu99VlPFGOO0O43GEuP4Gwpe5Eyqteh1XAu3ZOZSo93Bav+h+0G/cWChkJn5grHR
i/VmTGyIL14f9S/BFC/cCoNSQuwCaoPkOmFmH/lMQlFm3fIcG9ju12L82laj3NaV
PrABvGhnJ/5UZmJN+D4+LIhN8AthA9qeVvRLjsxoUFS281ippsNLndl3egrGNA0p
/UqygHn17xGTTEWiidiL3pP4Jbzyu99/qUo6k+36Tfy9rMth0+XbQzyKqX8MUPKF
OEEClRyM3hs+l17Gjp2su4C8qbGn4W83F/u6SnnVE5RRix2UyecoqtOmNC8fn4PO
K1G/cAyDRP2hWKxa1OwfF5l/wFpAzMpuZoCCe42OhFor0i88G6sTETS6qFhhInpp
uNPqOacki8Rpxb7kgCNRHPV+cxzB/y+fFviQLkxpVtyB2NvL9ZpXgKssu14pb6sf
zMWq1VZVrBbH79XjpdaNDkxK9sFtAwguN8Cg4pUvqbPU/6rmaniZKeZlqKv8TOfz
RAQwJRvmiupYkn0HVQzxk5/c+VEyrQ3Wo6sWCgm36bZ7DqrorhFLFRHJjRUnxdLP
iJvhNTGz2JcoA5ceJWbosOMejd4w+usl8E5zON4vq39FwfCqFgL8TtYAtuQrNR5M
2Ik9+P5qyqY/REMAw8UqN/hVElraglLfIZUaQRt9Pry/uPmZjcgJ6YgPSOAbQirB
m2We5KAAU0H9FHMruOnJeq4ZZadBYmQmPnW80ZpxHBMkflLEw/1scobtPT8cqnem
PNdD0uhygkUR89LhWTa8P+cMbk9NPZlh1LZQLR7zaE2mVPbrjYI/trUtDAFtGQkB
eYxBEEmECoArnoQLJYv/LWS6TT8LFXqqya4ikSVCX0C0TDVrwWpnzJHoB1piwuqY
eZEQBSKv6mOP4KCbEq1wX2S286WDSAiPUdqvsUBXz8lEOjnz+TKbqW1gsktlHiMM
3sRSHqWZZwhFpoBYwAsabYEyNWrQAg/3UASIwAqdJjVC0p6XHdS4IO52/j/Z7FyP
OAZMa/fbTZClqlVGhFCqtlsnYoznxkDMlcdUGc8gibO+0AB+UmdnmNolIeh/E+XJ
djMob6z5qcooADQZrIltB1d+dNKY78iWdl8uxjE7pfn09gqR6J21mAt7PPjH85zo
rB28q0nPSm1rNFksG+CAYHhQ1P2oz/4ECXgodjiptRKdbil1alhUCZh3dwW+nR+Q
UTPzUg2eM+pokwZZnu+RZFnbahhyYGI5T+LOH/mxri6JF9/gza/dn6+wvFdAPhev
KTCeNNkKWvcM82cabykLSvTsTvjlBmD94dYy8YXqyjuwANJCxsiHYvWnjA8WW8BB
nHCiMzusrJUxSZV3U1NF5L9QTGTfMiWLoRaaElOqTCnMkzKZi4DAGCFPriS70y4i
d69sVZ4t080IP8zDjx8yCmt0Hlh8oOE4epTMbIICWBNQh6DN3Vcp6EKIlyen/L47
KBFquVV7WyrDSNtUcFXspBcfCPidu7j7wL5Y1zFipZlLhIKUQlZERrl/QwG2maZf
O3ArAzgXZqnkJB311xyXfqVuDcLRgnHWi7HXcnOyiDMMJlHg/pEnnRd/UUC4bOZ6
cf+iYmwY81zBFK8PekictJdkQmmZWz+w8vowZL4XES/KTchgLEbNeFhHlEABu/WU
HF8jLhq2yooMLvz0E0KHPQVlkaQgSHn9Xt1LKFCe+wNjnamT1WA6hKXIN2vs1Awl
7MESO6YBtec2BoXZDDHpwpnarrZ+gyfE54J23FvZoQp9K+yrUT9eTlDFwRyVDVUP
En3DMgqikFQG+HUyEBWk34dniicndh28ewM6tqpGJKuT0gNtYpbD+X5febi7tOeL
OVPqypj94cn9UbjgtZpxDHOGO/8CL+5uOsRivY+fUi2uhmogD6Qi/BI0xKXdGeN+
WNslck4xdXv8h5V1GgxSDA8ZWuJsafMGJW99yo+YDwYIKokV50yiozbBjsUGAf7u
TbY7JaUGN6GUCke63It1jJnFWt9QNdV+3eNZd4vWpWDwVVhwONAL3mZwWGqYUI3Z
QH6ymGUqmIH10hqAw8AysboiJAcxIezhiwNZHpkZjZ3rf0ADGUZh514G6JxfhNPT
RII3tkrhgx+8UuME/8cCVFqSpffQUmK3T0IIXKsdyEBTVhu168ADf4EUM6k8bcnh
mXookAImvI0SIZPEWY7vGOHGhwWbMCtoHycaVSzQZrPwocuTrZTnaiWeBIl7X5z+
+piCHelxAFw8RaDtL11QdasCFm7LnpAwmR2qou+fYJCke/2Hf0bHVxSaXp6OjbZk
QNSQpK+rEHdm77QPSRhwqtL8Q151RFSGAnT6X32L/rHpFpRMNeLVcXal2N41T3F+
hdxwEXqz+EX7RCnMWGzinJSYKMz0jeOi2LNyiR31CQGK0FOMYWlNfr+XCipkwIlF
W8u+ZDdN0gIYucnmcY3Z3CTsQHGy0vl0eKgxlM8p1tK9MFZZbfWVwrZ0nIHXBWm7
M8o7TVEAXCCXyOEgARsIpjUpwSo/H4tDat8EdaNul8KKL8i/6SGiwWwu6A2RbNuR
HSpllZbq+0Mjakn32vpFGPDgxDTggzia/8P/m2Fze9uGLQFOurVI6JAD03fIrvQj
sYe/C9DaWDi1QEj1d8YN1jmjjikwWPIQzHjDnYy2uYskdAloWNmvxUy5LnaZVeNe
6ql0B1oFJ/+FtQpyC4ee33rHiCmQpuq1bUtS8dym4u5V/LubZ9R6aK6gRwg5bwbm
JUSqs1MK70n2vl+MgvacwUk+ZdfZj5gFFNASpbzuWGmRN/7tFJGP5xXL+Vt4Km/Y
vRlayesN2fyN1XFEG0FiZYSzRRXragOXW6U26nKhweYG3Ld2Y+R4s2sdAXXnXxje
gOhsQA9n3Dxt8owIJNxqo1FbNAqDAzhtC6esl3zSG955iNzhQZMUa6jKXhdPa09g
nnWMCJ2I9BJDXLj+aDMG7BP5266ebtA/TTY9jYoAJRSGdWaOdO5ZzbDFnmY1GZpy
3Oy29xR+IVv4aj+2uENCFU6p9l0bAzYOrSGXRhGpKbB3k80XAb/iMdadhF7+d2Uw
35Uv57WSqHsLoBbXU56YT15MxdxX+4BSbXgtmr4rcgBgVTR97dDr9/lqsyitgQ1B
2FAKvThYfn02J5qoUnfmtlW6LIQggcdMYwwLaL4ZrXztMX+3C/XgzAKyYdQHcByO
0wns1KH7wiBo3bAswxf+/C04iXbpgzp7ZnB7OdYyNh+M01WvpaVy6RDxE/BiamEU
TZzTaApGvHLgN+iS5TIJXY6NRujqdrBWgSFJkFbGAnjAOWKbhH+qJr7bBlZ0O0kQ
1DAZmFsQ47plHt8G9MBfgU6zWEQ45bnSQkBP+qUAM3Cp3BJNKbdEYc9rmBNgCqmz
smdnE5FcNdZ7R0SPIMCu8/CMBEEbFrY/wak/HpOzcxrBrwFRo0wE8zh6c3uAWRYG
EZd6HSf520yZI4VQTPv0x1J257gOSIrkTBiD1tUDx57l0wIt3+o5rFgasUeh36eJ
BLP/khU463mDKluYc0yWJdtVT223dtKl9d3c48hIDN9OgMLscbK36I6xxTa1+7Px
MoetziN9h3FS1OHmBhwuJKN7yEO1vhqNtNW6oQLgZLBV/8lPgiKWzY9uNeEttpnw
rsXA2PHEOSWutY5zstLwstoOEmeqxfCKdMjJXTuXxHYA3UxqZPKKiF4MVadUN3R2
+vnwAYMYpJ81UlirF64M9mI9ayDEMcK/tTbN5OpaNT3vjQlhrcGBvdjCp+Gzfwl5
9DmU+/AKI0e45nZh342LuJJc7vEs4I/NCnEY2G3R6j8VjCtNaaA+WiAScM46Bua+
Dn/9R8nzkMEA6/FUSRFFu1TZaJAmwsNAvFltcTpu8pVHHjIvn3JHoXUkdWw6iJNn
Imki2PSh0HwMWkMwsHvP3ew9+UVI0gwhvTr1HzcKwm0tWHvB6AwfWSrVsFeK9V2Q
1KUwrj08TuKW8EzOXRUuQ5Fc9W41GWCiGpN3xC94eZiNsbCGdW+UjcxAlYy+Mygl
4b1T1HuGqf4uooLZRCQnkixu22KCFL7v+/PIekQ1u7u7u2F0sADV/IlZspod2gAT
NbZ19HASru6Gg+BT1Q6D8f9jmU/73RYO0FlngBczuPhR9JQ/9tm7E642rC97QTe2
AD6TCJn/yEjC7nEAJUyADlyplpKA0gSo0KZ5hLI0m4qSoGYsnbSqtDt/ECgiYAnx
Asm96b2asUCCCOjqeEXXRGyGYm8qGrhmVzY7XqcobNta64lRSr+fhjp1INf+cqzj
BDzGOF9m+uEj5dlzMb8MO5E2AxNo2hpHOkx8morqDcCXMn/wMSD6TIguZM/wfVZs
d4znadQFbo+g1QwVvn5ov5EHZNTPUpaA/AAasURsgyT6krSh8N7VTXXgPrBIiHRL
9mN8yyT2DPG90/TRawzcaSsvZYBov6WDfTUX5mVGwCwXe3CiSkPuhYBwDK8itLcI
1lEQkAQS1ZMec62fNoZQSDWiMSy8MMgpPvxxN40F7HnoeSGCYKc+EM7M16LQeFC1
T14NBXFaqst9DI0ZPxM0if5iR05rwXMvVyXrRGJwJxu/OoZ0zugiP78vgpSZEFyd
/htLzHtR0SU6J+g7fjenYreJ/hbdwrtudOoaNWoZO9Wv7Roh0vPCJCOx5swKE6D7
wF/Fwz1JTIxpcJvK7M9x2SUPrNdJUb251GV6Yz5hqwmdZ1+811ZuE+vtZd+G+qu3
CAMHqnQ9cq8rys5D0jmmZbOj1nmF+eiHF0A9Qkrz9fC6QLZYiufp78NiqQV3iL+L
HcWW4vaKbSjWfXVEsidiLICKAPR7VOiwxQw52wNUBLU8MyHq7yXJy0/S+4iy7Ugd
abxwdMz5H1CYmloJxoEMcOFjYt+RFH4PBigGQ0eYL5lyIVeXQ2jXHq+pMftLF5Qj
qO6E8nFBdCfx7aE1NlQVthM4NRJuOtDK8cQ+CXoxzT3P8svhLDjbPgocXkTbKTdC
yqFf3bBEi8S4jQGEa+VblYCCCdNTfiukD+oCsklXmsDH/ZhdfO9MowHlfQUAMur1
Qnu/+8RApAsedt3YX6YDozQNnoy++p4FSaoP6nzuptIj221oNi3eJ9PsjRbkb+xT
UylvCz3synRNc8cD+XOt2JVxs1sp+SVFzz0zlKEySaJxF3aabczCDJ6BOkCryLjR
VjrKa3EzpiqzQNtU37h4F9/h3NcKOJNBsPIT8KCSyFpagPJomwEgc1GWBCTOFNor
xb8nezyjCckxNNrXIoXAHb3kHHkf6aObmYuvqFCqvouvpes40HXJBvzylKJEWUyh
hpZKoP3P5hn0xyua22zMO7rHGtccmgptI8EvwuHDE1cyIw12N5tezbZzI+zXgFGi
eM2VZBIAuVcy1j39zwslMHOOiub4D0iqALLh3jAyRVFy9CSkJPFiVo5TW48j2ny7
GdCdPJx5abbp8S3CPR/du2IwnS/9+No2UaqbjuT8fQFD27Fe7wwIAF1CnWHQQq1W
Y0Ky8ClWKSSa7FnjV4ph7iwLtnmgpNks64SxajDc8b9HeQxHRb89BExfsjl9QqwP
qJSWvOsiCUBwOmDlRACl3wmf62MIWJyn6KwC2DerLcCTZWcSOpuNYNIYIx8s6XCi
4NUXQTRZcBw7xSkY4WyzAG45cgCpS3oS5pesH4HlSSEC7qH/O5BRygnpUxMEEeds
29mqxeMOrTrrysJ3E9HUFw207TarqkY6RAoqmLckyrRwOhrvo8M4mn+mnC/Wmtjn
lS0Lvhj4qwf5j1JOLtavTqe3o0nToVbpfCRrish/ZPtDLuIwIE36uzBWpZNw0FvP
THFHd576Jjt9uU+8tsJ1taMFpptJfhIMVpEAf1Kem3/7240XDhsaa9T8W7WdxjEc
9blaBTQR8zc7yunzMX1T3xhauy+VoTvvVi33K/uhD0pxLNpEHpEVdn1l7oJsvmaH
5N+YYXPDv37QU1ogw9vxd52eFdnLtdd9JjKnhP5ybj+KO5udRbhIiP2I4AH+D9Xl
wFo2r0ZJ3cGJpBxJn7bA9XhckKlYSIwcbm05IZIRyzD+csmNvZsrJWC1eUE1/ntD
I2oaDL2FJLV2fZ4UjorN8XCT7GChURcIYDjeOtA8H1VzVhJnZ7nfHbvATzsPogsL
IKqbENOKrIyknZ5ptD3ouS2SJyRobJ21f9OK8EEQs2co12lV6iplLK1WQpboDdwf
g2/WrUMq3SSxnsYNIQaag/1ctC1uw2u0o57Ucd/Js7PsRpjijkt8fohBvLwv5KKH
amA6Do6BPbktFEjyM1hFzQblut5sad/vVIEP8XRF+nsm14aQ9BNPxVQYSAz5FlF1
0F9VG5pV7/x4+lIfCA4abP29+PXPDMQxH6GT4vEoSo+f5y6XfPBBroYNe0YIZcNw
4jyWcf4WET+mjn+VbuzvffE8LsC1ClRXqq9/8EKI1BEZqmBdsKx2ZAG9FklcASyb
SUc1NvzvgTTMPeJMcPly5C5yC1J1hES/Nn1TX1JKIVO5YijpeXxha4GCB47Cdbnm
EARWLmz0yQhfA/GQuiRhMDoa12xlpt0B/xJcCTm8Xt2+hrvZwKI/9I6bLwVaZvhE
AJrvytl+eFkf2Spl3cd8rk1LIZbhjWJNhha/gjOUD5x1cH+Ic+ETxizKbE9tRCDe
tFg2WkZEoRl7Y+NU+8zAknr+OaGuDb1CCgFKMCpY/FRE5xztv7rEJlEvQ+wNKPrD
eOb+5LVCHTcjeKCNZzb+7i+ukdDxp8IYYog1Pms/3GTZc9KPUNvo+0T8tOCp5p3E
q8vYyRBhP13Ea9J0XJzdqCTUxKl8CJKaSCgrA7ZCLpl5jRNpS4Cjsygx38d5xr6C
bUg4GzfrxThsnNSdw7EaJxKwigMyDn61OVtb9FaoCYr7YHoWS/LFVDyDeztk86ir
usx3Wfu3tl04Qh6OsvADQv/Pr5AehJat0lBRcChY/Nvd1L7BDS+Oj8tMBYMpJRoW
1OyzocJXqCSX52s4eDp4JxCEvzn1oU+WYkkig2/p9UAiU86E81ZQJNdsrn39R+c3
u58jmz7w9CVzkTLDuQByHF25csi59tM02H4RY5TQhsFwOqdeq9m80m0asTKNHYJB
8vgB++0ZlrUlduaPjNZeFaJe+3PJlAtlR9GcBrQ5LskXrImcH14HnsdT0dphDMuF
R0+D3xWMNxB7dsigsrUr3hqDe0xEmyIwG6DxTP2SD5oW6iuNllFpkFHGwMIjWbJX
UtMer32HOLDMqw6TZAvMAd8nBLlRyB5NZPLCUXLHFl58fLux1Dh0kdvYv+IDZvSa
VZPfqUsBwt/MI5b+9txX/X3QlGnlh5cKH8UZUO1aK29S3CNPOnmIohLq4Ogvd//W
rmn/ZNjpEwg36g/5Cb8Bw6wSbMoZBuLY/uYORyeaoVg0kz4onU5lBb69sX8Ol2bC
6nCe1QymPgjF5A9TwWrDQvmlu6C6VbWD7S/1lbIHYsIWZw4bh8C25jwNQ+pyYERd
2PHd9kd7mD41vdnkGscbJSo2vBvP3prFqBQaux788X25sBYKj4dNz8uFcTIM/tXZ
5EH+RjHBcpeWjyjOkqU+hhDlvfNtBkNc4GPhVChogGDiyqId+ArmNZIFKFvgTxeG
ph/QmszSfX8rPbQr4+CNhExdE36BYV+qo9fbLllwT4HnQo+lBH8OENy+kgNzrPwN
TVXpsOmPnEf6ulzcVglzgF76Gq0ySnCDuVgZS0Fw9tsBQ0a23KR1VHxg/SjyVEVV
TcV7AVBmSf0a8EPqOySfUOdMM2fUZq3cQGX2gcjwtA6Yqiqy/04/mlz6nEJbTt5X
c068jQL4PzJTbzvt3u0sZu55WmEj7vB22MTz/quX13Ydww7UWKW14rxbFny3lQOG
1QqvjSw9GiUOYOYGvhjTRLnohxVRJ55LGElctuFPDT4a8dMOYjqk5MJndlxuNy2c
72Efa3Ihhy1DX006y3cje8oor9pOQhoVlnU4h5+1kMFpEZidQslT+McrRsTPzLiB
nkPwQZSIglPdgH6eVppZPa8V1snE/uThH5Vj24X+/NP/3rVO0xjnYCONuwzAMQmg
GXWWDZ2cvSzN5iaMl4ssfggKMtI+8pzmAEm7QVdZaH+XuoEXJgcAjAeZDN4ol2F+
f/xu/l2ANi5rq8sVogD1MAQhqNct0vqhkD+O+WcoNhSY0zjxlazCwJVjE0a1eYhi
r5SI3RFmswO2NFQ6elRs83U8X0DWMqFwJeLgPGidf3EAswDw/PJiTOOTTi+VS0WB
uTfwMZ9BAQ1r0o1hTbNT4UJD5SzFDeiHSgknPey8BKx8iLu71tNGc87PZTGZfF5I
pgduBKb9TgVz9xhfVa7cRQBBxk6IgFzL0/Tgv4FNbZI4ovCZPQbjbcymdxGjXKOK
0v/7aTQ/eCj597EkiEl1pj0IIRFBNHcIBpQTHkE23OKZBmo8guNsofxrLWZs0gX9
N7pEZVB7PNkT9nm2w6YJIMfcL/0WSiKKR3t1emEkTjBvFZgMLseUg3sCH2NJaHtp
+mYNCywXliIvFiV7+EOHoiecq2uWIUaAIFM8tIdFPokpypANDRh5rCXgUBJGojhI
YuZZBA1/8rjQBi+mrmmlz/dnHsYxk+NoaHjj8UyYrScqnZhgwXYmmBAJNRRQCy/F
FJlbMftre8EuMaKlB3qW9IhezRGPaXXVVhI1yUwMRSVG681S4FMv/udO0tgINSIe
yv9s+CaeNoqOaBPtHEPl1I0+Iqp42Inwgt/TyWvkYYyr96VUnlIBMMbIZlEtuKj/
3QecQtdWQjmFgt+nsb8N04Xk2kCZ3xQpPm+ZkITFtfv2FQ5a2WWdC4EIUKmNzmEu
RBiTT1NNg1G2PLQpxaqfsZATJSqImrPEFpuEUK8xRv0w8rxS0cFsjiT2JLO+BfR8
J+uToU1yAPus50MasRApQM/St52oMz0a2jSK+IADB2+1WpxUzMGVnu3U4kDGyid9
ZaU3zs+ihUjwk/1KOLyGPeFSDiMXnNIH+CXXOdjlsiG/2uQaDY4HwC31s7qXO9i2
bEQNvshESfba7hjAAUkIs/lNcvGBJn80wEYdc0whA09NhsbSvt/Yi6TJVMqNA8IQ
YdgpxCAhizoXgUtublyufE2YMPgBTTfFi2otofVadNDph+61//6OHTIr3XJYG1F3
WwBMos4TluWrL8VyuilsCFib5w4+TF8+JIti9MejQh0EFukyn+c9g0SWXCaYBz2H
UOOna6w86DbkPnO3AEx0gZWhK6KJTc80EUnYyS+R+pyJc6m42O4jDa/lX+fAoPyr
Y7UO+woMDWCocgpy+EGF593w45GnmG0u6GZHtEVwpE5FCkXGy2wXC1o9K7utsSuY
wGLbm/bMPgDKIHl7DaGOjUzjrx1qr1OX4jZJFMOSo+GCmnvtDh3n5ddfdw1al9vN
LAgrW2wh6NHNqBNtVMa+5tSIrphs3bjcYoc23ipNtUTfN8PuBgvRfUu7LVvqyrGz
Ky3kV7eJkZW2RnkTqs41JOS8A63WXKIzBMXbLoFemUYcbzUmQBcrSVhxhU2Llx+R
OiC898zO1bp/PatCs5i214/bRu36pUxq1V9VWZjg+e0253qV7zH5U0sdXTX9+qfK
E0QiNtEXuo3JVBh73VrH7nWig/IaB0nWMukjSRHAvjp0hUtG+A33jT3nEuhRsyvY
cC6ZiXXySzcKEocQ+UghQqCKPk46L9jJv+a8OknFhVIVPjnvcXHHmB8mn8u4rk/u
NatsAfZfvaKt5jMoECPg5wuBTpHC7BfqNqtdG2vAn1MV40Ix2RKyAXjD5QoMolLb
+V0BHO5fya/p+X2tfGF3OcvvpIk+BtldXX0boSIG9XPRHUGGinPX/KmvOzP0FMHV
xcoUARaAIbTa2LppU6PNqmFRNVHx6ATryh5KpVz/GLUU80Jf7bL45okumgh1hjpl
7H8dEZeLmiRbWYvoy8H96Z6zIIyWJfzxNljwtP1/JSh5DqyOqYSHdtnQmRV9IuFu
F20yw57uXLqwGvruEY7wZ1AgRcSSK5PvIzrjxMwNnT21qDtxlLqEpqSMnWwY00qL
NpxYujS/m8gD7TXi6gJn/1iXQgwdRBWf2eTZ0ugCvY7kzsH2remnRbzQxpxnh/hg
pRwsiJMiNgPO7oSvqUV8d0ei8xia9g3tt1h2stBd746gNtVsdy0RrU0fO+g8Du2k
OX1lUY0ckSm2S4MpOl/ao3leiUGyz/GK9Q7253zGQjVYvFD/rZG+ZSNth+zLiPgE
LX+/CwzajM7N4/ZylwjCC76RKJM5XlHjEwHVLLkoqBj0ickUDbxPKKVuL1aCTBiJ
NAXnqipPbeLqW0cJF5tLFX797CQ/pIYBbyybysK2B7DNxTVEqXKCpJu9WyitVNEq
tGa2P7N5+9X0po+jEkYOFp1tTZzR/lXzrVBTKEswcaaUET8uWBJcoyGAUNsk3piX
pOiKWT++bfXytMNdmvp4TcpnOLa1h+1Y7cQnloUOxFKAvqPBZhFIDCVwoLWOImJ4
JajRH4CKh5NHl3s7GihBpeo/46mU9re7b0nLNPvSWM04e04HhMlPXKmM3QEda3Rb
iVqiMhEEgrrXeDtz6BQCvQnWDIqeccy9Psw8BotsGvUK6FNEu6KOG7jqM0IgOE75
0PKE9ROLT8R+ZAKSWG202lD3Auvkd2r2b66xSYAMgmmPxNI55f8JTIp5S1Vk0pvW
YaTGAGm5/7wDPNzPUkvBXmr/sdY9F5NoV+faivWj4BnBnHb1V+0TgvpnfasxGSwL
NexAdPBZpGdl3b/arVkwSKoeXJqqyIcUK6RXPV12BnIxe2PBz60LHwJd77/DMd/D
przaELS8SXkEz/BYueiXMP+fq0ib8TfuJIYBD6JLYmZd4wnPJxykdLAYMthN+Zmn
9fWBzenkj8mXYMAg7asFOVbh15U48cYHpjf+nKTRKRxtGX8thlufDNo4qgUnSRQo
Ncr19FVAoj3kTH+ytC+5eitv3osg6rW4o70WtGRBWP1baljeuwIs3JPLHyvW99h8
Py9qUKTZYN9G//nJ7G8rHX2foDGCVQIcLyxtxCalw3M1bVFMQKhBoL1Jlf6xR3JS
hzIHHNSDnuxB89TEEvx2AxEs9hF51kq+r1C7KfTt+oYVAtF6iUbpnmrnPitNVUaY
w4dY6ipr5Th838h9poUpGUuo1PlH8LpLgKoOxYn0yapGUA1CniGW1GIrW3vA+vpS
viaRFGFSsXZrLcy2qslz8TNc6uoexJ73+EOvC4qHHk9VXW5y4rtIssD/OE0bMN2h
Xni18Nxr4NXq4Z/Awc1sOpjRO+KzZhcR8YBnko95MWZTziYnkVjiT+k+0C3hWnot
mT4lehnX69AWnD7ol++W1htW4cL4iPKyMKKkB8FEdW49k7q4a8TLDRphphHd8lQE
+aru1dzNr826I8C6TwPDVz08E5vAow7qg0w9s7k0Kw2j2LXq4t8e02NFJtuV4h70
ij5P+6QzHQWWKZ2vDuniyQ/qipLEuGfZfS+86N2Fi5ZWF0vuB8PcoanKi2vzQ5FN
MTeEeqZEXOWaKF+7qXPEDVb2c0SK7IA1P5Q2gUk5CwPyfMv6JW4OiLCvkazEvfka
MuJPcW8egJikisTQka7J5nA7rCB+EBTNgZC/S2e9XuuOME/3ClPRsmdj9w5Lq2P2
w1KsXqvGoPLPIS+YAC12ZIGV9BGk83GcJxD7VRkgivS072Ex1+7cOf3XbOjrIPZ8
ttxQ88fdRTlaU8I4wk3DM9zEqzKROhD1VB/NfPcw74R7iyd8lEDxMmIlz81o1+YV
gUnyVkXDk0scZLoP6HJFPNKzaoFHZPJDdboM2WkK9s+zKgc9Zu4g78fLtiJBLHAO
afJXiGIbno0HgsGTNxrDK2ZGwpjb0Ozvmdwfts4UoEy60fFsaxyP2cWCBThR5I8E
nxIF5aKSD5Rg0C33QRVwfljOTk8oDgQB7NupdeP0x799FrdBXB+ySkBm4Xx4NMYl
0ZFH3T8gQJVIIuTZqFsP3JIzDevLj1WGkBskAtH8CdsiRxO32dbSeywsojVFLj+R
/Fu/59c/jbQuqu8T7e2yI4RV3XM3n/ZfjS6Z3yWfnUpS7mm0MoydsKavdNZuhkm9
WoT/EBZP+grbU7WxeApq0Wq7X2O3i+6MuAq6clWBNk2H5xXR42V0xSJ7VaDLM+pj
rlB+dh9I1lQmUhN+sZQGcyRjoUzS4cNcHn7u2qPTKcfaQ5Jd/hl2cKYFpJKTefSd
SG6Bs2Zz8O68AwX65NbkzS3xR4xIG3/RKlPB1GG7TVWVzK2qAiw+xbi0BiXT54dJ
S0ZFH8Qj6W3/yZc5rXIJHVgqqksZ0C96hF+s+0fI0f/5Rhxp7KI6VV/ThrksUmJq
TaKrT4BDyKojvnbHJrE9AT/V2Ctcg7/cE5N/dewxWi7T4i52Pa5vT2krUzVFo563
v5oLOUoVFCSmRcP0hqK2kgTGqsPaqW6s4iF5yrtZ14hCVDOvwIwqVRVcYvRmq977
pyB3kVnOw4jdSuKmlCiCGxcqqLDcQQZOGWhXWcDyIOJx2tD74Vp0QYVQXeBt4DVR
EUJmKd4pegKzKFI5dNMMVjwvxgrNkqEXiT7YLDPBhdhtt7SjNRWSEBCAIRsH9Cc7
16F/rxagz3s8CaCdfAOiGn2U+7wcC6KkqmjuuJiMkqIkSZFinAiLrbmqd3VHykmb
42NFPPKiSfFI5i1YHV81i7L9DSaPYEPy+BsB21dfIPjusfD4+h8PWBXjS7KJetsX
ex4DmHPn+kaWSU0WtUm5a0KcwMa4Ms1xiPv5atf2lnf0FL0ZCfkoY0Tt2TsC+jNt
rOD5MNy4GRrH0S36a9bBF7ZLW6BMmVSoRtYDqOKi7335os7dTMwiLmCGxarzXERp
VkZLvB/TEc8zNGq2d1XxSW2Gvl5I8AJchqqBBVpbNQpZmE8LS8m2PlDHXcOmib81
G1BnMSSme1y9RzT60gq1yErJ8peSP4FMnErnFMFYL/2qnIWX8y84Y40I3s4uFib2
mq9GmLUkLCG8nak6EtwP3MFkZPKGvSn0mertYH7+Qbgi54THPYug1FknmavH44Ow
6L6MozEWTekYsTMcCOofI9pFTTQDhWkezvcI/w/WgeXAk/2+0qmFg3FwX5sp/4Gu
BCv+kb1s1eoVhfKk4FZQnWgONzI+QdNgyl/mor5CwA3TtV+yce5XoglDBlHafBBI
dBkiT9AP4+fhE8T2+Am3KfNVTxu8nnDVysDc99NVy5HO1UJLtquiZJA+kqd5f6oP
JXBt35+sqIXLrlnquyw/74+oqYnCCSPWZ9UL8s5XXgdToGJH3uFef+ahZn69m+K/
PmO4GJNTar6qnIJq5a9Uux7h70AYMOppwzZIaRDOyTGomSNG5rofNaP1u919KQzp
HqplGBeLdeT0WAP0cOMI7DwTkqCMEG6XW2B9fh6+XCsmcS40qtOwrj3lIlwvKGtJ
nHkEG+XztnoEOfJoVT+RuZc3v8jA4p0Zz8NALdSEKeTZqSeaqqJMQ0faPPaxA++i
OfApabvPBaOi1CxVhOHtIWEMuc0wsDk2hGJ78Pqg+aPYJKUSePPNSC+ASA2WohoA
xoqIiHh0O3tNXeLFY7+lajrDnQ7MQ27nUMKLCladSr5jZbUmCWp8n4CH0APhP+UJ
vFf9a1OoBXnQf3yh11S/f1XguEQ6+WaZ5b2+rrIof2/Z4myGTCb8Z+hJCTZARVsB
e7DUgU5Hi0WaYUXm3DwdnnB5mYSnDsQUKpoYhckIlG+rkxJzPwFfjrRjTo9Gu4Ib
kge0s78nLs4qHwgOJk+AvfS0zuDqRP5QtWf+k8xwwF4Wl+UtTlLnv5ca71L7uHWU
lvqe7Bn5+khvejBcx36ccaOdZghDVaXjRcrOAIy4DkOvtuVcnmgiSziqgEnXp9fa
e0SFtjfP8eFEsx9EkH9Gr5ezFTOeT6RJiD86xO6xiaGeSIOTd8fU+dcWeIFqj/4D
rBu3lIFrk0eu/CCIlPOPQOnH2+JbFYY1vpc+Ue+MlnFjDjb6bNjm+kh1EjPXXVwD
FCPlF7B149oubit/2M9oIPepCts7OSoK3/nlDIZwsm7qM9rNpxv+8ehoz3jOH7Nz
N1x0NlLDeNTzRtFzOp85WhKE6MXyTl59IuplE3OhgfpZ0MlrjzyhUZ2H2gps+RRB
1eKPMQG77CzO8V2oToB87pzy8/pIH74EIBL8Cg5uaDeb5ly5kSF68nICbrSyu2Fn
a9BX5lBJgEqcK02sBcFrJAj+jn3GzN7XfIvGdj4MGDOmxcwPPmZg43qo/8+N93eY
j+oL0qxaq4vwyBTUliZF5VQU6SOCLWpU4HW5N3Qz1fKCSI5vZQQD/eIq4NxWHHy1
B85TAdvp/DqfUQkVhWeHMxaUSniWBubU80qlY2qzBhfjuTmjSBNmq5xh+aaZQPMA
albjC29+KF6dwgabygySxtV3ad89DZjsAmaa2Lu6y1c8L0Bm4m0dJ1+sIibGvQwY
SD9QPwRn5xVVpoP+qZM3jQSYt0MUOvICEA8nu9iE5pJFDDZB9KzSuf9RLJIL/KIs
XafP/OK46IsUKnzp4w2XWjRH+pVPxNYBei9icoucqR6flehMX86iYKGIdGdYP480
LfYPa1qqzJf/hSs7xzDS0oITzFUZdfbDD/S0GeS08ixS9vL4ryrHmNXM/Qfd4+jj
y6QvZUEuGV4kCvV+xl3ogjrTpw17XT7mRS//5PCDN2hnVjLQoRGR/ctyPSC17OzB
16zmZRv5m3a9QUjZ69yXNq1s7nKoesgcjHZb7uxAO4mCxmnBQ/7RfJRJ1hBRjFAh
2s9pZUYE+E0nTsKOVET3V6ejnb6CC+5nTZ7BbxCRbf/nqrE0jU/8ro1ZBpBX+Lqc
C5KZaz5TZ+BMiZIiJJ55p7G9qF5XF0gLnZOhoT4lZ79YwM22AkD8ERbjWJgEwvDl
13Fn01ZnNmd3xVWRPmDEaqKFL8zf9Jp9OTlRQE/pSsAtwS3vnS6a75WPGVapJBBS
NKknL7ZWLxAuaBUoidFCsjajTiCXc9p+jdKTG8/MGsQFdRw1whT+PsEoWo5+n9MP
gEEipBr9P8TgwintQt+i/YMWMzzT6dCKihUIP5SReRCqRiwhiccoJgOhyYyscJZl
32QdkcjJYF5DBcoMPLihwTLMMQ+foEa9VKvDBxaIk9H/5XgInl21RyubxAXZsdfW
iHoAKIMkN1tJ6Py1NJBQ2Uk1tbT+Uvzog3PN0vswFKxH9NvxPBmt1wURfinnTHBV
yZ76etbDYSSw+6ImlFI7a8I4MwpSnCkEzDeR3AEyUNergX0MRIYmoK4vRNynfyOy
nM0R/BQxpEw9IRtNEC8nI5bTFhacwMzB0UXBhBryORxYdLtQ2m8jvwRQvo71BQo7
xaoFGAjFdYoUXWQpRVAQYJjJ0+Y/YDdGkYEsFS8YEnnhq/ZKI6+VMJo5Sj4EIOkH
wlzGGICMFRI8OgfKO60JtiqF6KvMAWDdELRYj0HLs9PFTl5SuJvrbGILJWh/9Fkf
PWCQggSe494CzqPMwLFYfn2taDe7bn+fFEFUhmUCoenCsJiQGVKZVkcFr562/bDM
L0BVYbVoJBYBFqT4PKxmL6RWrA2y/zIirfBgwdlrt5S61l78tbtTZbq7LbuGW0uU
MTj44YuhRGT59MHqZndlXGq5gU3KbKx8ajXYf/3nNF2GOSbee3OGnVKPtHq6VzsO
jYkCMDAvONwp4rQDktYm4CxQ2T4IQpPmEHHx5ESjLKwfhDKWC66y/pTx2rNZIsuA
Qe+sEGU2ZQOJQfnUk2l8TxUOG/Z1vSu8akKIjoRBDf//3X35lHnkdS7y9/sSsh0i
pHcHyDjeT0zNVz5IvPM8RHD6vF+t8tfl1yjtLqqM/UdHTm0hwQzslZzUIIeeATEx
FyQIOC3I0hjvXWDdcVFjMM/F08yWChv95L7GE3ZxuzxplFYFoeaxhBbmXjHp7l+O
aYnL0Ni/sItgDjeCRaNUvZc1i9dcBoxv6te0R+3G1HeNE57v8gG+NGWEFXdeSCYU
hJEvj86zPZ59TZ5+sXZlMvMOl63ZGhfiNgco/knqYJZq1gEq3j5jqrDPZjQKxirG
ZiyVwKiwEfgWDqlaDIPkwaF/Wi9xQ0JBsyxMTn3YpO2wu/Bsdd5NyRQCzGRsXNgx
lm8SEwcaoZt/gtdZb3fNNjWkf+ySHrLXaYh8/9zDYmdZcI4uNHOH/C7rl0p71EG1
g4RladnFAi+IonFXF//DKAN8Gh9OSeQMgKX4B4gQLPoDE9Rjk0PVEbI2lRZRcH+U
jZ9FqYYLX+VMlm3JJ3UX16518k5Fb+nQHicqo8rbvhm6Iytd0OtjPiq2b695MXMY
ZpNolRIITGKcklU1RKqgGYJHSNGkUCLo14oVWzbGV7UyU/jzM/OVZDxe79emw7mR
UNGCvNCATAs+lyPkZe/dr7E0IFqOig+mkTSBtpMBs3I25wS5fVNAlHI9YgjDnn1d
66LstNMTSPXraxqgl5AtdUdIYfNbgU2xLPTTJOZen4nqBR7YfqrL2xYzSvQlvltr
5sxyx+1neK2rSgzVCW6W7TUI+2fU7uWpzEjQ3So9TzQ3ZjVAlctbcJaI6Kt9fKSR
w6IsZXXNAw1eQt33sevLJnxyMKKG8waPntYSXrJUNh51U5m0BfHqH+eCN7YUkDWg
UGlgxwDbRq5psNn8kivCVwnCu53GCdzmWUFguL34nXHHoILkZYQFBCtGboHYaIN2
TfssOgDcjw0y4N8bOLbFkHdgA8j1GXwaoOqZOPgLJf1Km1N0VrSobWYbKLwqr7gN
txuMAajhuipoPacQ7oKZI9ryOxy7LDLWvVpSrRs9fEYvaK1f0sMacF39ppk+2mjN
02eXH9TRsLsxH5W6dxU+APRcocwHzBbuvdFx3dvzuglAgaBriklj3l6LaN7SU70y
FOz/b/F9G3+I/UQmoVibAkgeo1yIvTc6qMmiVO0ipylXizPh3rFbRTyjucvNyTos
e9+/mBpsMVEwFiDaFhyIxXAjJDd/tyOF+Uc7L6TKYJTTtpGo9uiEsXLWEpE29+u7
TK1ojqw9cDtkc0rfN49yoSzvJLHEv/wTwRC0NdbafeLMozPDJSXKx67Roy2smb8A
bQEmLea8HyfziM6GubI5+k4kjb0fNfi62hbKNkdkCGC1UICTsa685n5D2+PIQsPo
fdV+eQV9f3fiwJw+JmuC57P1rkB/S3ETfwZ72n+Qv17SyknTXBvMvRZCeAGvH3h8
q3aJ/jlMT4/n0fPI9E7XPct3GMHdNpLLn+CQAl8SzdUcG+HF/3UQ6kfUiwYzj4me
XvLDVu/ix+O5w1C0y1Izf/MrYQJBig7X4P8lr0nL3+bZPG89HlPiqPbaWoFKuR2U
npyKtHgCQjPW/+yM0bM2aNy8Kf79HJhBr/7dohIsPxoDCoQ61SapfuD6+WXoWcpF
rV5x6uU2qaTQnPSwp6BONZnrHVq9xZzaQ56XX/kciviz5TM3uxwtB4gSAk3I7kyz
UzvjzoNzecdXwcERe9fGeK6x3B4maiV5HBSOaf6HrMpCehAg2xTIK5SyaezfD0OC
smZ1Fba7q/5Oz3VfcW+H1QeX5I5/bYpn51FsnhMRkBlzdsBIARKOygFHeQXV8MfM
N3lYcyRmHdTPlGeJQSMhjnHqL6j4liZi/D5ZickCCmWBB3DzJmuYL4fuOnIa2XX5
E9K9OLtpU3QonYEPZ6/e2a1NiwXojVvvju5+Bbv2jNubOmUUxHpL0azGuGT5WRiL
slKK5TruTvrWrCAk9vn/MAkMPdBYoYgKjldS8OzLHu+KAbM8I+g//B1iT5aeUjaP
6woJhQoJS/nCFc0CNwjqDvFN07PCLJ/le8l+3kIxOX7LZ3FrTeuMGaSRa/DMYEUT
PC7ad29T/eFaVcnNi6huzAJ4kEurdaqI5NiIZfxpSF0q7nsUvvo7kGx9/BurudYI
C8MRgb8rzHeoHbevysp33EGzZ2NImmpJ+MiMfrv2ZmgwVkw/Hp4MmKPJFAa6p32n
56xuGck+Ab5CdbJUZ1XFJCzglPQys6GhW7jipTAGLmfBuNSqKs9oKfX4NH6pqfIk
ZTb9raGjaU/pnI3zQDNBGIXzl+rr/y+j2kzHrvvTyPvd92xWp8DqXO2uR66eevaX
abt0TlwiI3kXTPkMepeLJyY2gA3jQTiBxSNo/fR+Od562MU8Hq6Ag/qAAkVRg/Xs
FqZ2YUk1SsCHr11/arZmnVOMjo/4scs6VIxCZ8eD1pNKgCayjIdywutGH7chlUxY
qLDeoAOixpwBbVCRFuGoupTrdKPP5pBDMxb4V+XoQiS718Gxza/ucExc2AMPcuQy
rHs1pUfNGfhFXUNCxtvO69UJgImDQsTnmGumHIh8hhGq/swkPl7SWkoL2GUAagPv
rROtTOTea3QyF46zdwp7Tb91GI3DG9gn9iXDnVxz81xG7bjDUavYPA6jqbC9rbSu
gs1uuBn5GP/9+6Z6p/4l6lCno+GVzXoNqMFInCpFsWDaCupfReSQRbCVD3TI42Qp
Hm8WvWNTrQwYuibxt3KRI4VxACi+M0g6DQiiE1fm5BJQe4R+3dBEUB+NBUte1cWn
mD7YTIC5sie0Aa8Et+ujqr/jglwCLQBdzwQBXwz8i8+7rDCRbTMrCkP7LrBCQIoK
Vpvppn122O0C5dnJtccKGYMwz/aIsGo7F4EN9ZBMdKZRtTZaz8ZJLiidbVvHOl4U
AQjX/Zc/6uHzICAh7t8gAXUofc9eoOWrBSkWZErFWGdlBn2GEBdpvfiYjfTRWlSb
cI+JfBjnQCa4idQdGFTLLpQTdJpW/1LkAA35rGPfdM1cBC/3Z00o0ufLIWzrNko2
AaeKiX97DA94+k2NJhbQxsOQCwUfJjydnn1Bi++iYPnzPOCMvWUyf1hpOGqcb0bk
rhkELsg28GTaJ1Q8QypNd2lJJRqZ2EWk9SsFdZEMd7R0tPgkGMI4fbvxUvIcXQWw
1jwP8Gr7Sov9GOf26rWcbu3cSG/WCH+3DFL0KsCt3wkFPFvBdnuKUK3scVkc1SsO
OQAN+PjP1I/3iSIGEuVyjRY29OmLYf8KZvB6B2sLGjrjTTSw9YqS3rjRcY9GRJww
YP9wnLtAPpbvf5PzpsVkwv3yxFY7rDbuMLHWvl1mDBOgi1ZNDuLRAkC0hW60scsu
xeL4bDxVr+fFB/lZzQlbvR+kFdgG3YgZO3IKyQXO9FdpsP+vCO612qyG4r+dlV40
ZnICaefBRCO+pC6ZnjN9Y+uvZEZTKHG1A2gmgCbqvg+5SH8iulBztB+IehsF+XEs
4mNmA05ctyR2s4ZKVs2v16jrDkICvgQTdxOnUj9I6EVkE9cNZkkUD//Rs5UIM2hI
d2XHxV4KChKhbln0GASeZ+ndm1/41Ilhtem4pmzVBLCfgsS10Ms0IfZMMw4OMPyv
Y9XRN3uxYtYqH+6g8Cd8psf1cGj0zzzvREwymAXKLChljlIObNKcmk9iZpo5joZT
tC+LJyhVRlpNjtpJPvgrX+6d1++fS1jqFE0MRB4h/+VFoVVYQ/2/Vhh864eEVt8y
cfVb81VktuU+6hZ6w0F1T6e8faNH90i0XP8csgmxp2GWnzdieFNV6VkjqiGzpvus
f7sALAHpGogCbNJl5mUEDzJg+5vhS9SpUPeEpUed7BeOGAfQb3BQxQMRbH1g+38s
RUFbyjH5I+a5SpwdXB3y5hExFQYS9zf/LOzweaAco0p2/+DR2ANwT7BmVM00Obo2
bEiaH8dFcit3bq5TAqi0MD96/1u6vdJU7pgFuwm7vgFF5UdFhQtJwoONVICmJPuL
ZcIa02uwL2GFp8Zj64YGsD5sIS9X2zMvKe7GhQ8p1tgBMX3GC8sObIinfYK63x+Q
7NkMP5Fhl303BBr1jf4Wx8X6xGqlj6IKIywGFKahwn2Se9WvF/f3uKhoThVd01A/
BAPQe0KRMZbgJdeCn1QE9eHDX9fRgBiEzU+kM7Lk6bj3B+yId/42JuFlGetPfDQD
Feq4ADTp+SXLuw9w81ky+KptZn1qqbJpf65hKVqH+Gj5Qdya3514jo4CP58ZXmSe
kgwnrDo4agGtLFTv+r4kNCX0bSesbneJhn2OvQusnlTeMRis/npBHdrNPIbe4bnP
EbEd3ue+4/hkYYA/ds/LVco6Nz4TsCJGcuzVdE+ektufy7YjYe6xctqQtivuLoxa
u4zp0l+fsKxKYUNYUpGqheJmWTIMEbQ1vnkxvS0K8MWl0AN7RZgxeGXEL01DRf5D
7c/AE+Tjs2z2JJ8sJ68EIb7d4+0gNQqjfia0xrisfvY9LnZHbVJKY4iHM+P3B68I
l3otVne2Au8QFRQlMO4RpRiNV32UzwcTRK/6Qkn527lhaAw/JmUW/sMcdhVodbUx
MPZyQ3nXTJEzz/6PzDiytdz6XnO7ojPcYaX0VQ9yrO19OnLn3+A9vtOqFY7razo+
79F5QH7PpzLx34wMq9Mg0zI6fm7x/MR+qgywpe4qwTD8dbOOAcr62etpPD4GMjUN
pcywctji9qTTXeiwxDXs0lhWq3K710/hlvpd16sNnhqnqLiUuzPXF++plKOoB01L
pFKUkyKJQzQhudo72ZTnwu8F3Uwr6LhRaeCw6/HKjxee5Hcay6+z6xZHVAyBZ0c8
NmgU/4Daj+xxvLoib8dex+iWKGvTxN1YJNoucaQhOqLj/ESv91OUfFc/WffrLuQF
gbdHD1QqSohScTNsTezM1fCul2XE2XAKSg+HLGdz186vCdeSVc94NN++8jS59Z01
YfILga1uGzN41V8TIJi+32BVCWoeW6zhL5WTobJLseSVwbCdfCI/jAqQTrrxQu1I
m6eVg8bg+dSMsTgXy38qZ6CERNQES/zQgW2wySVRBO6v6LPpjY/GVi7oZUoZ3pKV
LNbyAFyFhLwO/TSiXy0BQwlIH0KI9k4WtDDKTXu/+LIE4eXnOLmje6DNVOv3VOVK
Ll9tvMVl2BpD2qW5nYHYvBi8BY/nQK5vxv9GvO/wgO7OwcUg3ZJFID3IstwwjV7P
IPeCFzRK6moK/7fx0bDY4C7nmueZry/6I0CgOmRxfrVHL2u9qHoyrMse93RscVf2
G901XmfQTCNIO+70l9spDqKBZuDr71BaaqRNTxUMbqR8k2MIoK7u7ewuskGUMsOF
8r53sUHebs7JP690TEzZHcAbjwHdW8Bl1/qpM0HdNiqkJ7HkqY0pA+W60k+xX8sY
S78EaCSjyx5lGE6JKW1OLRzWW5icR08u2VK8Ji8CPbUZkEvwVMCZmYzXgqxnwlRp
fgUoPSCHUgAaFFj2uTN9MFwQzZpbSFNYu33yUyo4IwfJF5icq/qXsGclQGZ6nupa
8coT3Z6vSSYjI5SA3HldRgWaean9yUvr6uEgssellcUVc8CT3Ngax/ldRPUj7drh
AjZKoIWyQNtBswDlJm1tXUQ0eU+OIU27WPZBiAF2qL6kQ1MD6tfxAh8tJSMZ4OwC
pFtk7l4v4t//uQ5/6S3OeUtzBdh8DjUjFBzX6e/16bdyn5nHfP15neMtoKZDjS7j
EaNjHfZIwIDFuiAfbkFKFNuGcMFmDpxEBjDublklnzI0CW2jYJuJsv+i9HIZL9GS
Qh/fTLU5QB09JVX6ZNloQke2LCz071H++ffrV79MwDXELX2+jLS1BnvUwcOu0Eyq
emhlmZ3e5qcrRlHxZBGcc4yoESKb68I+5+KGDZY/fBVAzViQqnY7dUO4Qz9JTexO
fXZLjTtWlZKnZkimNe4+ZQLhUUCkPKiBGPnfgvSCdiONbO4bkoesEz+/u93t4hoG
hDO7xRrFCGwCSZD0dSXDx3E5gA8A6E4kNS4tQUe9jrH+HxYVEPPtYGPGeJPeLl5j
PkOpsEW8Okwd+5ycpnkvt/e732dN5d6mD6kdukLfvcUwr+C11PpaHBf9c+CtPXrQ
U2pAZvmt4UMLvffJjJ/vq0CPkFU/DgRF4dMba1jCMaqOqSne/ORt2VVLyDu/Qlpr
u2sPIahIRORC1v3noRWgXzkqS7OzViU8y2vf0l7ssGGIfyohyBdJQs8TQgEn2pk9
pIcKEogLcZWwWc5ySLyerSnCtzd/BW+MUkJcY8YWr+vJlUx5QhwCHEvI0qgBYZ8V
b55uSIS/V2AOQOAByj/QHBclduqRxovWs/mvTPVQg8dHUsRUg7wDORFTFKCPaWbC
AF8BxD5x9itckN212OW4HC8yziwkfC6PUuxTvKGF0e9wCwv4JNVm2njVWXk0wkKJ
+VMCghFDdrACUFvYwAiz+MHpouENBuhmdaDFAx75U5Kb0IXuUwKJ7ry5mnlvLyEZ
s1xPyLLpSgUoRJQeZu77Ubtr9skLSQQ1gZN+0GP+v9lFmxnc4dGSmpwF4TJDDO89
Qsj/EgTv5STiVn9gcBUi5anfGyrcvcChQJG9PtaMd/UvfMgOmWt2rB/m5TL1QM3c
hi7is18U0s5ruqZjVYxONEx4h/dNua81epJeHREgV7bJZr4MjBDTwxZ7QRyaidiG
P2nexH+yPLanmQLOnigGUTddOn9umuB+9A+cIA+FRORusJza71KlKzm3jMg9R27w
mIMcNwJSYoWC9CYL9rKaEaw/nE6DDHPxK4+w0mNRciEU8Q5yD2qEmoJ8KorKezQJ
yWogyga1dKpdCg0U0e4RUgjBtNpZEasyfaS8OfAKapf6E6fIho5TGZbjT+YsYd3B
w1SmkD6s0bcn7GrByIQmKmZfZSmio0fDsaepAbOEB7ZrellAgn56HSIqcK8p6Lo2
fzHn02aLX8OFYfEk2fH49qDsJVGS/raZYw4qH/mUAw2v1uk+YRe63FhFF0NMDXPT
1F0LO8tDcKcfSPdu/43/J43XyYTkW9JOiG9Hv6hqe9NX19bUzAx7rT9Xozz1r/E4
gteovg7JA7rs2CLe2IlN+AWGsb8iYqHrvFNXO2d39dYUz/mN+U6eQ4Lwk1gaPETO
RmdAKMv6TOD49X+GGEpk1oiadD8a0tpEnTnJRJ3/ASPFpRyf5fxosNZQj4rJZQXL
0cX+ZZFzKW/6oeDeVkfThDo9f0svLwohcoID0/FkbFsYOAs594nRCi/E4BZ0aiYl
eSMdJuC/R4I5pEkeEO3scjPYqqtiFJdRAYxP1GUt36aG13i6ZmvExJHmnsVGl33V
D0JXfqs+zIJtP7VGvzGBXHACdA2yvNHhmE6/SYIAWED0HSykPlTFwKHapnLOM5Et
oqS07Jphvz6SZOdAknLyGXbSex01YbtCAbJI+V1aC2x6FS5XClYHUzj3Yva9Slql
nEnP+PnWdNmbByfYCau8x/PNz8+SAltOov9TLcbZ2+TXQVmO4QyaC/W4lSDN3vf2
pSzR/IQR3sF0SXRk9zbh3cYX9Oc1Arf98HuXL9eiOf1yZaSlz5ainkWEnU40ntea
+zV/pLVPVddle2Zl5jGlYZihPa2FyyyLnOS/UwH6fsqBLmw50twgFKwIG6C9Qe+e
VFN2hIJlDjjE/MXCIzBeInKRHd/JOJA9So/zdnJxGZxw9vhTyUJFNlEF7QP94RTL
NujYjDZgWks6V37sXp01tt2KOVNQWXwUy5IZzwdI3mrSwC5dpNXpBVNy+ro4ky0P
d5S2f7IIj4bsUmUmsqBjcPlI11x8OIcb/SiCUTvYtTJZA3Tlw3n0TnQR2JXPrPUO
A0JnGmN6MavSBvmQFQgPo/NdasX5/97WW1GCItPISsyhP2Aiqfz1lu+eVHBS+Om9
VOfsm2jaPGu78V6Ncd4k+Vp1ucRL4t10kX9KEc2cOYgJOAWSbW8EX29szezP6ARi
OfbTZlm5HGeg1dNRvL5q1Tm5/E9BnGE/HkvcW+F8D8GMccbp3pdkBc4TS7OK8cIm
oEw4ByE6BMieEEPTXfecmHIzexlmnkFICw6t9hgPtE6nqGmQdFKiyfsCyUNyxnXE
36VM1ENDKL6k2TKo1HvUGWbV41k/Ct9zOdX7p00NCJjLboFF4Qz7CdBnazK/mSsV
wvuNIgwG3DKpG3pgW+aQ0oJh6YLcvJRWZ4nKr7Nwt2b+JIHjghRyenC4+x6nV3xz
gyTpPWNC5biny+wPvSsJjOSq/Dgva71iS8Zu+xvsHyauakmRhk9+a1Imi0rkRf8+
ItXTaONnsBbLWnDA1VSEtaR5VfdWZW3YQ4nEndv1Y5+yoP/Sh+7DJQjVOOnzvZJN
JdPNCMdbqt8u7KIRU4s0WMB/a1x1GtYC5YsgR2ip2edzep4F7cKGC+UgJ23IHkob
PKXRnFn7+3Z7ZOYp4ySiwh+PmplZ1MKg0CFK0sBlV4QKHx8P1+3DH96cn6xDaHxy
teUcVN2M3QKcMeABoKGMrpDpECGv1U8LnvinbSJt1twIANKRYuFxIc+Khik2Rvq3
L/f8YIzp2hKuU+Ic64QxJHbkOCuq4Mlw0BixbJJcnef/Gqkn2x7fEPqGLKlo6wOk
+i5kb4oLAw1aqMGZJKOW/OO+04ScZ+mEXYWV2FJui4oE7Ysxuz2uPAuv5xFh7SrW
yrvDKhCxx7xOTkobfI1b4RlKRpI7rlrpuf237J9UW4uirgM057TJM9Ib/4zEggIV
XGPFv/rcNLYbtszvTAMramQm/UOI5bmCSFuGaOLyXm8Ds2e0Jd5di7hruq7ih7kh
CQR3luSLjIql64ODqp5LLXxzU30KjsaT1uW7JJvWaPbqM+GQ/HdtR7Sf7qXnF2N5
D7SagWUOmUw6VLhUrHRXJcZ6wI3SlUqoFCK/4pjWN/Y5TWT9COXfYH7XnkxaaL6U
4ae+zt/SOIIfiHA+1Z2q+NwwYOu44rzIFCdzGaWKpF0b9eF4V+hSH7iyMi2H2mQ+
Dso/dVp2ZNjNWxGpnaWZvs4oAAPmiI6V/pXznyAJZX7o5ppKnrRQ8brsKgxe6TWx
21Aiz8DEOEDkKHubcdGLtoUQP9zXeCeTEEYoULBIn1NJ6VRuqLT1+ZtGX2djBJSn
E1wev8zqAHiC5toSRB1LpbzL13p+yYcsflKbbW4EHnj+oVvUbvTdr96ufX3e491r
QKo4Ki1f32ypQ2rQZOvLFMVPpq9B+zJeXr3TubJdlyJxShvIX6eUiguTFAROzVB8
dS5ofhMKPZlG3WU45u1jY/HU2uKdVmTSDq+C4A0UKA1Ls/GV4tQPt4ZCzzHhRtj6
1rI+WfXSmVZ0whl3GfTeNnKC3zQ3CPbiLF4QaJlHs209QLxkkIvm5GwVKuqcDpXJ
9KYZKoyaJy5ikK/qHt1xeMNQf9e1ClGPp8+jQyjYs2qWPwUkATPspFXu6zwc6G+I
ncG4LuqWFZCKYrjrdY6vohMWJSMf/Ao3eTWMJ2UoSzVAHYYuOO7rGgCHIA3gwF5N
F1MGYSFYq7PgExS9wySw1CuQqenptKZ3eubuyiWAD7sStmTThbty+wDhogv6ghvE
YNyAxe/3ICrJe+mJnBwzseC9eh2+8BjwVz19J8Vlneg0F6HLulRUrbbCaZAzHzyp
PzItgm9z7d6u9curwSoNbifqmneNsxIGO++urDoi/+nf5NwodiDpcwA+lzd5kFmt
Q9PmCP+SPaSa05rxQpu7KsJIwkG15+P67COuZWRZtGne0cZW3RyNmtGPFPyu0IG5
YhXITAq5MtEwez5E/B4eXcJRvNdEHcJSEomKDqcJjZPMGtLzsv+GFuY3sSnq9BWV
3tLTMJxdmQvRvLe1F9LGtBf3+CADw1Hy8BvfdXmRtMFBbPEcTtLPgYTWsd44JOTz
SH/YTxGNdZEBrQ+KKo+y5mk7ZrXOmagzatpbLB0sMSxUUaeSeUETpAOSFtib2tM2
ive/VEZXFNUhB9SfrhhMVaxVG8O/7Tr8VgTvK0I5E0ZPgPOj5/EAgMyZ+Od9JszT
9bYV+g/Ha5898DrJzkkIw1Ib5kq36uogjjsNEGaS7f4L8tCYPhVm3DlfJ3SWRsOv
8kUgGNip5SHI+Q721CvEUoJVKxsM71hY9aQco273rlgPpqVX1BIP/2VS567ih87E
H+bqkgkxc/anOkbFLh8KIphIBeueoJevpjnfgfxDxeJsrBRZSo/fYug7gUG3s73d
imoalfHEqFe4LfgX0fxg3csgkXszSE93/zWMIEgpZbLq6/7/yRs1b5GJy+cNjdzz
fGVdvniqidqUHtpZT1HhqVPiS5UDm1+wuCEaL/9Cl7pQvDFXU5CQAp+XZiQpekPJ
UFVe1wTUakUoS81F4LUsUf9h1mCFuCCs11wMKsQpPavA1CGEhcUAuzYj18U8HjUr
1aGKUnhDIq4rIRMU05KMj+F6uhd5SMA3ouptfM7YSkGq1D4alno19UzOKEQffD83
TbpXSWzqFHkpKuUPlalIZUpDiGaTpDu06lPsA6PsLcIONOeMZ2JP6zt682zZLr9S
7bki6h9lo42qDzZLYiuWEtUJvmrpnLSEJc5y/GQUe+5PMMUB+YxQ8AuDykhyRLjW
ft9gSqTQCCgqqI6whYl/1nF/MjG6Abr7LkXkfjS4BYypDvvjeD3QAEcFX12jECb7
n3Rb1zU3M3tlViw1ZK90TpPo1iv1gMH0wOGjS854ygoXYH282coHDgGxAVmqWoNz
ToHmgHHezqom6Ucx4nWPPG5sAhgRJg/qGC5I1YLSEd82tDR1gwSbvSQ6ORG9lYur
u/gRp2f06riPZwE7Ln5A5+pj3d5F/b4CcSMTqWfU4THEDuvOYdPGOpeFHIaZMtjn
TVJYoJq0U0Zcz8hLWIgLC/vMYS91CK0da1Gukvz5HvvH6jV2RUcyoDfJHOfjB0v3
ckL79LLI2FlN/TS/3UykDx1/Hi33bTp8Iofry3cSsTo66lPV6In2AvpwXqUX4/hW
akva+0PN7JSoRR6BRNhxH9q/I2VgFRR/Z9vLOy8/t2PVZJNaB/DELfElKGiDXK0e
Wu7PZ25mIRVEIz2jO+NCQy+Dv9Gv6kaIej+blysI4cCTCAiazOvE7VvXrzODytUU
dtGZ3iroN/C/+orAXpX06ljQ55Zw16NOVH6Bb/IyNXIQgm0aUHjkhaWy1rKyVnF1
xbmbBobCwYxg6kz8UecYctJOCado1m/gxvznVK6341d2rdBpGjgQr2pD3QoD/+XE
Pdh9bZd0DvbvUl5uuiamxAy6iCgDHOsdd5g1jbysLDQzYA1883Qeld11moepjoQ+
YUCtiZOS2Wb2craqK3KQgHrlQYxi9+aVfn6mKEyaBkQh5mxlABoxFybxIL4REX8a
8iJv0U7DpYumND5O9jmwnu+YiBdQwLo+gIJLcr6FAibhP8EB5MbUvt+No6oe72VS
XQHSpaoqHoeXAP+8WFnfB7S7JAr6EL3fBDj2/z3yh2Pcsuj7Id31TaDATHwG1axA
1WHu618uumgjqB0ZobnzkPlJ2iSMhtd7vIiV4C/fhFVxeauMJMrY+w+YfbUrCZUX
e60MaHPgrwWCSya3WuB/X1fl4WXlZ6YapmfY+o1/6FC/vECDOp0hsDPAtJMI0Ja0
wN8cNOrTAdeF4bNtSAEcC/o70dGBypneH2H2cEQdaAzPb/OJ19HL4C1FLoj/HQ7D
qIsfi7dAvKG8AYFz3jKRU54TDBO+EUcxJ8RFfVzODODi8nR/pZkr2nx5diq/SzsT
v0SSNvuYVHQVpHPTIgrmCt7AR74UwSYo3FVchpeHUcHIpIIRXI/LK7Sczojpji8d
uQ6oZWQQYa4WOQ+s+2Bg2uaM63D47DwmPevuxrc6nH4C4JOcFHKG5eiYWbhcuKSK
XfOlkvqPEt0+ZIWFJUrMuvc+EZXXg2h/EBEGKASTxNVVLIzToWXLRghallU486+Y
QoxmQ8jXdMTGr7aAVSKA1G2JUN8x27jP2crmsFg5xFF5vFVU7w8us8cPt6f5cv2E
vIchEaYdR90i9psOjejQW0qHnZLqg49cahHB5ctSgZOtHWgQ2jEJiPucUe2Aceb9
3UnNfbMe8YQOmEZGt65cCeQ9dmmxaEuAEWArNxoGgSxLKgf3zfp4jZ2dDm9LueaI
o5GZLhoD7UWmy3Qd2XQC4UMTm/x3UFTYgpsKL0t5RH7HldSErmOyjv/g52ksCkh1
h1JHw0MosJ878P2ON2gb/zVrxXTqNgTZq0YYXafRufVyVP7JHDubfJ+D5+DrqNZX
WTF5cRX/54EnoRn4+0FZrKSz9OM04fnLj477MFu4AGrV16r9vT9K0ZW38K8eWOQ/
09MfXsHfJYV/UM5itTolBkWQGrnqoj8Lw2KR/WzICMIyf05W4PI5WmZi+DoPEFZ0
2yKg9P+Mqv/Et8VShyfzH0yLr4NrF+araguFgduHAICQ33LB5sML9aVt7dQSTQF3
j7pBS9kdBslYdGJsXQLE26ia24JKD32w+y0NBcfu5z46Sk0dVDH2UveDUcLhW6b0
slFGtkN0wolU+zBA2nj0IF1VBdTp8Z42yE4e9Epdj402gImUKKCJTYxr4FmmghTT
S6bVxYXyyJXYQGN7QevcXNIJ9BEJW0Am++7PLOTrQkYKgJF+oEhexDWN9iJmlDMo
CX7ExAxsZ1uwEgkjFGD4uMxdQPpBE8ylqUGI+0yiJOSi7tOYfRnCqVAzktouRdZw
BG+wUhKtsZdXnbzxJR0HY8b4RqqxP3qjm9gPpcxzdYZzhDZQQusqW/v6BDIem2y5
5lfDmiEisfrJa46+so65OLrsehLsr8MI3Ja6gN42yhAeSX0QUx8TgLI2SwhPHaFd
pcK4PVjnhtOzZ1yKj5PDCAvxvcICta4TmaQnF0jIrhd9tH9PqB9qoJckCFj15tqN
Af+LX6nrvY0itM11Bthzgp8TjHWu3VI8cu0w6IOKn+FKHrhKrfNtQADOULQW/8wH
r9T/H1CgltkKCbEMsonVKfRAE/ONhFR0Gs+bWsNOZJip7T/9O9ON9R8UCUUVZ00S
OuaVM66q2CxqYa610KmaZCgO2lFQlDhY7+sUSzQ3BBge/e71Jr2bxsuLaHNx2bWE
2QGacx6ElXKMNyUcrlPzMuokmi/+Fu7fg+0Ytkdc0ssJ8gHhKeRPvfeK51M7Kvl/
rgkuAws1iZcuyZTzkt7o4IIlW+RjiMq8UImIBqWeX+rUKwYIofFreS1prKUr5Ic/
GPjL+kW0UAk3kWwiOPAva3Tgo9tKBlKNJIX6A7isTWuaMp2rL0uvSxvGaC7+jB/T
zw1vDfGstRZVGm2XI0DvpoL+nRUZDWkWYTnxrbtEN2E1VhJuME+HBGUWl5sI8mBS
dLPSHXBIJVULzto+H7xJIUY2roBCZWkRxeDYERbWlHT0WawYomS0xiXh2AFXvoGN
Yni3fvYJ8aQO5xDRii5aOaZ4kAXdm+9muRpRbyYKRPoSjmQbknBT4eIz5UYXM8lS
oTdI8gfoyNZOA/okdlZWJPXGHzUbyvCbe2pgLgNu5Eo7mDSpAM0cePAA5+Vpjk+t
EIuODmWySfTrHrn+k2uu3SW2d260WpHT5W6PoM9bWzXgSIKaMuPkj4QFhBOToY7k
7whDYZV8EHb37VvRsQuF6pEa4mVGq4xlkOSq7dwcXPvRrf3r+wT1s73tbOKVZcnI
0LNfdepksFHWd+vPGRIAg+H44AnHIIuAlpislcCo5FvG9X+CHveegGv8jaXwqZs/
1TO7xrr9tzpE5PHIgEeVra2rUWwxnG9wxYw3nX9IuB0YYJ25HqHQq+yqxUy/Q5Ag
h6Jep2QXtxjDOzDQO7MU0WI+LQ9yG3QcQGELe4r1tr5xddAW3gp+RhIFUFdHJv9J
ViN1nQHJVIR1gAez3IoWAz4SbepGOe8HVbEi3XKpjO3StEsU36c6+c69j9EE5HHT
1PubIQeifqJZJc+NjUYgfC46sSNuw1JPnw0kZhurZt96nOSyJfw6XwAJ3T10RQ56
0Izb6nRZDzuqUB102bzHEo+kK1LPx/HxncPUfofvyCDeLTKhE9CpWqMP/JZXwqbf
kajtiBZ2oa8kuuE83W8/nX+gu1EbViKUiAo8x770ucA1YkOkcARtmKfdtnVNx8yZ
IvnjWUSJIcu4dSFeWtbkTd56pfgLalRJUgBcUFgEO8z5iFfqPpKfDoJM1IOiA9Rs
jM0DwA4CHzvGwOpbdkMT63OoPKrV2T3VOBY4ylb7kYO90kO5V0n7XtBkp9Madmif
NJuyukaYeFUoVIhT15MClqhxiFAcU4t4xObY2bR+MlXtllWrvOYEJCv7HinJqs5+
6q/O9QF782MrU8Niu/qkRx2cnlaW1TOiT9u7aIhkYOvDiqgspdMIJng7NSEhNvEI
Le1I4W1DOuZrIoIjgVdA4jIrFah4D4bVzltGZfIVbUs7UnLHZVXHxQF+JgZxEJuj
8dNBOg4Cc0j235ZhceX610F8p84RcYdzsNMs9+4nqUrrJHhgBKT5QsAkT5kvFVf/
kYQJA1/yYGnaOw2Ezv6lmFgpU42nVpw6V8LiAZFuY7TP5M+dt+FX1qVjAHaLBvzz
Tn04I7vkCbqEAbLp2bj/dHNUkm77ktqKJ8ij7AoS1v4GodltXR/4xm8I3qKVb+Y4
mwcpD4eYwcDGL+T2gePy205KeLCvrnSNHiQyVNU3l8ONxJnVSjPBVhTzPoxwXMTo
37CfSotqadx/3JLIjGSm35VdWcpJgTN+H8Nn2YisYO4AgbCGkSvhqvSd3keu4G+1
2boGFPcNQn898/2E5+mNrgqTDJO2wWcm6V6ntVTZ2hOLGBi0i/YCV5Ph1+BvgwMD
gMtwp2vwewR+e8nGyRfG7DNUreiayWwyWQSgzZHJ0PnN6d0mopBHvoBmJ9k6REkX
xyFiuSF35IR6MfIxnQlqzK/i1FuRoTrJDyxE2IZGhUmQnaULo4jEVZ6R/Rfu1OGl
YO7pe4Tbz/+0wSeys7thk1nSdVetpK6YikO4WQT6r9MwGf44JArwK4oT7Ygcsrwi
hpqfGbj1kIfv8lxi/9n59ndjTUMbKhX7wzpmJ5J7A70Bjfkg7QfeBtfoOIueS1KF
LcY6HFsHFcZBQtwxxg/nFGQ62r0h92We2M59LFHe6/jxHXDjPkksjgDc8o4+CLdK
vBGeKK7YynavA1j7H1nKtOL81dvZIum+c+Bvrm5m6M2r9RKlac8g+a0v+vkfd6vq
vqrX4rmuMgpifJuJpdfVq/3x9rfau5h3frtl+vHv6FylVc3rhaHOS5Z4xU7b44ms
GPMIMVJh2U6dMKAqhUGWej1yXz3MnjLFkJKdj0lHtb0BgqRDZeBQGQr6STMpgqu4
xFvqBE/4twhYLrsUoCv1TGwhACTMDHTJ71tbzsnbkG108sHzMB4ywFhjVUmQQzTi
RhF0nXMyrKuPIYFvRrKmpI0YGVmcUvNJtxzM1q1/usupVPqRm5JRQX2kaASgo+N7
Sf6Af2+KchlDldJgu4CiGgDsYPdmLqO6+w0Ic5qcDrgvfJvJU7sSfxw3cy4Q8K1s
IFluxu2ajfV/tRxAmlmOYeqjJy7cnsixJTZTizVK4GJCgMZfdi6G6Mep8iUegDl/
2J1K0q+vPaRDIMuYt1hel+7F4cBKKMRwtyEhwIkae5OMFbBo0hCMt0tcF5jiACfG
QeGZ6602LOktoo9722zAwErXhn4ShKx36R+lC3hnEnLrpL2i8FC65svUlUBx2wKh
GuEwvvFVQRqk0mahXICN5RFWfgi+9Kxn8gLfzLFVe4idlGvias9vEutaJp/sDN70
vule32QGkqEJUoAJre7BxxLvZuNFMilO19OPkVMM99eU2LTnS5rk99Vf3Wbkq/X5
wRBU9qMM0Nt5r6XW51JDVBTzgflY+QubR53W4ldksbwjNU+mBV0Cn01roo0nyR8l
1rWBjIaHRYf97VRHPHPozuOqxeukMRtIvosifD/ckBMjiGKVTgVkV8rNgFyzse13
xcvyjMVm4fywTYrx3ocwtVhoyXAWtvBdPJsDDmjOlrkSwF3tmzFgUnj1QSy0l5Gs
ToDWZ+J71v6K8s5HT8SG73KrQRsgTrehb9TOnghvGMNPWHZH81H3FkHM4e8BpFtV
aX3XZCEGwSIR7FRmY0x0iulm2FuLA+KkPO6a2sjuDf/NTIIVKgmkRfuUEUQgllQ4
I9nnZDcKRU87DLHsvN4fOjIGnlwlEDbJhdgFtBJigIkh3OvSsUZAHEovcJBeAE7o
ckGefDJleL7Q+X1T/xS9ulehVqctH/RGIZHz5xIi7RC3v/6bn2Z8tqE/2WiHxd42
hdMJgtqLXqmzWCNBW+lDiT6OiknK2BNi1dQnP+dnVaHA1nwbjrndiRGfKfe2tLg4
DuG6kEittJlin4mEHq/Pff6B3s33J1FU/BSoQkuknLYGjYlBPqODt5Htsni5W+KK
kPDlUDWoMQCd5ltu6CexuricVNbPSBdo/Uuy3BTZAM8RVxNbXZY12q4SwqyCULHO
Cb+eRBED8jeL5b8NKWSVlo7wROFgzfg0R/8W3TsU7anvZ9koWLVXjAny9u97yU9I
MRZHp/+T3SgM8tSYTtSqrID7KNxV6ZRNS3fbMGc8mPOxnK6Yec8ZV7VHZiTu8RDI
dIsMzcpGyAPW7j5OdnmswFZv8wuX6KRs5xSXKTukMCSPIOq3dWl2rCfCGkCmI1Fu
4B2jMYWPf4cxFH3/QcKpsNEBuX/Jlh3eSA2+RwE/fUjTn68BmcaK6AgkFQWz/Bcy
+bcoayY+5LqB9NFFaGDZ2q01JqsHgV5LPh/A6HlkRW/e+EjjURbrgi4t3U13FIYa
TSLhPWZNfJwi/3pqYFavoMWkg/ngnlB8CIeUttt33yMFXTrB7SEqSbmomU+AnSIe
IXJhblZosgOFmpBj+QPnd6CPBBE+SQQIllIBsDocmtD72Y43i9Obmf4pLKUT8j+7
KGcob/TM8yr7UydxN3AbBS4q8KDL3EtDn+YY1n2pd+eeU1gILQqn8/HJn3rvhYrf
t+6/zEnEkJ3BQlv4Tqo9KflUsHaukWOt3qzxkq0VcPV75AJ6aasvlzK3RgEMLGyi
aeWGVU7kh7sAu75MVXsKEvL4LjYAr4t3WDJSDTwn+uNqDplnI2i6LqYXCAGTAI3F
7ODAfgKzk0Fg/BKZuDooQ2kaArW3orbyNkAS8Rm3jQ+32+LIknK4y2ODAZi1uf1t
grwTNk+w3heA848G5gjr7EsleUbRUKA0H5Vzii1ZQ6pdqNXjQ5kDttk5L2qsWx/+
hCuQmoyyyYjQNFpEVh8lG0eYJGYZag5UxkahsNbgvkW6KXf1xrv6lr7z+GaPLFux
/ImBZSXPU7T2L0tAmAgh5cJUJzcNNbPnjMpcOZXNaBIObyq9kk7sDBRVv3G6Y+Ku
z0hVBtLYpUoSoEEUc7UcLkZ/SkSQb/AQmzHMkJWsHIa3xBCIh3P84wEokkD/FiJP
oIRDDw0D1Bti9DAf33US7E9jeHCDDdUdDP9/xvGDC/PT3qZu430s3Nc27kOYwAyD
xynsXS5hAfzgugUDWJAbouj5og+aCdeoq1Ke+ZitZmKoBzY8LRV0qQ3dK/rIqlvg
9xx4SD7HIUGfXd0qLYcyrFyM6+4IRGUtiYARP0XhvoA1aqZRvNFAw9DLUNpgPIjR
fIpHk0z2fUqwb+e1gyiUENpZ5S+bbvd0qOqTyj/6qQ+RvbY16W0uUtW/6o5aAL3s
KuvydIPXxGc51CgxrFmwSkEuu34A/OLxQl9KXD3XSvQcUABmDEraE9koA20vOE2A
5JI3VW8bl3okquuVy0Zy3Y1e0QsPFhMnoH8Gn7U12x+EDbvVgCBsR+LcX+xfQcnp
4pxlLJxEKwQN1ov+c3exkTDU7je26l5LZgSgsEHGYo8Z9GnDWJjFbThnepqAnxEl
CCpBMog86ZlomzkL7MO6G59BreeMyd5N6PKryqjqcZreUGNhry14B9cLuZIttFpw
Hauqpcy1cgjGtqIeYPmf2Pyk86Yk7g0ICbDqLTgQNaCiQKBLtVFYzUzgTesxfCgl
bFjXHUlYr3tOPHCGgIX7i0hPnIW7PLo5qJ+TkIHHD81jVgjZCpK9DNFjzxaThsX2
ZxhVTiBD2lzOYtebA6D/LgiWtiGKLIMVL/qNP/BHPm6axDzjpsA8QKj2qpD/8WIw
kMrwBiicscpSYWbMdbspuSL/x+eo9gGYHb5Xr7XQUf+dP/7XFs5yJ1GCoZj8PLiB
y1U8Ec+YTIN6pLDbneSnecgpBan45DudjJRMf7rb1Km8DarDg72+4vqXCw/2rP7v
pitepxQ4gU3aqFaBClXdy6yGOKRR3ZnKWzCFur40xvRCQ+YPHR+9L+BdokYMAE4/
7Ijl/pXVLg3DyiwknBYlwghpUodN3YlRNBS0WxYdtoyZSbwgdl6CqN2eNnmXAw73
86/NU/07zTfVYwdJpHq5/GicvhnCzefInyENHC5JFhvzm0e75/TSOKG3Sh9ydB8v
4ibtlD/VrNgsvaorAUIUfBH/aRJwb0aYahfsagcG0AurBnIpuzaDcN2bq8FCW3eE
WjME80WQGJ1dxRgpf41jy7lXC2LKpvi/1SWFvJJL2Ftz5UTncpbH6/BcnTtTVIyL
aN/jWequR+t5YILLI8Knv2s1GmAVWfvSuNHzymYSd2Wn04uBGiN8fGdesLKJo1P/
RHnJc2a3wxNfZ4qkiXzUjZrXCeX4IVBME20/D5YNMnH9qvapQ1yRVy53dozTob3l
PN5Nc5Rqu4nyREUyWamM0euqLQSZGmK1cotRKj/IwclwyToOgHc/dEU2eBjx55KE
Zey4tv+fwdNEu9aZv4igDJzP1Jb4ghG1cvoIDHd7RL3Z0Vemxc8vGJl0fJ20MFAk
atljjNrJ/xgxhdWKCNUUEIMEsufg28D44ja+YPEQ53XPhxebctkLPCBzYWx0UZyf
bh/Y6dUSuIOcUm6LeyuRp72WP3iQjDmID2G4+FBXDnXdQQGGPgcjLkGGEhfej4EB
7fXdUxUJoS+wRRXThZQaBkga/NyAbKTGGakSPnW/FZDsUrv62l0N5/FTZRWLUc+g
i5+OJnX7qK1XMiF0TlHG8VBj3NVf5vrbUFNB4awki9GLr4CKQOdIVPlRsobXh7aq
fHiVcmqaT+ju2m5KrvnAlXle3pWfgUm4vboOmg9WuB+P2qeCXaGMxbkfrIIdd/Sx
DIfYQUq5PHzvI8qww4htDBIUrIhCz7xHdMtvBhlcXFVNJPpugalzNNNpkHS8/gmT
+OQRO9IIsr1mBlrlhD8y7wLvGOWOpcEk/rSN6cqxctoCXri9mlp8uT9tD9544LdF
mFTA0MUZSYwV2OAzJ4NhR/DekWkG85UlRlE/m36k5aiYfcwYI0R7DXlmR/YxjXex
Q1gEMMvRdlLb8TpgR5qUtNEaMXXOtYWqudeblnGFd8tugVNZ42ATW4tn4icdsHDs
reSIH2i1t2qddJSAwuYE/tWGONytfRip1RYr+T0g5TOKxIPs8KCDroX8kRUZM2Sn
bn0KpFir8zoeoAEHOrnwxqtOsMEhtWMeXJdRvtuUf5qWr5rmI7ilQnxjyZR63ZzL
+1DUvy3tDweOiaZLwL8rjtRqZozhTkFTr5QTZXmNAgg1Gi78MfU/tBXzY2FCfb7W
p5wORQlUpT+rzkce2lh+aTuK9/ssVm63+WPG230fF4eDt35vOQRX0EkMm+qMsaot
LtWZWP7ZXO6TPRAA5B3wGAxBBF1ILkaIyCFO65BHaTR7J0W4zdvG8cFqOKm1OLhR
vLA93nptT+F5hxcdP4nkMfgG5l7EffVYTUYo033eypAvDy/S+o4m2kSG5Ps3KboM
MautD7yxI1A+lHiSXXXlZ/Tu2V08mz4OzuZJYYVs2QQWAnu2yvRncEyaBW8EnHGa
0oB6UzRFCiACARQUY7q1NVL04DMXvIPk0EDCtslBA9F6pMC6PXvUwo5jTrjU5/Tz
ryAf1Tfjf1futycS6gAAqyjKep0Ns6a6FseoF9PdEdkTz3vZEFKVKDHGr5ZUmbl5
GL/CvXM/Hd633xhk44B+asjyxfzZc5ZizEhbx6RtxbVldfJ01zZy5rimaU5cL1IN
/RhEIDqE5jtzFuy2RxvQXLqKLY2FuuHSiHbrSA0/SAc7km0mGH5ouWu7QQLaPFXS
1jNZ5Z/6bgRgiOcdCbZ7FLwuIC30BsBYqs5qwFHHFST32dRgBPICU9sIDXqcOxSu
u/10QKV3XYsF1bSRndmD+wnikuYbdOdL3oa2+l17LgP0IwMesBnDqJyyHARiYPOF
trqoeibG53GpJGkcdbjjc1YQvm0pp+qyMAQ699olBuch37Uv41L+434eeLn9BbBl
T5dlXrk1m5MMlYt3OsGXQD4IxwsLgnVHIx7OE/9OUmYNxLwOv8rgVYB1/TDPg31m
A6xTZ1uJx22iZ5E+PPKqqFX7EN6D03kyj1zBKqV8x46tXtJchzk6mL09hzVLHMiQ
vR5GICui0vD7hjuSFQssqMYUfxmEdKLt7ioMTO2AyKN70cg8D/L3Q5Q8/UR/t9UR
clcKRBLK+miitLBP51AbpjRW/U4Y348HtvnmqcBKcBwmJNI4brWYSS1i1PMlixc7
xVPilaUKogYUBsekgXIYoilpOksR95XkJs97XdK/6sZoYePXR28LIz/JXLNuS6qh
iwAnY59P1u+iUTgTKjpOl2sOCtJYIZ0z0R5Xeyc4Bbhvb09T4OF9XwRItFdL6NhY
9TY2vDx6941IgdVQB/Q+SMyXJvQndiF+9udYWljMzD1mTJlLl+rA0dEaGaVBoQG1
siKk4wFrkvxelwD1toxTLnTd/20BOh0MvDmZb61Fn+obzFqSsta49l699sraisVb
yrsBUYkuYxcJtBiYn8nq0VjSSnWoDMLdGHIHT9d7aTWXgvebN4fmHXIxQIjPv/4+
i4fClHAcA8HYEqCREhmv1n24UPIUi6eO5/kxYcuXUxowUI+QsT4S+JBeJTBSArra
Dv4JpB+9nG0HBF05Jt9fJpizgAMB/8R3XRcs0OHGzeWgcyNbdAsPtEYBqML8TtyW
kpZVKAx4OOyixRzoL+W//jOnsp7e+ZEf7E83OGfggs6K87uSUwIaHHxVvu9z2drK
BLnSrPSiruXbCKKfUNYY1TLls2sHEFOPQVI7KX5VXgU+6WHyD1vTH2pDmsZGoEJA
obYBNfpMP2lcFSCu6Pj6alD2EG2pydMZ83JW4Yur3pTiK+nFY0QXXBZFzVlkCEkV
VXlzPKHgbn9pTHYH2WJ22VjpLKQBg3DxfDX7e/HY9yr9gRNmzhXztjVX92fzI7P0
F8PGtPkqWJNGvb8H7yGFUs7QKh1Z1U+39VZOSgj34sKOlhKLNlJ3fxBCe0DdGok0
GmU69LKmKVrCPdyEj7LTGPhBqWJ+GdcXxQ/3J+AcEcW4oP9c1zUN4+XBNAh+4xHd
/2uC2aIXGq2dhS7zw9hRlYWEtJNoQBbfNIu7odgDMqulwpn4ghzM1MSOxA5oAEOa
QGUBHpDEzoGQTaD35Xo9UgxNW011OVy/WNbD+mW5entvgJTVLkwHu1TeLF0ctxUw
1Vh8UOYfpVcfjqM13XJ5vS2GWAaGdXUkMITDvxNTLh2Aw+af+LmdoY451uDdQi1l
MJG+dCduv8tfctl3iCaiDI4uqLn8KD5+RARcf9Vigp+/OsbDscfhxpjHA2ELIUPO
YAqpa3iZWxIyfCb3p2As6pFZymaccTNncjU3Pqo5Hnh0Dqc4dtEzEPQKmwsTUSNR
3indtAEsBK4/VepG3itPCSrCDhgahvebQagLclLMIQ/qutsrH4SQGYWay7EEfz19
ulnyc7iaohXuPEPpbEnaWNUP7Q5tIWMzm1Ld2WHquYkYzg6S/0V20AqLmFLMNnDR
fvQQ7FLrTwxZYgGRKqBY4qvuiAaVWYBr4cSy4bwYmY9B+maD4BWuzxNseX3wrJUu
D6nglUsMKHSUoKX4HLBaMg7cCck8PLY7yxJ0xTGvV0tT8NXMU2Z5YH7yv+cYjwa6
Qxq1GGNTdkvYTq70f5wf+C9GJk+HTpH20pTGIwc0kAPJZxe3iPSn6eDoK1s/nzLR
RxYdhd8EW03KFpGe4yU0xjcv7sycXfa79EMZ11zrQIgtkD7bjEFB2wc6CX54Pa6B
PP4PkE54T0fiG/dFsVUXGRZB5F9HQD1iqD+OBEir5xkxWzAXL+GCpo1w/stAzklf
j1xuCok98KPSGOlW4bnLNmXXEb72OjfU26z8v7kdLErCW2gPJEjf7NefRRp3330i
0jL4ssbCJ/RhC3IbuRjYUHpPac1HKsQsZk8hYv8NJiMCzINvNoTdYiY38VFfIRdH
KWT3TQuPvpn50+PzugdZClln0QivDuMupbgo9hmmpYMMIiTK6mODhtEzLsiVCE3Y
Db8q8CZpgBxjdI7NULg085EeHi5eOgJKQMUys86s7VobzmIrEJrrwZJSC8JGdKWu
nMeWzQOboHzKuOfwtZV2oanKS8yoR8cE3coiaDSbBl41aP3pL/+TG8mL9a4oQ8L9
+KJB4gDaavDXjnPT2DOYgufY6biOoTiU14+AoRSWyVZYRIP6+AqWMXuMqzUnsza6
L6M7WSzHHOK/o0jcHsaQ0/ZbbMjRR+d5jbOeptjI3o7c/1wYGl5IO/mAH9RgCDWb
TMCjuq/ULzZu1YeEiihpUcGRPG6IN9xNClN9L8pnAQqDisnO//6N5FCxKkiutwYA
4Jl9sMuW1O+m85nayRREpAvM2PMSzhenApPEMkCCvZRO7rMoNV4NoXy+moGY5yli
1bc008jiedKB7fyrZHY4dSlh5rEs2g+aWTQ5HH44ySh5bFO90ePTwWeSr70a+cLA
Y4ZvQVOUgO3bnHEan7XoiaYg6qNW5k8iK1TJRJS/NjsqGaIK7QTKNTcMCx0czA3p
tVIpH3jt99qy80QWLDY9/aZ5bltN8RGj7pChjFVlro8TduOPdje61gpUAu8uIjB3
HcLNdtrJKoPlMlDNOaHmbGrWHG0BJYjhg8v3sjdNZoGGW+AZ5LaX/6BlTWiLmTm2
bWxUEYPxz9uRXTJkDrZuxDElayKYVpYN8YCPK7epudOQ1q+saNT86CQDpPFoB08z
at9q2G5MSlTEAbnt8tLH2sjXJqHfyug5cCsM/OdH2T5RWkH/KOEo9yaizCl7UwZJ
JO9W1t1IVkzNgYoDCuke3daSw+skZHhaFomY88M5daZLFDoWwyPhHucF/E6IuZ8T
tV5M8K+sSmxjVsKOM6J66Au4wRzy1H5GYkLVHfNB3aBb1R0fzOFGSdgQpsZrUxLE
G9INTZ1B2PKSwO8TVbfNcdqt4iOjI1t+BTlcdQYlKqqjI9gc/s5XJlIhlnshWc5y
Hz6ypQpdDhiiWDxDt/mQ9pf5ejZMgVTzFTWvW3/GvJWI/eOE8g07vzvIwVTxEVwf
bkCNsNTd1UShU7JAJUssXbBp5ui0fLQIrqY4He/0bKDGRM7KEvL2DBg7JheypmNm
ELnvqep5W12uPhZRde7bnhOppUOacwdDUN6etONQrcm1m3KDB8ucpBHM2IbLJJzU
CwpSY/SbsialAM7coXPsg/Y7r4J7j7EIMcXI31tQM1jaKMH2MM2YFHOmaPifJ1vA
5dEtQfKYBc/qSn66b4G10pbnre0N4wFC67VF5c8EiUu3D//oLd/N7WDi3Car//bD
ITB5MrPSvroZBpRPl3UO17ejDh8p4ZN5YLtXE5jG8pH9Fl8TUE9UEjXCq+0mW4xt
ybqCvCg3MVDzzFpBF0vC3/3mUg6EbYhH9BB6GQ1uoJfusjXffDHI7dNxrAxHEaRN
ZRQx0K6AWCvnPRn7oMOWMp6XlBBsqr/+7ARkCQqWaHoNxHCCJ4IsLEANot2TrdEy
XyEOijzrhHMJkzVXSMPKLCrHKD3Gaj/EWJNwDE1MQgJkwZ7rsTTxDN31xRi9jRbE
EZtuvk6dDRNTHThvlPXybwBqPOKGF4uyY844ABVtS+r42KxT0KQOBxBqG4Z0fjKx
mIwUxZisnbwQleXIoHIsEDPYAmv7+kGKWBKztJhMFkNH+04eRe3OBD9X9IlgYs7r
ka23pMP0whrSBK4nf24L0u4YPz8xqt+nV9RuFiS42+yd23f//dS+OlOXAkuVFFPP
DvSv8vco6NanueWJRU/bmDWxGvYe8sHspP4bWQ3OnjO/PyqI3UKc14eCMEZDXS/e
pi2O8fAiYPrd0RXIpDlLufSOdS8Nygc+LrWfwF0t6k9UNqpqDXWbFv/H/ryH/Mlz
3vJipn3M/gPU83yAseXZnKM4zOluRQpRjxVDJtg0k+8e/FtmM/UyWW4ElHPQMWwr
DV8ROcuN+w8lkRB9unJfmPI3Bhuxh/Ibrozj3+SK+PCxNbc9A2iTtzqHlp86y7cg
fJsk6mNBrSkkg9ADbzN2KFHJofeJF+eZGAgOmQLd0pwIicbF19V6MYZiBW1fAHZ9
N9BmPrEC7m7X/EJx95cnaaVQo0mlHmPZymhdvFbaPEArgxB1heEds5Xkop8XZImA
uBPDzLj8idBbI4yF7VQgXydks1uS40w6XD16OAugnROIn6ZhAjrvnpazYfpgyWj2
oPwJoDJ+SXFwjQ+7cdw69DhBZROvfNtjENGkTtjrlUJogAyc7JjjUHTUnvH5Vscr
duU5HPjXcP9WuYNcCqIR2HRt1Rfzjrowjxttp1N+Y5LJlhB8gd+l/WV8+7UgQPNH
eQ4NQiyJb14DTNL55r+Pubwvx6Sm/WCTahJOX4sBGu2nod273/HOvTDEzYdbkdne
JVhc1HtRfzcjmYTK3OcdadkdRiehrUbKvXbxdbVe9bsOu7MClhzQwAho6spVDZdR
RzNYcbXkWIL+VfW/0/xd2CxquFqomi6ryNbd7U48kDzOrb53j5heGCZO30DL85kO
ankmUY6Xt9Qpq+HXvLMQGjKyO2L3/wLPdVhdzd/iekJihISCSf0pJC7wrbErD3yx
33UpBDg1FZzF4joAgZLSoWFf5EbqU3RI8YVsjPFnMBuEzjCuPfmZPPfsO7/jCANa
WJogA4s8fYljZ6UEcqxD0zkwtdtbry4pjhU7O3NRs1IBKsCSAzZ2TusGsFM3xdNM
owHA/4Kr6wwypKzLopP4pKPRcyT5w9FNLLpjU/yFBFi6CgfBg1U6BxvCEvSa6Omn
LqEsD5lLddxMvNu9hj4e92562kuaJ3g6uriFyWnlxVHmaEKBM2lYvHJIKbvFrlhE
qLPckq3vTgQZntFbRQcoW0ulu+2zu3Iet3kRlByT71zT6GKcudjMt9+rW/PZABGs
dmiXecfV2wF27Bf6XGxLkpTGPyXIsNm03JAl0M1XUE4+pGDswGWOPuJ8kKdQPhQ6
S7E8W52a/Ccg3y8sZvpxQUJP7Og2dYRjZGaNJ17PzFxhKjinKKUuVMzQrZH4onTx
KVvLRu2UWwvat9GBIyrw3tN3W02Ndaq6Wdtd2c1LMNRfndLJa6l49NrzwX0TCbIn
4OCDETC3nHObHFJveSqQ/vlGr2N35ZQCcAXefBQDNmKs5sq5hD4qqKEy0sunBew3
ZITbMCNtDxzU8JF/ZU4a0Fr1KFR8H+YGK+TfAy3fDqwjzEgQ7/Yf2Rs73SsgBh8x
SY69dnQ/ys4B9Wznw2clpY5GwA+iulX8FMu8Rg+Gp55c2UU4VxqkxgUGSFsP+AB7
ubZCWRmU53IlNj4GSgJzbFEy1XtiK4e2DvuxaYCxSKM0zc0ewjLCshp5MhgHyLOi
HriihvP7Hc9FfNi4ib97J0g78A3oJr+J2SlnfMVrGnsGBiqb/pzXbZLbz/aDf+pt
M1z2HAj2wbHZindNvUa1SVdDaq1iXalkznxCN1WyO0YfXFy1c5bJoYwA9z+KWTP2
nryMuP8iVcukZK19srIuIhm8xAPYonBeG+xsWxBiofCLh2KUHixQuc395pb7YDb0
WT0pq0FXuw/8v10khfPupNhBYtMCmDLPBrKLgKzWAR/oOlg5aw0axbZyMERZ3y6H
tXHABaFp0lgXkZUlAu7TF2X6FYXAauKLw1r4y8HQ1ddIjoRe/FRYNY6Nu5kH1Sgd
e9rW2dg6YHj6XsPK6zMXF/gZ43f6r5xn60Rfo0kCirUJb2AvrFdUOEY4py0SUB0p
jHkKq8NjseoiW4UJjVWqH+2mS5JFRlJEMY0qvlSNsRC0jyvR3FKJjCDwHlfDg1/o
FCwUUeB54xe1T41QepGPTSEDE442UnzJfO8Vyn7ZsLTn5dmEgsyTdFHzbAqQzV9d
nLVmQIOGaQxV5sUEIh3DPE+rc62yex4uI8XlsUpUp1alktK/jK1fJrVNU8LBe5RM
iITw6prl1lqQHLSv/Xf+qj6fC4I2UmnzHP6hB+tr0UrTWaw9gQYDEou+YUojY4c3
0AWd4li18/s7fNuG/Ua9NanotPm6vzKXxX0VQEJDJiXhNpf2AZ7TJA7OdtfE61Jl
Xjq9K+IQfMdwpHVmMICw7T9IYltxMW38g17ieHvakPaGuVdRnxvWJrNVCIpn2thS
gBkW7zso6j4gWtOmSZAU2blamqRmlx8kIP9KdmmBBtJ2t5TiL/LaW83WzHi3v96i
pPSLm93eDDKZIvlpQgjBExHofpiM/zIab/bAoHzuLnQOTe4OQzybyKJQ7fnCEP48
9ZuWprxiwYBRJgyDcNXiW34fi0PvLJ+qS53rYmAqmSfzQMa2p3h3xHBP2H4FdMtG
GYIs4DJ1L93iMoF+BaDJz9yEDiETemY9JEJVdYUjD++JTXCC0mpXgDIC//PgLQW9
CGqYBBogzQhz8t22lio+aaSKnmIEOWqZQUTiGB4nsh6OlPK8b9C0PqfYm4qjSf7X
cShcCShySHdAVJX/Qk7QN7X1a7Dm9pGd21gdE+IipGVvFGDTnPm5NtE6F2p1FfuJ
Csgaa0XyrnYWP0V8C4pEtCRKZmZvwuWDogtBCOyRK00UW4CGwtn5wgGoQGQu6Evs
7pxjKa1+1pcxPmrnJ5fZGW+bSOZDoOVOGB4C0ihQjNa+WIct+u01uLirFtM3Jb5r
lsc464mOZlG9KfgdVCCFjh5Kzy4ZIaZfjGyukcks8Hr8VZVSwoeLKTB03gKZKOfC
aXcUafzGiHfNP7aZori24dyNqZq9sZir0D6qT6tbFwO6P7QMuN1rtRT3EXvetMP1
9ZO22JZEhvmBGHGAA3OsEMDnD0qso1GK1Q9UgJh8JGYo7Xg2BgQsRomgaJjK1GBp
QAbu2TVk2sM/Gp6ULd9lbIBPlfmzf6ZZ7MlgHyohs2ybcfedHO6GjD3Vd8pjxzfy
YTDgd2RwKLnXJ5+P750UaiWbOGNaDB9OPsu4wdhCHSNnybxNggk6RVwkRLeMjMuA
JLTOPamsHcJuQySVdHVgitK5CVKhNAB491hEebwEZV55JJoHMw8EMf6zlUrMoTyi
hdOo8pBLKBzmwYl7RWGxJMefuZMKdTukUj66ua4ZJwnXqj4v7YNF/IS9aEK1CiVv
rUqLgsIPgoO5pUbJR0pHARiNI6qfYT3hXxGFAGUjd/eU7DLBux1dwpntPk6azypM
AGCYLC/C9bUvHm/Jo46r7zmMEAJs0J5aywP5tfZmds5PlhSJJ8bjkxmBIvSw+xVH
Grj9Cazp5U29TWJQTjeVqneqPXrpKakQVQoo6puha7JnvVoQ6n1g0UekxnSHubVG
xfQPElqStWwgtdjdTzUi9mYKjSquCexZwc2hs5UDL7ctExy2eL8UmoL3ZxLAI7+K
y3PfGEsYufKgI1M5MfnNIW3VJna+UGUtbdl8RH5aDuLXBvRNo5qIddgpPxJSIWmp
20AzL8TmrmgjPWnNqANW6dMJAhhrRAdPSeCj3IRubaCgGLx6MPB9yfjGGuO2M1/o
mBN1QZU9zH2gxFPDHNyifqTugaRQK+8S6Ti6k8fcP3aC/46HyEZTcasTxkywJ4fr
pChSA/7b4qGQGqNDUsuzwMc6KLNnvV2cYlpjnUKQEM47FpHeSh+4NPzsEn0dn87N
oEHQbMvty+Vit5o/SyYdFXFXUl2ZiDt+wEs9tmUnAXCMHIgcSpvKYz/3tSC226fv
vpy+iwVzU9bTC2eWjsZSVna94cKQbJtLR3dTu7Renu3oBWYpxYvMtCbDk0NobC94
F4KPW7x0v5k9RS1avfKhyFHuZEG5fDz9xTKLC9auh4FLUc46EDFWTIiNWWim42hi
KSgjtBnehiG6MJfc4yF292B9o/f0oT1bkX6rUR6NjC2COBGEnRurmvqGst0eR6iF
M5ugxbOpQdbCgqF/BYvJwUm50dajq9YYvjn3Y0pP9WhgYkpMUKfIXKcurlvXtL5R
zPwEfXpb7+gLZK6RYhhsHZabyjQPHZxraTuHIbSOPdtcSPvpoCeaDDxZX2Kv0a+C
aNqwiuJUcFoT12uezPWykxD72SIhVHE2mrGxIMPCBqsW7mP8AhSBJ/YNj56PqmbM
vULmDN/hecvKWtgLZoNHXFSpGZwGraZE1Tjpnq2X536mnkmvht9/zVnGnAzf+5qk
+SjspQ+9RMwiZgCd2AJzL7y0J0F99Z2fwj0SgQnGn5w9JlqXzJjNYJ/uMIIpIuvu
e5FhaaIT3sPSEz8xsto5PnCejXh2gijJzYMtS3Aqab39tmyzNnmUwPFlOSxyTgFf
vi1YGRSTLRDaQbRxwsQWWtQ99xh+hgpNdbwssHFRV0OA4ND05FOo/GNXdiM7p+rT
lHHZ2JcQ3fBiq0K2WP9Pzzu4my6Hgeknghsyg27lT7HoOoNPIhvbrXC9CAO2gC2Z
fxMpvUNLc9hVXhWgUruqSEfuNe+iPOI/BK3HBFXze+LYHnABifMO3XCxuwKA9Kza
aq+MDVHb3OIGnGYd+Jgm2ln4orRmH3H30hpek6pcYVRt3QDa1WLWTgWzF72v9CJA
HALVkTUSM44sTtWfqheliuNQ2qgNURehoFpHTqKcMQCFjcOB31be1SFoR0JxjrqI
YX4uIGDuVtv33wlB1zMo6CZC4mEc6TJt98EX0PHWViRWmhpryuetkU8Fxo+zT3Fe
fOu4Ce1p57AH7dqoENkAup4abH8AMHUl4D/XAedWikBXmMhjM7tQhq0Sog1fptme
z6FfkN8qPy2UG5pne60CslqeTMcFhnEATPzR6l7mJ0Ii5KKjv7k6UaqM9nhMpg12
QJbtVqVh0S0HZTNEe+L+YTz6ht/LAJrplJWxFDuXET/4zaAEcmrl2iH6+8vZ8bQV
D0fOfTbwAmhClVUpai8gvu1QccH6fRGpA+aAY0NDTYn7JovpEsyCY6ko/BLh6s0q
8m26sYfFwc0ZAE1RJ330m290xpu3xl0paoKpvadHs1rqMF9gTRm4vOlA77t7+Kxp
QYlRo5GOZoZ2uz0stUlSlmizM8rBV/pMkcKPrBmfu6QbtIW9aDCMwYnJG7R7+8Vn
faPoy+kzXaHAXiJzir4tuF9ckjc2ON8qtMdVuJ5QOm7EQdqjHRRolA7cKEq4SCxl
ZPjHUXkI1BIk9Llijy/V40B1MQ2j1U3f3aLB3vPudvmg/VoztnZd5GWRSm5pnGY3
RN5TN6rU58dmY+aqofb79oeTKxZiPHOm7ynAHuV2xxNUoRPQQeEz1+v+xHb43+bS
imEgSXR/lvNNlhF0dxzBzB+sCSO98y/v565MfOPYE/QoLuKL47ENKs8WDD97y0lJ
7PZmZF6N2/Je+Ax9fwn46iF+R3EHDRr0wZ6QMo0crOcmDk95AaDjtZ7/qsjTGBjR
Ho9I9kkr3dO5NW4fMuHf2MkF274sZAnClrj6596ImsKoCFFLktK6UdHREBlSj19X
L6LrA82CRhVxXZ0yTFqhxEE5hfq9KnamU9+nIi2k+mdpXfBAe6CKgiY/PYuU+Avt
WmGHwMCv553PHTHZD3owDdcv7i5BTkwq8r3pAZZ5CVD2ShW1/BqVpFMBh3vVjZfq
W7a33llBSBO7xu/YBZDnCkRCcXmg7GIycaml6EBPPtJF19KzaZSA1sl9WdClhXse
GcbXbyDwiDS29by7ZhHgwY8kSQKQr837j8bCpDF1rmyHhxCuJECGXDv5//DOJX7Z
O4KIHDQArDOFIIkArQiEbVBP68SEIxmn8mPDM8aygNtCp2GrYm356srnIC8B1dtZ
og2K3KGEeHaAvpBAUCs01h/oMC0okuX3VAbRPUfCIYqFQ4k3yg//cb4qBUcJ6DHt
ZwGPs2KFSiuO45uG8+2P55l1LrGjKMt4Y8XnAD+vmwqG8ciL0qlyrTepBBgeFZ37
IUqYq6Jnn+dwJv9lHamsafC1J67Q+kRaxQtPzh7/uGLWsjz10146YzOKAp+7kJUL
5PDcU/jCdm2LA5HAi2vyCQehbFOKvJbRwDNvb/8Ubgr9Sf/dLAVDxB5kFUowmI81
A32TLMYBp6GCirLyMhXQio29aFCADYK76JTtEfFtd+OR1MTtnwZXke1wxYaGa7N7
ffY5riW/btxq4wT2B+FE5xU322lz38kAeWP4lxn4c+vGgH4IsG18mLK4GeFFRoSr
3fKBM9inYS0f80wIUSedmu7BwgAR8F+WNN271BZMcACSeZ/g9bEvejl2Ej/Hkn3Y
Q/7Y4WYXA8C63XEl8robbgPCH1zYkOLW8nxvwEt2X/wIVp5YT/UiYiiby/NK80MH
YdSkj/3g16MNPDicnGyvPp+KddcgagczC1cH6tYEBufyjg+FtkT0fea7Srld1r8o
gtcCrJHiS28YyXgyiQULh67ElcKkp7N2c7bANrk+0uXVsNz98Fvv3T1P3vIZ3OQo
Kx358M+6muery6pBg+xA7oSu9HvNOO1bRcn/lFpVnUff7ilMxeHvgNbclNUXqZE9
qzpE8ARFz4DtmVLRVlUDAnigNYO0d4o/9lZUeRZO++vqA4omhWCfSvIOK0AcvyWn
pLlueAjTcdwA6JOcqByhWcOMpZchfJ+YQ2T/gvfK61lhJCogGS5h3IFXr78ks0h9
ADRYvVYwgV7eGRDnoqGp0bzuuQWju4cPj8M7nxT5vzbdsUVNSIZmwmCOE+LxqAQM
Ylshfdv4BoyYwgh2q/ARvBopy7HHY1KS6XIbFyxe32FrlRmkucjOUy+JIXMPkShb
RUG/UdXYFky7sjKFcb9+D6yC5SHhzclv0sSnU5Mh6t+hGeQIgagmLPK1j2uAUDNR
ujsb/Nl7csms0wfWeKjTyPFsrzGMOUe1iZYLXUyz1rSF4ASls+DZzJlwxHTYk+ym
H/vV0zu1mLWTS7p3V8r8YVSUHz/sjTUAK53EE6BvEOOZ0XPG+6U4HunEfFcOI8jn
H6/6zWXGONLL7G43J3trWqpVL2MSFMesHw9rGdF+44gDZoL7BEOOwClZIbA4XSqS
VJMm4ZLeo5rCtJWVdB47u9FuQ2dLxlCbnx/wX8Fljt7ZyE0qBmkO0+jRlc1mxYfd
aoU8jY9rBuqAa9V0xDMGnM3uHdnOKN5dTtHiJpuffncbN8QQZkvxFZrIzkbPO+Bu
XqDOwheSiuLOsKTWs/Om8Ow7UtRmT/jCg41gskdgr1Fptuv8On7vGPCcTZmcKi++
H+qpUpF8RIXC6taOnbQ/Cgi8nVQWvwm/Qs/h0+nhx0FG8VR5ufpItBP0cZMA5nY4
K1dxi5xuuhxmsEVkdZAyOAyW1P1zRij5noE2Ya8SLZbIEWxu+/QHk2enQdSZWkuK
DcS1QOE6VL6lb/pceHZ30uxhxfI0DHkM+eTfantp1OlUyKj3lQBfkL9OI9jJ5fDh
FLjk9ZBtLVmNSfscq/8jki9gWf3MsbFYNbI8xIuzX79MV4oNt6N9dpX7+AJXzCbi
hdS/8CQXH0plTRYw4sobM97cRduHfMzDluPpqZvOOehLYpi00+rznUEmCl9RKuQk
Vq3mfa5XNwX2y1ljni5Ggb0y4XBlpcOOx0DmXQ8vBMbE25koAmIUfbwEZdifQ/re
VSp2eib1VdcIfG/A19CF+ePsF07kIFXyF61kZGYD6k5lFNTM+3Zak9hBLYCgKm6B
eyr1hyPyGQkuTFsfdhuvr+ih00GqD7wol5fVWpEwUeVhHSjYSlyeIn9ykoPKuyfK
ZmETfoyGbs0X9l3Ys8ZwnlKNOKKvG/FgnE2s+r3ZA3FDB3dyKhq4mjt7BKeNGR5s
n9UPhx2i2qvlbh4m/Ds5AjtNW0DACpKKcJ+DqWhVanKGCJw39rh8kU38Nb1Zx34F
6eSiUrlYwXjtZ9K46bkHmddA0zNwMOJ9C004jcvci95HPBUj4TDzRQIYIKeRNdj+
7apbOHsir6oLrNh1EqsDaIzBbeCvp6BViZQ29fmb2vVbCQqAgLkJekJRxZt8PtPO
Em/3Zj8aMZQTN5H4EkZpmUjTHdjYUkVqhYVx8lfVF72vUOPUecTrQMEixwBHVd9s
B14SiFtvcMfSiinLq8k7QfUbTIBoRQpqO5HwEpc0Dw/aiEY2muhE7rg9/dbkEmuB
5fI6w+cJWGa6GUCrxzb+XRsWQ8AJkLbuFZFvLn3dS0vNJxX5bOCq0x/cK0XNeIur
yuJWwDZ6LGDs3o4vmrbZmKIbWz8ia9n+k+5j3oNgje5HuuT2cyO5+qulhNga5Ghk
jzPFZDWv6XgD7QrFTcS7uioArajGVdUB99F5RGQkNyU+ncDidP2VXvf8v7TkBd8B
QUAxFkX2GJGwx6cFoQXH9SrigD+pLkfOjEiLG8kLh4P5Ct7/jXxitDHkakgVGLX6
VUj81hXHZDfoUzsRVzn4qPcr3+PEE6zuVj3ozW662ByuNKA6rUJTILsHCUcRWkJz
HxOMlHiiXU1Nckhs+pIDZ05TvlvvsXS8Qv6Si255Wx1kvK8i5YG30uwrpyOjKpe7
FbSPyVCPUuoB5w19KnJi1/viYqRHITAXHVRyhY4pbPD/KwWDtzZznhJeUOLZyweT
2wZVLdF33w9XC6V/DRl32OatSrKpCLOjvtlPTzig/OByiXjmZj3FGQyNYo/pR8bt
wEAs+X2ChQVsQ0dTLVq5hCuHKWlCypX1eiOssDW/HY8jYx9oksxdcWJuJ9RkgZ2N
Efg0b0oXrpruatG4ZBy5ESirZQI5+fwWIzPF8r3jFwDfSKZ22rA/4uKh8YyWFRRv
A1rGZZaexmddaKkIuXtPaW1Oak4HgG+3VjUaW++TzMK+q1TaflCZh7w5xo2QexDb
aCDxMyzDQAZPRuJzGUfVryFJsXw8/wXjlhdII0c9HYVeIyr5vqa/UamcJ+GV8jdH
esfSKkYdAfF/clZ63NjeCSOYhbt9pyE2xh2mJL9GVb/nlpNm8UITE0xUtMHhaUqb
nUBsXJIp5Sx68t93zob4BDjWdFGLPUg2Snh0/efAoirRzZTz0ggnHNjXdr6J897X
QBOt2y5vld1I9Tict4rm4gNoyBQlzbOlVPSVCFMAkJ2Gx7/XISZvh+kFSa43pER8
0podBja6yU1jvCeRe/27+vAeCgzE5Gd+HkuSrmbmlmfiNd1zTOVGtMPMYSimre7P
Xoeqfr9CBcNKFc1Ac3bzIYaxbKF361uilsQwzfwrzq8isd8qtweHIG1Al8L1UDVH
2cR3uPO5b6KW4o891wygY4xAB2xxy4ucEZJM/PjHFqix7mKwhKDqCqUWHYEPcFt0
xWCwRJ4En9pnlJUY6C34aNELa/BJDBGEVp97VJxbJ3Thf1jHphTRDjDOrPwDKnPZ
uYdo/qY+9RQ9L5g5slOIL+c8BH3ORelQPry39XYi6h0lwl93hOYdptp5ii9xvX1X
g7NWlQMjMm3adeRo4+OErjQvIqqLILDnE4e8F7YV9vKuybBIgn+RmZc4o+rRMHxy
hB885p1x7xq54aU3qYwgCQgogqIE3lChGWWyYJXwA9H/OoRopZisxNf5nUEA8z6R
lg80537CPPd1WAVJth/MYQUqQfXaV0Lcl+473DzAFbSK6VC+ny6+nZTybatHvxkn
ZS1doktbeZ4pg2+Q1KmtaKEEIAPv8RwWXGIy+BFERgw4lY+7fKJ5jlVRry0PEllE
Y2Ui7ytKnlipVH+FL7rsBmnvUCMjPD9FolLj+m/S5l2PZxOGkCKMRgRVvH95y9hf
yWpudMdY0L5OH2EOIXWFBr7U+GNuu2318flG/Z6AiAr4TjEiW/I7q+oNodjoefvZ
HCwkO/zn0vjallT7GxQNGtsixUILLuW3tH4H2CpzJ7ASClFqMaolizfYUGYoCAeW
7bzJV2hIa5a0zxdXuUozjZJRNuDGizhQVfM0DOVuihh5vink4pLy8+bnrzZ3Q+uw
kO9mTX5ZGW++0nPk0JIVGTSfioX+ZeP1cwbJm9eGWgcW57sL7c1rp34KmoxwOe4y
qsaxDQPhkaQAZE1rvnursT3fB0SVX6gqE0FtEqFjJnAfMcXDeSElkStldEK1q91K
ZDdS0uSMEa8VlK+ABH1Ufb6VmEMpMQUG+O0DlDGm6Qwe74k6l7ZhQxpqTSqMY+nC
sk5Yr9KiYf5Yt32Q6n6vd2GQ+Aw7Br/pCJdHZXGAlngnLhXOyykOH5qJlz6L0aaB
ZofI/y2BIudMZiUvxvk4p/SUppV4lmtnUpUb5NDM+Nf6CLpIRiV+81b72SaHEPGX
sz8UgMGLHAlNB12Yvne9nwIsjDsO1/f9bNDYqrAks1cI4BeoPsxmA7DHGyOA+8o3
8Ekb45auF4AU46HjZfcKA8anOLfTJpUcQV/pHZBHFs+jg1fUhwMDuEBoDTGPBbz9
lgAkMTufk/Vqmr4AdfA6O2c1MrmGd69r3V/9ue1lb+4ML3x9r4ig81ifsuv+0yPM
GN8pU9CBMovbTpS7eT8i4ol+buYKw8emp8Kv7r5B+T+Muw/Y+tEILez/6dbEi3Zw
xkdRkgleE/V1Utif0elhrkYBsVk9MczdxCNOG+eBKCiIVm041h+a6Sm5vBScvub7
pA0NzTYWzK9NJySbYtaiDtmZuQwgzkiWLAY85er2KuNovsldmO65I25mgZRUzqZ5
l0lt5pAxJIwaDGtI434EVoo4XqFi6zbPgO+jizzSlUvGYaEPK6ORzx2VxtC4+b6S
DvjklT6l/eEI8wm6OskjoILoy5Acdg+ed9NOyg9DmKgBLsPXKQ0ppwVBDje3+zdW
pCu3F7kuOpMDwYB/1Zyatn32GsPlu6/u8X2zr2RwQOqtC1ATuwUpGBqNU4y9XL0W
PSsFw32p5ffKUti9gQ7SisG3T9JX1B74r3AxWFZhJ1GSWI6jXvigDk35zgz1Rflj
hjbVzl2dXKYtwWMITmB3h28rundJDX6q+3Gd9C4gv1q/gOK0MBDSSzC4BtJPbgij
2XdZlXBtKnxW94kaWD7zSs19AZprGS87S7FSS7IJi+2OLjbvsQtk6fpeuixqOZNn
042f/gCgxVolTUlVQ+PopmhCcg6A46l5wbE5LoCWzCwiwqdqZg7uU+U6QNK88EoG
Mxb81dfaASU+6bdC3d9DLRY2yj6UUhAeIamswZaakyJ0YQv4YTaW319ehWHJDOya
BH8Y+Q24Gqwf5/ZLHRJ01kKoXtQo92U6R7/ra2UqRwlt4FcHQEsyoZGBqRwIlhHI
aRS17djRqtACRFdPTBwaX6Vu7q6Udh4YMmO2n8u6ch7jVmtGDgKR6NWI/90ukXMH
QBalVAF1xH8lQZMlrbbYIn+rcgseMi+v6aYk+qYOiSiRFMvqo8UcaHmwLaE1V816
ccyzONNtwhEPbON7jGLacDwM/3gSrJ2ROJN7ASl4+NOorCvCj1uAtvQVcp0TgqMR
2FsrGN1RE2hwFotJVWLS7lh7k0n0CPAM7jAPXI8w8WCiGx1PM65Ftqa6s9m461+2
GmcuNvs3c6Dx3NpmwFfabzRi4+pCgFu2GFn/PdhfVaaGCgEK5sYDcZe0CtXmBmmR
R0AiLdL9fb1IPCDJwqc+gcqza2D46dKBabalg7UJZYMtta/jVzx+noDiv1wS8a1H
dWevvNg3Z172mj4QmCAsOmbl9IQK5Bir+vbACymzVpujM6LJNPZoZGFbJSTd6aOC
B9CBowCDcx836qBWzPDYDdlEWSkD+XCYuml08G1owgURJYZzoW6FNn1vmoS1Gp2U
OmYosLFCKE8y1nAP3rUBh9W6YTQVBphCkTyWgmVaNTNuRJEkLGlbAEM7jVpCyDdC
0BoA/VO1slFTDtJ0BXzVrNjDEf2fDhf1yrJbuLKwr/PjUocgxoc0Gfl+UE3z1adu
1G2flrbTV/GTMY7LlxP6dr4X7qoY+vLuJHyUdJ5m+8FTeZpOtDBwwa4k0W8lQJP1
s9NioBaIYjIXn8pf49wt9lif45zab/hNVI4a0PjEEWKFMrJ0eiIQfetMjYov/vx+
KGC0jtOdJOLKmXUsk2C6U2s3jbG1ry/JH1fSWTlpbi+Ke+AoxiHc32yYFL1CnDhZ
r7YGEHXXb2XUgPE9PpPCi61w65ruRblYfyDs9BRnyCtf+hjHQsRj7B6EnW8OHUvI
HNAmjZbFLBT6KNhEodYVw+rdYNwDiWLwt8qSPzNOtmE6JOLkyRxjH8HlabMvojuA
NeZI1NahaKzoC4epYfpx6VQMubBh8Hm/8G29vtwcTLb1mHFAJx9IbQtuA8U1+iof
7ImHGc6UafEPR+p/+IS3mKJc+mHx9u6IiFzWclTlGGHWcR1+wLBnWwZUAru9u/KW
zU6+YeamJ4b0t6axJwgRwAbg2RrCdn3ZJRJeH5zWGGc83mKLvxEFR2cSMswq4PZv
DniSs/WA0LHpq+LbY4tWJcZRcXAA/MaafZuvX1DXQ1uDkZMg1JjXDqsx3Emg3Dxt
uYbLCWqvLuBj64wCYTkRfsZ0whH+gnjgG0DThYf49rqxy8BZMC6giGHbgZFc+Hg5
XPsx7c+T6sXcAHCNwe9SoSihVv3tiUlsVUl0DA1bXAlFlg0mOa5xcVIB0f5AA+mo
uNAfYIAeKo728KzEIfYQZ2dd8Khij6xUlHtBGe/qpCm/xpczweq34guwsQihzAP2
zepkp8YZfGzDVxsAIX+1SgPMGYLWnSSVN3RfhhTggshFju4eQcHW1oSWNcxjv/nn
JT9JtEVDwmJXOWCfUmkslhD7McuXyCUO03BHXz4JJPFsVfHqisHIBe2TAkAAeup6
+OPulMTn3xeiFS6tLfbs1ScnAJvqGb/2lPF1Q4cHa5nrM/w3gg3KoOhGwqPQRHST
XmQjnP5U0ItWm6iuSlhGIvnzS6Xs1BAnxzXFAlOdtSuqcp31/Jx7MtwPjF66wxsh
b2oNk7RQr1ea+4FtC0cI1FG2tSPt/5hgWNmP62yz0TWkoH50X25+mCNXbOEYx11X
1LBJRcNBCgxaHj/qCbLzkQFNcPSTBONfgg3DsMFafYvtHg8h1FmVXZRgIlOPiuJU
s8YIbOTQW4mdtHObz8VOHH+qljU2Uc7OiNS3rDJkWkyYH1l2LqxsneYez1wnSHrc
uGQ7L1rSzl18dQB2XSVFMdZnbBDaGZey+u9yEUrPBTT8nL5BM2VJRryEt4YevsTx
mDJyMGIGaFwnyd/Rla6O94gichxn7ul15w4CpfJwPpwX0DrQ1d2F760HPJ0diHf1
oJTY3uVLHbuAWxtq2/ynlm7V3slXggaRYgbgLZ6UKIYUuPTIRXHyEPlhky04AR8n
CoVKDLBofJP2thG4JSufN8ubGB9bNtFoarrSoF3MsjMrw9ZPe4wIbop3199yUYGB
qQhyo0yxoraekFUZU7RXUf6FMn6Fq4xoHJNVutDQPMukHAEBz2GFPRYsuh49SaFX
ZtzByfLNwPwT2o7/w3BF09vmjOXAgfcre7ohK/A6kwDmUxBdvU3AKEYuOVRkWxDT
fL6fp719QYDexdbpfW6T1ZBhPzsUuuxjPnwjLfz3cAdwHgXZd8qx8CYIM9h97zM8
qLMQgDD7T7WdHsxbyk6DaWEgOIetxOPXALWMVU4w7M7+38Wn8E7E0UrcC3wv6iIt
1Xd5hwVHZWqzkal+kaaHnQarduM6l93bQtqjTbGLUVlrgulkOmUt8FTM172WO+jb
FWkoY/T0jnuusDT4tzea6xnTDGiCzbpStHwF99UwyDsTI3mYSISyQE8MxWhTEllL
64oCDVeNOb7hPp78pUdPsL9aGqaDTA6pyjRKMyq8qgJt3LRz/dnK1IEafgfKYdqb
oLf5R8cFMWc2INYTIOe9LEfj3kfK+GM1tJAB02G/QM77LPfDRPRX6T63XrGK9JHR
r1aFko0Xp5zABkg6viJS3ZP6mZe2xHUrHkVhknUsadpZbmkYCi1bLw41UT+2qk/o
/HIcvwVMMsQibRNP+uVC0MNAsU6bj8WKwrbOY6MBn0JXSLmQqrPMjLroT/mG3IvU
FJUd06Tg0vnMDZAY6PQD1b1gs6tE0UwJIBt/9p9WpcvGBe1EQuungx6TydQVjJ4c
8LurQVdu7SZGSLfUCeANRb6GiYd6OkuSnEXTn1xGY+A2kGADyTRH1qpjH3kNEvYM
vF5oGEXWRQ3BDwfRIII7rvFZk2paVfP1eE5/CHWikYxCSRY6vsPGWK9QEhYjjrc2
cCUAt1FMD/XajgzWdujy/0L9IgLGcbOCWHNyYOf4RPmneKsfJquzQ7son43TBx63
0HsSGyAMloNDIthyyzFdj0si7+yxfPivWrLr0nerDrtRK1omQV2T+TPr+tWK3V4B
DstF5zcusOPW1d8pJwug9n+9/RddEdjAPJGpFJ1JVmDI8itjsaYs/ToVz1oI1mI9
CraZCGnf1ckM7c7/l1CmWLvS3ld8Y+aiIP1fslaW1qHjLhX0jNsEL0R+51SMWESP
NIzbbbSwhhyQXvW3Gt+4GhhXY9QVXfEznHvPJn5VVXeztYGoJSdnesnr+6QrzZXe
BHcAMx95db3IIjFStVgZEnappslnozN453LsJr83YU5M9gyC+2/kwcxn/ZZwuphq
AgjIeYOqEJeOZY7jXLGL8xZ1LnjIkaDOuYHlVBvjLKN1NzJKnwnDUnRz6tHLuDkD
NoMxK2dJwMeBFKqN9K2H2e9ikUG/fny1dZ/1gOHHmJ3ikkP3VO2C2bsvquWHOpJ8
kL7rNXhKOzoidHufWIe3eFFtngZCa+yWSFn7grl/QmOWEBaqx5lREtvZP9QPmK1T
T0V9pQjeoxxRfSa7OyLASWvaCLfqrHBUI19JL2FWuD5aILTDIFjogca7bZTkdWuO
Xv+iiv6GY0DjX97Lz5hOPfyYxFcrKZrZwgypyVRmnqBTR3n5ZUV8Ki/VM/LJFcU7
DU6QarDpleX/EwB+CCA97khLbi3uXB/9XqYicwwvg6ko8Pvgz6VOTvBdhoHXV9xS
0zk6gwQmiXdrBVpoZqAlo1oKsaiH7CozpxZOTZ1ssdP2DVoHg/Wtbt9a5plnNH6x
SwHOHKoIKwLhW2BBF74Fx0yJ5bJKzas/lHHrQGD7TfIoJ8Zp/I/GjUZ0m20AaRC3
xM1hajYEoQOcgcf/eMUPwfxSljBOiyCGqdkTmiUX8o8d/5gNbpZeo4pCiuwIo03X
MLHWKAKHpJDRmXs6aTS1Xd1E4sy8xHjFthI2QHLIlsyEX1WP+XrshWb7ggAt5Qob
MY3FAJwfwVeDiR5kF8Tk5jXId8kHilSEo0v3ACq2aJiGgYuNReT4l+Q1G/FAwUY0
ZdvrMfOM6VcfsKX67DslUG/fMieAbqcRUjMpNJER8Sld5q8/HC57LUECklLjQLtK
9zdZDMqPO13D3yec6SbluLerh1HRNq40L1fhifzIKg6U2h9/o1o1AXsHF2uV5B2E
WT2sxxuyib0FEZmYhRLJlmcCVz/QkRtBuP3QqGBgqAuABiodYdkndhTdhtjgsvPV
qqTLoES9SgHd5RMU/IK+MXUy9eASuqTbBFqfpTtKyG+Vq7hA17QY0Mgmh/evOZAz
qaAB9hZqvQLc+2RoncbM23wvR7h7Q8i9vd/eg023b0EluVDrR97xaAmNAu0nEaWd
8Mwp7H+/cBo9BIu6oQrWD38IXXNwJR3tZi1H4EIJjDfKrBPdj0KevxHhRozP3HnP
elApglebEnWPYHlVmkooWm04uc6s5Ko+YJilDG0ZHbQg6e/04tOhGWqKr8rH/Y7E
NwWeWTgEb6A9lWmdxiXZpUf5ciZStZLG1g4cQ34u/vFFQzumGETTUVXk/sjNFZ8+
oscYvh+MHh/aEQD8GoTmUhFKNcsOilp5axtZzfQOboC+R45WvWeixKM+eTc67LDD
IdvCGIlv21tuBtJEByTxbYDrGx8KdwfLGjxW1/xwp1oToJRnmrOJuaQvwsQwVGpw
9+pBOL5jSsgyg6Wo4CTDbk4ruOKT9C2qdKaA5c7f2bb7IH5BBhsTrJvyjEZa9njU
hqQNI661/dOixOkPU+y7wjBu8dvywgPF1TejWEFCXhbKIcwytCK/sPWRIjs78x3c
50EVwN+ZrhKpHQr+C9uz7aL/aXlQDdpSumdtfWYDRmvIH68ShDeQ3Pkgr5MW7les
Pifjvhh9qubArxS7dLE03AFQERWlKxExj2sVcUPEMFlwFi0C4y6HhW4k8LpwOuZj
44oCvGVn+Jfo1t1h4QGTrh/GHnwRt4s+MTqkgHY/sRRpXpzbFBx4IE+a790cG1my
tw0ifVK7pL48gc9oxkyDDob/3hGosM6e9Yn4hp/ewlaF1JhzhyRCrExmAr598Vh1
V6GTnsBwVJslStPzrJuBKb21JOgl2fQl0Z8QGbEVTh1I0ABSPKGm672XFM0Vc+yJ
uqKD5CwFUymPq++j/GTEf4Wihg7N08ZxmOYrr2hombFUwU+KT5dJppD88si0fDBW
NtJuM6cquKjcWhnFseQagSHOvn8vdE9IahAlZCUNSIBV8RLYiuvlOiH5mDk2jwCn
fK9gPJVJCxlDkUbUOHbollfqWyDNxVxP9DBT2kDm/KNlxvCHjjYyBplmX+6hO0R/
9VtvuUFar3KgEowkpiukI7qG/f54hXsBecehfYpHGl16t+r50tn2D59eDg+EETnT
4DbwWXl38E79MDqr8r8HQR9e0bDgO8Zhfwd0cgtaelsXo0e1clCavd++AQrsbz91
WDLEbL0Cdqhrgd1wcvMEAT88V//v2ILPm0HqQD+pj0/ROXLU27aVeGUmTWEUY+FR
Vocni8kUmB51iXWtsYQArgXrC8FrfTc7jnV7qmNdDV7dgJI7ka3Dxsi7162rbTK2
IjZA+GIAzrTu3xh+2iw2K5Idvtswmk0njB85Dg/Usi836tHl6WcxrndQYwDStcam
VSiPMEBEWEKgxPGwMQFNbcu9RQHnTgDYO1fRISFZAneVcNWtothoY/LUAXiSqmi+
fi2GWZs6gWxXo/oGN07VlgGvaFcKhipdQqRXtkGGr4mLk7UcLTjBhQcQ+c8Mv5++
tJMRN/UzK49WTvgPuSuKa99NjTmBvPUGECTVatWC8o1YIkcFJy3pZjMsgTkPVzpv
8Am4kho3aZeCPukVLRQA/MJT8vsU24QVSOLDi1uDRSRunBCEXCuMDWAfBuX07t1D
+yeOHuaVTeNGJ3a5kbu9pqZY1QbkdNC2GsHT2WexVzMS84PFY7eE2MREW5PW74Hc
vjSVZMB2PTqD1K6Z8hsZpI5GVIzXzmb8ljFMwjKHWn2WY3F4veBp+wKLYKC4A5Y6
2sqGVaKp5j8Wl57fv7pEdhE1XeF6Phhg82V1W+JFHvUxEGdOEQ2GdFcArc+yn0+2
cNVotkmmuhYJn0Px/mKtUP7s4iEUp9IaRUUJ3hCxO8PhLzUg5V+a3KIfiZYyqVMo
OhhLPN2aUbvHDMe4u0LBl8Bj6nq5xI7m4LZpRcJEoymo6iSX9JU9knN0gr0XelBV
H1em1/1qm8zStVbOvRL+jDM7Mvk/RRUFE4XFryBd2AMuBE+tX6v7miwCZYF9KG0c
sejKfKhkNG/VhNRWbmDExDV9esgPrDwXHs+c3peEQsNmixeyOYpK7hufDFFFO5/v
weLsGSiLu9ZaFFk3UPmX2hE5ZzEzXGZHv2pcUSn93KRHIVYmLaX1kHvIgbJt1BGO
ngw1dinUoq49TR1Lt5zNJmYfZlrNrQR7ra3yR5WKub/9IKocTUWPlJ5lh3iBOMRn
tFUO29dFdBDwMQObSnAkqxLBmis4wkUu/KzIc1PrG3iIditSbdziZ21Y+ejye933
vwpXI0NtRNslTyWii2hWwQo6moO0Ob29wfMN4hgGm5c8Aze9ZtdFe29fXsq28/5D
LS4QaqK13aatLzzd52YDIezj5QrjJ9fJ12aSN+r+oGWMd8YlkNro6RAc17oS3MB3
5fVtbDK65ODaYkPA3GvdOKK/Krv+Bknm1Zpw33I76HJ/8HiMMDgy1GGVYhnr56AG
srG3x0h7JtScNptSEqxNI7lEbZZxovqrkmiy/gli73t3Q/plKUxXiIkV7ltGJJcu
gwauUKi6F1U1HSg99B+UbatHFgicJNYnHSU9sigHXMS/sTTDaSKfZasDGySy+Lk0
VnGMMdGtrJ2ZPkkr2vaAH+7tZwORo7Rid/21AQ1+tRcXlSkuHo7Y/OdxHTG05u52
ca24iRSYZn0SmwgpZcimhPiJxAVn9nQkAOwcxJMXFmrWsOEWeog4455NB3Y8+san
TD9U+kJycjazCe2+gVguuvBAbtN2GuwQ4wmtfvCCriRRaTkR9lFhxBDnr8lVB7x2
sMtObgKMjpb5EIwtjgtEjrtYy45H3nSgEk1DuyF/Uu5U3PLXc+dOgTvMk5ObTMpd
knyhkrGxr6vbn2oMY2yBKqnI8plFCCV9X8MB/vVSLghww7hkFNokmnzYnyrASb6L
JFVlFeCDm/aMIb5HjQ1fRT0E36iSWnMcORCjzy4+o5u/w0FBV2SohhhNbyTlYfhX
LW3Ml4iwbrUbcfmKyo5hFWoNpzZVQx2RcDFVqzGHhzKmgb/XhqOkoUF8b0NfeQTh
8TiXTSIPC8ZX03sUyw8/ZZ+onMO4hsIteBAas7ye81A4KvJT1dwha3zuqL7UFVoB
R0BZx44ezONergO4mSnCPv0UIwnEmWIOY/fXMOl7gYJCqrNLqstVq+5qEy3bYGI0
LlO+7mpEz8TZs2ahbpzsXNWldK7ralaKyp/hmUklNqNC0AINitABjWedDYIlOW+K
e9PXy/znVV2HJ7sbBcgJzAJtVRXpzP6lHABH9u9bTpEYde/QGAjzr8+dQhki+OA4
6KFoC2ZvIvGDb5FFa3XkWKFERTmNiEgCr4T+uaok4vx/DLPwggizgBlAp68DMdKv
4sNT/orrZ+7WyinUNsSbU8pjhFp1NudTSxOAsO58ni3XuRpQVtYMEICenDVKozb7
ysM5Pb5V66kqZ0d+ByYMN89gWONYi5QqK5vncQ/30G4V5BaGQoyaYNQY8caWzYrP
nfHg5QoxrhyGXmW+7cilFzbVWcHt+arWkZA8pxcD36DuiLE0VQD9lhg/J8QFpOna
SDCF9WTAQFfWUVMPcKsKlwqa87Z1wgoZ4hjBsFU+LIkmLuvaebr/XahG2U/uE7T3
sNnrTBo3+PZ5gYYyRxx4CbLkQxDrp+4UlV+hqMyL7J6x1Y1bPqrAi+LnZS+Al55O
CZ8cpB1fPeFYJtspFLP8JMGUcsQhCEZOr/fNfoeELx0Yw1Xh6KCK8Nshah8/vCrT
BHG7eqEbgItJIuuuJCYgELifBA8ugq2Ir1ha9oQtrphghMpPgH/T7kNajpjX8tdT
X7/PCBcTJRo54t5cveuayTrwnygvxARp6QAqz3QHi5R1g2mYJuxM/r/KbcNlGAWS
yAl/KXS9QZSoZb2VpZrVYFDKlhDyt97ULrh2K4Ztn8Fp6JHeCdyx0JrgBiotb27F
zkXuPG2XZIaHTE8C8T6fKQGpCbehhC9lzUnkJxsYvFKLPbxHVIaOGcuycVSTYfoH
eHPixw0pUDvQc/yMNVMA1KWmYJjcCynXr8vLrGbZ7i8wBAfAhaW99ryK24m13Ik2
y954Fdmz66vO4/MbjrcYJjzsAUoIWgTUJBCCWrnTKKpr8Sh1fJRLPrOp+XOYSRKH
2bC4bjTUgDB9eU7fVkjuza/NhrVDTqZe/W14qhnBHAAp82sy/s7zzuQpGBRIpZ7L
aMgaMmDjAoa7eMOMHqSUXMPgMLAzy9stX3h3cth64YTQ5MGAkb995/j8NV1cOnb+
uRqi4p8bIe2z4GRVeK62WgGR4DFmdYJqB+E1oXsBgUfHluBQPwbXcnwK5VzzuhyK
oPO4XWK2nL0Mfzew1z+k8RoN3fmzl57dAvNkxmuEVoXYe/KeW4lkFP7mCAXjg756
jwc4aGoyj4NmcBC94BQ2d//3f4UNPEwz2fcgq69vWk0Xpr3a+shb/goHu7vFdoe5
0IRHu5uf29e9OdICol+MNbMTzDzN1+58PaIG9CjjD/izhPigvmGswprX7nyuppxj
6Yq4RXFsUF4vrpDUiSsW2QiZAs9RnEjXx+Gi07F4D2N+Yn3OE6yonLsKPQDa2Sti
YZBMeETdsvLlNlxXQWoBAgdvVkQWyXULPOfjn8jhb9y47wXtknt6ACN2xTPAqAQW
200uIoHB3W7QMgE9R8zsRO0GwWGqv6FrMni+wEE6o0oAXbWokzVs7+k885aSfjci
B/YBodSntMdxRTYsZnjqRq/HzJMWcfuz59TWr217uLBc0mnz8n7QvrifkdsYwfIT
yETSADmBinehU3GsPxNLfg1z1NadgxfSSanSkicYfA07wGXyF3PXF/68OrwBnNkq
69YSMUkGMZoCm8tA1fuzSfWjfv308M2JMFISKY5kUe4CILT4bVVTuA4U8t9mns1J
+vsrZpJFS5FDVZ48LvpCps/KuZpFtf8WYghL9DU0xDz5E1KdRmeACaa6pDqJuDVv
iJRc6ZE41OlwbJT/1DYUV7Yn06WIcwBeckgL22ZIYzxvHOr3X8pToj9wb/osdjXp
17bj6rz2X+46qXkVqxGvQjtOCBCUOuSwt9Y7lPBRSb/0ujiUTU5d+NHWvIkVwmgR
ItrMsF4r6I38iG7hjTAoafMuKA4biXFzuTEv6h6ipfb7ADPtKlshoTr1tpCcKsZV
VxYQzw+LCQgr4rJU2ukJQIIqdp5mH87kgeXa3njxoh0Sj+qJOaOJ1izUbzwNDDRU
rmyEUvpGdWDOKhcPnbR615w7Js2aUghZ+NNF2zJ02KNhYJBQuDiZNgLtawdBV1gh
Cj77iFYppiOiX+8AK8Ib2p2WCKm/zBuxKYT7yJSA3/tEa+tRaEQa+hFYcCUqnhMA
M9Fe+nX65D2PG3X3IqLKbRuCDkZkGiCGV3N41Wd0Fn1PixZcbvcdTkLi4zi0fSdc
pc55XhebIWPfN0M7qM6rEIPyvCFwUU+E66rrLDd1G2qWqzgRb2QNefkXE9facydg
CpWB4iWaGG54E0MGHsRz+1XuYgx2oBXgKIl0zTyQkQkNsD4byCBBwK2YJI56C18U
4Dm5+s9oMTP/p5gx0VCkuFTNfFrZWFgKQWyUc4JwD/+6oLALfr388jlL3IIvBgKd
iCB9jPqHBKQsvgSovuDSspX+979qTW5kAO+CJfJQMDkE1KN7iuMP0HyiM3/XLJ6z
0fGfdduMV45a7W4GfqfTN3O6Y/x8rkW2vx32/eeNVClrqqvP6sbEktf6MBND5rCq
9ukP2c/Er11BeX76MOYv50O5npaPULz379vfcCko3i10nud9hS34GYqG9ZbACEIy
mv4UFHW2uMsAmQ7pnDxKcb9yBopyA2en4WXfzR9HsO/cAHlKoghezFsBLImRlmPe
YT9vMMolYCkIwnER3CGGavZaV0vldQAT6GhTJNe1I/k1htUvpcnT3s+wYKpmtnhI
12Hy0AiUIeF0mjioSr2VydHs+wUP4STrGRuMnxO/6OxlPPT4F6403FAVDBNFwDye
y+hIqMPEKPSsEtce3b/kcUwhxxkiBHgDLS1jQvT2mbyQJtsrOpNivqdZMs/TzDGI
+aG6FZYM2XOtyYEqntYyiODwvhnLTZL7tuC5fnrMZtx3dQeT1+YoDULqZexAlGZ0
IWjZAigoZI1k5mPn03i8xwrVVb0hXDfg+vJD16lEnKLK5JrKqM0PtlofaQwiTZ0s
0GLjOytSwaXUpiyCg9wpAyHWHJKH4HzbJiH2vbmBdJeaUR2zdTNxYGBd3bZljehH
FeWN4f+2HOgUO0e5x7YvpYZZCKj2aMG/EqFQ+UqxzGLz9PfZr41rn9P2hL99YSx6
QhH4AkacnsLSOgxUGUvkr/Tlyec5rEOg0htQUDm2T4Awh0MzgM8UYiwIUU30YsPv
XFeJmQWCCiJw+LvQRfb2QBzRtKAU5AqZnWaSJOpld3TZS6oiO1ae0fM9nOe5aB6u
e24MwoaQ2G6Sux1TKJcACXkXtoroZDP3q9lb68FRGefYUnNhoJHTA/TgxW06Nfvg
7SR5yaarxczgbcj/RVa5TxXSIh1M6g3kSB5F6j9FSKB/B27mOL89Kb6mFGvTtVeY
0C5RJu/daGUcMdEiZi/W44iPZH2u6cFW27shTB1KKIHeCOna+JZ+yRkibgFe7xDJ
2TpW/duqRJLBNE9bPsqMKqfAHOtfC0rbUETHASpS0xZFMnECMLkype3scNuEdKUP
oeN1b9cQPXo7SVnHLrna2njIGTMU+AeTzZ24yccxsud8frYI+zHNNGN2gVSh8uW/
c0+4eAH52N1EuywxQ2KOPP399c9QbXXOMyH9BChIW59ZCNWzxUk3LxsgNfwJKjao
df3M/tOn8cKG4399P2sXEozwCHGk2h/uNvILOPvLpoNpZfxvxApJk+mE2SXLdE5n
biCl4WyhmWxHi3qGdm8ULJ9N1U8FxB5mf8CVDZRElm1Wqsc9vDgY6lz+gZmRjmAB
ObQ9v8RRKJHCKjrX3gRXrK3I6PVaAdi7DuqcTulrDphZBh/pSxKao1/OI32x0pJc
wCCI+Fy2VcV2rYOPQRbJGg0MYsLsKjUDjQte2DBfg6ax0dicuHbzYoWUqQuGJxTs
nNzxDxFSblTKPLwf1UOQSfOjhlhwLQv2PTNM41Er8EwOK5O+0qN+63urw7/vd6H1
oqVyZbWdJrT5xCH+5UqyaAD8rvirvjz6tuJW2ZWcKS8h9hnS3yu2UhXWkPDJcSEo
YH7pECQsTg3V57k4CbdV+y2L2M7UsrKRPWhj3fxkJB+hHZJp9knIIwaSWEz4EKXl
hxiY3qPlGoMRuapafdMl+EAIhw/kFvqqH8Ng6yu03W3gVBnrYshhg3ws/6X+nsrE
k306nhXcQaCJiQuoruSSALfc7qwTf7tWE7oqubYhvME4V7AaBgNAEcyN+9a2eAmh
Gy/D4V0UNXPR1Bwi8704/SpwpuQMR99LAtnTBvsNMBbamC/ZHMiQbgKz4vNJQ1wz
tqh24kyzKz1OL5z0vJHwCV5kLRwXf0CJDsppP4RtuYG86CWBLMVFwUksVNw5gJkb
w5aE9NZg32Woms5fible2hnAWvLgR5rZac6RwucBBXOJ3j3CtosYbZZunsUZZkbx
kP6fBrC7OmOwEpSQQLppoySQEZJa0BQ+CTb3Cjz6S7uhLkCOVw3QRuODtMre1BS8
15rutAif3cBlDkc7qNFHY4f9AVDvQwNHMxh8VdpVj+xzlfogFnwk3vO/xV9mB/F2
5GQQygFFLkANZFqyzW56WTcPMK43/MoQB5Wi7WvRtnYUUVMcNZ8ukyZmFLBF24rj
cK5bQ8v/1zgzDF2agasx5hX26ls7QfYkRPowzdYca8Nl4aUGcQutNE+hMQyayOw9
ZOpzzyYtL85Wm1zzz5dk7eIx45KfRxRgunM+39HhgBnYRGPdw4drHHfH+Oy5u1YK
cvfOR1eaHAeDGcZia8i5ketL2aptbxdDezpi9J67gLcYA1t/x38PeXpsE4S8yeF8
suAm7P7ciZ4YCuo0IrQlX6Q69hDfz8VcJl/Ut+6GVTFjg+yX7mllHnHNbuQNpkRK
EQCWlPhCyN6ALyBzx1Sw1tv5y6ZI349QR1rkmwMo8oiI1fAMLYIEztC3N90RWPej
ZGooP5p5PV4Dmt/C6JBnKwm+LMq5zZQyHdxqzEwt17ThMlKGge54vDjqUXjpR8Fk
cRRCCPrEDZob7axJqB+/gCupeXR83w1uy1YC7AxEkC8wE4cv7ob4i3wYABrqugnN
rtqRNBXQ68MJP25mUa4uGNKp/nAW07vi2+5cU8DSqWB5l7JlwvFNzVNd4MKZVS5c
nGcLSRSAs2TT7oSgExd5eAtcK0wUc+TKk2BLDW9xVlnqW4wyx5CQ0kAC+R6FQ/gw
5Y1xonBFopFZ9Niw5hc8t+fyYsqSh4zEMxJa3GvVJkpI9+KTBRggOwclS87AHQia
AqY+ARjC7qry1eEHReIbTVogfFFd53bjWpfprMY2tRsyV/058RnhkZoaV9aYfFMa
lHu/x9wzNsa+/k0UCiGKo8ocqGa50+2LrxXRnD+I/pKuhf+stxDQV9XH28tsmNOt
Yu7Qtwv9Uyir9fi26eUElvO/fGtDtKEmozh4lkFnUzWHC59qiESB4RP82YYkHRYE
shDhF/EP8rCf2RtrmZAUVRbaFvYZWTpBn/HTbrcjLj/QwK1WYtOUebaIcvqnYqam
bDJTyMlOZyb1g1fAg1GOxyeddOa70nF44ffZT7y1ZwwLOLb3k43i88uRFtw3x6XD
NinFNNt7YfZIJjuPAUsYvAENAdY7ogwrnP+YDouOK7dvQ/Dd/0jyBarGo6blOend
BuKrmoV2d7aVg+fLoze6HUy/qT4TIL6yJcZ+XjJy4WXS+6WfiXqtw3LYhV5nm0pq
ZXWMW4omztzKP8xOf+oVsou9hJ311pLAkH8xBGi8kXVqTdjtbT7anKgo/zY/mvSX
hlrCpfDVPBxcb5gDMN21/5nXqma4TKiFBKiG1CuqSzWWZCRNmMBk0TjOFwOrJRBH
nAVb8NZBUIp4fL/Ih2/lb6AtqzmEIGDR+79XWU4gIcnSXwJqhQJJc5KgufEI8nPx
jkBmojd9pByJa6TItuBDgYE1vGyR7dWUMSvzMyJlv9JxTf4/0yxIaQ38aAV8LMRm
4yry2HIO6eIft9dTPYzvrUpiohQYZCpcSrfucirhaoqB+KmSODYsZoNMA2QbTm1s
BhIjrnanF05JVdzEJWWchdxuYtB3M6+xHVA5cplhe1+c+1mjvyHIic5nFKJVrBiI
/lVQKHLph5Ac+OSQ5nZtz7kPVXnnMEmMMMceo+4yze1acUXcpkW3zRKM+NuCkhe5
DHiy1M0yy3atxDCzpCgD7oJ2nBOikn2B5cwhZsmUx3sLulQnT/f7uVyEH5usxN/b
OBAqr4Dz7OMBDDPkcO/6pKsTCtjMXTLUK3z7voHpuId9ikUnSWyhcCN/1QDWQarR
/M7ol/rqB0MTo8rnbV5T25UY9KiwFJEdFkcHOmgob1g+M5lfDuyeDZ6JfZtxSWLO
25BFPSJgb7/f/jJrMCvPauPrB9FgTCqBxTxC9FjsA5+K9IkgGD41JZQjpWEA6Emg
EDYuu46j81B2oNpQ0cx+lCjv3dSDC6vrHkm47+W5LRUIiFikAQuTURnXfULGPdqP
jPWu1Ece8tJUOJNtzTC3q1vFWsNInac+SNeofjDGOwzV2Sc6mZvyhWXdCPusCDpf
nf57kyp1zL0uvIPHXUnlQGOraSQnBGhFyGmvqg4X6sf/RTzTQWdApis6J8ZwiBLj
0KmsO7tah4D4eLBf3yRoAlGSAV7Ke90xr7bAG8tyhpDnG7cvhC2fEZYuI9wwAZUo
x2wAvCmRtgOT0vxraseoxOg7uQz/4XGXoT0TE3FT3QPKPcjBkfU0SlCy3v0R/gF3
YxQR2Aqv1Q3yCpXK6I9e+DWWIrUit/zkAacoQBUyYL3tDhLFKGJnRLCDfLc99k27
rLWRU0XmItjbod5xdJHY8g/vA59wCGEXZyAzQmFshPTVl0NuUnI69LYa1QTmArFy
6xNc8B5YvfJJgBcgf3FIww0H8HCLfL+UNsTczZxoEsCf5w5js+hUTkOPBKfVa+u8
epPNs10KUZOBYdXTvdw2XgUIqKiaVk7D1sLUbLA7hLoxZhgPpGQxtkOf5eUAgWNI
TZozBiZCreSy0BGFT4mFyYTxFuR6XuBHXAdLUrSNRoRC7Syk9anfSxzXJPHCxWuh
/QUTGmsHV0dBNX5jAOOibUAk2ikqqLbsGOrg9fFlvifOJ/8myN719xBFei32yvr3
A5Pzm9tBPyIayiRE/GNS9n08uuJclBxJNKv3yaHEh6D7MRf+DTHol5odx9zD/Zt3
kkwCzAPJFCWEVkelZnWAo2Jhf1/HWDP6yhU/r+0NxQS5B2gSKjp7wpjhiLOCICMl
XXQ8lCYvPK457bTr3s8Ddgy0hbhWW/ZxibFKyQXIakWKxThK6yK8zCR8Aah/+I6l
mxwZlc00RArixu5u8UHohtPj9cswQh8QlNtoRkyRWdvgN95iGCIJEadWUiotwpuU
QO8cNiRl1xce409IMb7RmIpJ66wZ8X41RP6DRMA0i+gEEigHzWasmy2Zsk3tB6xQ
4fDZm/7gi2J80EzZQNPgpe61k/nKgdfYPH5bmdKEkdDzayvstGQ8jvXF3wLV0EVp
gOasBSYL2gKBgFCntXnUyyA7C1SmGZznQ4pgAkpJT25aoXtty6lpD01r5uxP3eKR
pby2OQGY7+c7LEKo5DBdeoZX9OOY7CBRmpiBxwYxamzWnRwoEKIPSMVPzk4HSt/f
fHrdRYeQkZu2hcb10KD7ge4NpOUUNqmjNqtSGAxnbXY2+2cF4zAdTBjuK0cqpiT8
60iQBM7XWMP/jcfDi3m3O1YqMa83mYYvYzJPD+KWPDeCsrmhyRzEUSYBvZYIUlDq
PBbB1gOrN8ajpSck5a4nCEGpCvmA2oojTgkzmS2YRZyZ2hNQZSrj/QCflUp6PH1W
uFHOmsDQUZjq5u1EPqvuqgcMUTtEwDWwkLzpKct6gW7CzW3ZR8EjfMz2/I4wTZ2A
4rs30nL09wbnPwr8odYSOi16e/EqzJjK5JxgRCAM1xvKvQOyR5F4q2JEzJKtovvT
fSCn0zk+fgt5jQMm0Bb+3sf7ud81PXdblAjTkhrOQPmsKIYStCKnYaw5mgTCYtNt
adny+x7IY0Ws0pLyYIsrVTcCIekWlc9fQQQ6K8rtI/dWe7elagIQIGrHF6pBlcUO
Pv4z2GsBa8sxbg2hXB43WzztJa9iZo/w+RVZfe4cf8eeQBoBtfiehgN6a/lLQNb8
FVggIPs2dvXP8uSVr/dEsPZXMDiBtRQtTGYBL+ifVGX/aBHKJGV9++dVEzsRHXkI
66Y6EuWKcIPDQLIXV28Z1vwUaBAZyaX80XFpHBryQBBA0YP+oAAfDR4M1MSR0PPm
1l28Fihy2VhdBDGjf+vaDG989bwjB0oJLSxqsaR0eKmx5OG+y6SPZZt/p4ViueXl
nTQPoXwV1Oa3KzdnC0IBkYBt3S6gqcbN1AmLTM7nDsvX8fquwNqymYRm9pCpXfX8
Zmu4ZHfBJp2TjNneIU/X/3C3x9GkkhWIqtGoc2fmIKo3ECwrDYDglkqXJCGGMjfI
y0QYNFkq83ftTUAIyHce3kdc6RcRO9eFcuY3fPN5eqr5A0HBFr0L7oHNo6XOXdcr
Q/tw0IeH1IA9bMOXjLrjbRYhioQV/D7WtPKogQ/uN/5BtOQVA3/XV8L30QGdpk01
Ok2jMEDtYWH4QVw+BsWyBvDH4l0EjMV74dw8eVnq6SdPeLMQxSMdMF0K46ZMary3
0ZUHGoCTBulpcWCF7G0/cBdQhYz7eCGWJ6mxi/guYI/890ZOs2YMEoPfer0k+AV/
GaiLvhNGO/mxhzFJOdCllMWt52ITjf7hwIlDjIhXBsZp2s7lz7DLjxFnRXGmrADj
M4YcMzhBM01enZSQKwPqnWPjJLVIwirNeUvMPLWssjUhpv1oRjUZzGWtOOhgOK9s
mMopphfg9tjGndBrjm/yoVw92g5jQ+5JTl05KUTqT57Q/CT8/HvO3P644WOyhJjD
18lZkOLsvqCGzVLL5Vt1p8MPBozpMZNe2IE9CgjW6HVzZX2G19InMLlMtdZXVTZS
o+8lvP0wBAnEZiC0N4/E4jL+Kv5fNewEgMKxrAwzvR/txKwivp3/fknJtAaVdPMu
3zBzzYfO+GfQppI5Z1MAByNT3HH/N9lVbv2R2hKQWeO9j3Wf792/gbmLPT9ufWl3
DFylp0DFbJQ2hHlAZU3+msK4i9+n9z2tx+RTjqciufY2pgzLtK+k2+/cNvenPr8I
n4Jr5r9pdk6zQb2Hnl+EI6wCXTcbjOeQwwxxqVsQh3hVgDm99FmrDO56JCTjzWqn
NVYajMdG9IiJKrIBNJSUX8sdBEj+LE6HFV3q9/3wV4R36byMS9tKxrTH3a6KypbG
VN0i4aN++ft1Q+3DhOxSszBsfSAzlQ81AS9fxSkH1EGhNWkrDd1ZR2kxrVISzT2c
WIwrfpBLZgNrL5GZdk1XDPi/HzjMAdMf1MajvDLYL0dj1OLFHTvk39HqWCHc6fT0
iRi75ZHA5e3+0AJ84b5YkYgaoFZtz8FNN0WYpZGqbH83GNrDvCfeUWhvmuVSI0Bl
pzhHEkXjLuc7xlF0Rltx2A56XMhsJ1Sney1sOxPoEzL93SPMtUBszS3Xua+3HEIi
/bhKMFYKb/3cANlmL81rxv8zRk3Fin4o8YbZkT0tJemy0u/00CTrt5YysG694t5O
Yrw3xBy/7WktbsgA7NR8HTuXp4pf2cN5SrhcpC3+8VJEh4QARycOmpVGR+E07kvH
WE/JzrB8loVQWFhFIJOMHWN+VF7ZSrmNnYJPd/Dy/5/CSeovJtd75gS6dp2kYLoy
3tGhEiOVwQLCROzxCFbdtCGlBb2TlT/e7Ec8tjFtDC1L/1K5DC0TiDR9rOoxLy3f
9pl/JRGzd6pDWgjqsCsiJkW9FrqtuZAwwRO1/9+AieXDuLpH7VMuxLK6bs8/uKx7
j5VJzXxREoAe2FcO1n4TuMcIpoQUuHuhc+tPYTbsIfTmizHBC69QLkIlvMNKeXLM
JhUY8DEyn+RpdlwymGdpf0Ql2EWSIUfsDAd3sG7ZGIU79HAlH/Qw/kiXv8QvexGH
ehL4q/cSON4iadwTgGTHtQ2lWlrWGfgYbcJL8bUpHkZS4dI749y7sKZClXWgLyLC
aavu84v00xdtlSag0zOU5+6CcH/GMPVRVVf7fWRu2yitvoIh/dw6XzowXFZqjanW
SL6Hwx5Y0XA9luAqDvNOXpPsR4lEn48AEU2Lzd3B4/YmkQqWaETzt2fKpzAXZdqD
ZeNPUfxbdN9owqi80SXrcq2L9nFTWgmlnCvdeXIWr+qJ17Pi4X7Wzj0TrmHKc4/0
JXfQEapCN49XDUYbR0XusiAgFT53qidrPB4ZIaXij7+nKWcxLI9o8sjSGFab4OJ/
4WhLsOUKoEXvppKSM/WudewcECdtpNlk8FGcnRD2/KrOXv2dWcr1qG9+KtB0BcaT
n+iEWb7tGOcFwkhTtrETl4N8Z7uK2NPYFnuOKShSFr0eIfxQkE40zpfjUTl6XtX5
VZWhfMVEL+G0Ja9oYB6R16rc2FGGO4NFZNkEaBS+1YNjxf8+O+3HYgjRBYLVd0zU
k1pjzRELbyeSZeiQyzAyaftUOokDNDrba5nktt+CAdO8RTVR2lCxkH3bEMOykFMn
DO7aJHv4k+jJH/MRi/e4cqi6LY8wrCH2DJ4GpimrwYx2O7X6L2u2h+SB/8QJIuxb
plczKhIYn7YEATam3gsekUbszevUy1o4z+2/z0LVR0ygkm/ft8D8B6dZBQIKuxVJ
OT80hPCZHbyuG6AuquykekKDIC3xIFzDAA5Wc/7ifLi8vkwluJ/jrC/NzMiG3AcM
EaNG/osW7fCXw3kFw9s6MgR+l1skDbFJBiTWTmoWIbWh/1s8iQeRoRlnyPcXjVss
1VeB7hIaQB/vY9JIZDDPyw+R6LUzKSdyGnTzaGkWXdt6JK+gfvKOyIv4NexacS/t
jMmvRUBFbasvx21LFWGpww2nTYHKjJo/VMQjm5dFvQ/bgWEK4+T3iU9IP08HxIIA
MAES4i6DIsLsC+tCWnO3UYE3SDKqsLpgLD6ISJmqZcxOUay3bKy8wsYtoBHsyjG/
qN33y/fl25UR5C5BWKeLVZWo4LOcNP5uHkyg3cxSW5QVvcyLCORZs/GO9pYwRxTd
c3VOHQQzLQc/bE+8reg7E7H1GmsaGV/sGbAdWr0mZ58djIIije7QboDRJs8bKnrP
euarCJ91k4xNI7e5AxIFhVv6A6WIAnQd+cQE9agaO/N4yB928asPQqO0GPPxbmIY
3smeMwvQzCeSr5bXg/T0wI/GbEU++h2XG9PPVPO6/ZMQlDS3kKyyqIWNbOgk4yOT
GbI6EUlT3vcmEK9UnHxH4cJyfjWRYlXVg9QvnUSSMXNaC9auCZIjesM7TCgTIw0w
bDabbrzc0j+yjwNUDpuGSFKXzK0kyG3rvIHGiQQWid1VUmWnmFNBGB8YZwZBFFFE
3t+7pdguhREEsBrjQxrd/5je5YxuD7DxHEd/VkhZhKHwQl4r8+veklEXDr54Xhsz
myBzaEMXAt6mgeb+8VwrzixHSYxql6q3ODmLIk5zOfd4h8SH0PSHCg926MNJ1jJ4
AXaucD4J3RxxJvDAg4afaRRVjPtGlNRNf3y5OvMOUxRDlsrAwngst49guzVm8qfq
a4FndD8jiobkzpwp1xORbuQGt1XOZyutlD4Eym0x+fd46blTw9HUSH9XwiyAsUZU
1X7LUDouW4gtkIS7sE1+NIcMM86o2hj9DCumWschplBzn1/yuOZ+JX2SUi881DEK
7mVlFHNJayfgSc4driTn7aefreDdtzKZtftyiad+RPM5oPIPn7piQkZbKaIviP1g
ikY9pFOWZ1LKcxZ6YT1ZOvZVpYm6a0PXgaO1NxOvmuwqnf2tGIUN5HmVyob7mbsw
8v5WkOV4RonwLwuTI++ceEOgsXk5jMQXCb6FZYYVdVQs6btGgwvcr2Vi8bru7sMV
V4GP+jz3VHLMHwb588jpf20nGgUjQpWM8CU6IWrJJPsFdJvsjX71w5UYeXVP2KYV
ASC0ULoq2lhvHJaCMdsrM9DvJ7ihkVtOmiIn0psJ8J68eAuMpZQdidKJW//eY6tg
SCq7G5N6dvWIGv50iNLVKa7XmNAyFZ811wKWW+HXuIbDgDJFk+m77j+6yeejwqAK
j82R2E63hgeyeNtwBLq1EPTEwXmsrq4vciFucE5Nsng3VPVinmY6NWGWs44r1AQw
DSfMTEU5krkgrMKKnT8t/FX66hAA2RRFZ+tJwszph4Ubbz2z8KR2FmjPycZT1MFZ
GPtHUUNVQd2HSR2UnyubXFxsf+92pxi8HgK2VUJ/FTXG5KC9lFRlKbbE2b1Ebttf
c/et9HohFUO6qk02iN1+f/Lc98koADg9X8p3jgKGSI9UnPVvXils8llPLepEaYDP
2YdvX3eO2TuOpTrvlr0+B+eEu5lId7L9fpEaGe5qcKkqcX/S22xZpZJtaEEK6OqZ
ICem3H4nd57TpqbpCwtsSOEXtJEpDrYEuIAGAdnlEzp3A8lzbj9hTfLxMcPWuGyt
uiJR1gJlxnihhbQC9i5yUHcghp0Q7keLgBYkaaW60i75Zyc6STq3ELURJX2Puy+v
wL1JjVzh3DrvKv98C+mi24KoeEZ8LGQJ/Vmu0tOlXsPF0hgxn/a1ygmPMe4KtNnW
DDa5C/1GBv7hABWIRUYDiWlb7JqSj4ShrMgl42NfkW21X/pLYIX0tx+SSpt+msGa
dOtGOvdVoHpO5P2vny3zt0AR/+Cbgr817NG/R99Ed+47GWM+Si7pdSQ/jTj5Uq3u
/nd7UR5uAeePKYisZzA15PRQ42DkHZ1LBkErC1JWeVtIJNqkrcRb97W5qr2+0zf9
epge976u2TCXauEIfBhcedk+Qb1xTlZ6dG7FBJS4ogkUkZ6R/i0u43gm+J1zD5kE
ZB0Lv0QI9T+7RHkjkZJeJEwh6e6A+y9x6fErUlMNW2RiKs8QQVblDfCwDM0MpOQC
lJ85E2ZuHgtv6MUzX+9qmFdwREC5JBn43TWT3GEs3cRZJn1YnmlRLY7r3BMO/sPO
T0zxUEttxg8gJtI//nPC6OoNR4+YBNEY/Kv4LHucuYwk40cxVIu8shlVBuUz6ufj
OA1FLwz5AGq2/zUhKD649b0+tlTlFqu8iV/Y++jWtZIuESK10IVkx3g1cvw2X+1/
TJ3Nnk2ffElsGtLfMSQI5xVXvC3B5KdqcpGJCyabGwAR7Iv4SmBxjhWml+sgJZRx
TWUX+tTsw5WxvEueK1MIwUYlaaODicD9pXp+bMNa8K4vCGSbUVo24U3xHeXnCxSt
390vq33xySWPxDIBYCH5xrBLJ4BGhrkAjjJyu/UqMRunUFay8jYHF5v3sGsJAGGv
t1jiCoG6t4kx9+YhkSAnqFQWpwrDO7wqXEjcKocB9vj0Pono3FSuN3qAQGRJFGAQ
zpstACx12AAmSDazhB7fbnK4J5U1kZwRbcKIOi8/TmJFfmzMbm8Uq7/43/WBvfzN
MzGv/HLPLv6vKLdmsA17wH0SHa1VtIjB2qe3LF84mAmR3sl/+v3bTurNJB54S6NT
zzVGsFey+f3BUAT2RV11kVbRRYey/hATRgnxOF6kAT31fF8Q5Dt8d1HsEAHJzGBd
d+TgPOoie0gHY20oIKq52ID/RaF+tx9zqzMRtWElw5Hf6tipfUAGRnJkyIy9xvpO
IslDoWhhEKC8eF249jdK2N7J0kntUveUxD36xHPceROWNp+ngCj1r/H6BL0LyC+q
HL2Jl7lmY3t9NY7AuILAHCJvP6VsR1vtKndg325Ucgb3vG9eeK2QqSEiATghO9aj
wJ9cEFNzBQSju8+vPIozPxQhTZuTLs+Y7463LYdOvj+4nh0avlI4FtvvFypE/gWc
o6bKvpVm72olRbw+v74Me2Rr2UdP/1eAXcLNrYf4edciddc5u9AokxkET/wUL50e
9EaUGIugNYg/YHWV9ojEg8z50ENX7n4/MH8DwanDlFI3jkrwSpACccIgcvSOq0XD
/xexthvihxEd4JFzTfKfkL4wt6ovp2KKHTkb9pG0o3lTrhSDzQf6viFSUxZgibxk
GEMAtEJAGmeJQDzY11wUW7Obu7fAQXgSI97l/sY5LtjVkyXHB9+yX/cPOiRglO/g
8xUPFzgYZbD253RPqkOBzX9v8kRtftsaA5KNxOirMK4m2ftfwNqi9Ct258USFcsH
+1x6ncYMYckzj636NXKyZYlQdF4NWxfyUnGpQrpeF6+A6EE6YMaCPvBxv/hMLO5B
Z1ujlAouXgoev+KtT6rwHQRwl7hE4RNWmrAAgb2c1gUashXn5hgqeYrzY2KwDJjO
i1Ie6yMcPykbwzMcCkCJNm8/+Hr/DVFZjV+gTaW2W3mbPvfNpRGjxoTX0UDpLthA
Aj4vGdgC6JydeiSJp+r5Rcz9gSMBFMw7f5dk/ZrNQqM9OGfW+ZGgOhlAlJVBzSHp
Fa6wgPMHUj3inUKTItSl0aBqn3vxhx9ozft/qGNDw+9k8shY9iBUbshBP9SE/L1P
FZeQMC/TStwsZKV8zUoS6nsZE7yU+hTAz5oF4Jh2Wl0LnA5ntlAI2SM745tTVQci
4qfy6Nze85i5oDjgimu+j4ELUuDdfE1gZeGvCsBAo3nAo8Kll0N1jBrg3ic5VgVO
4BSvT1Gs2qW0I4aN65RDq3EOTnfPsbUtMYQx3YwUaAMg3Zb65RvjF7kM4BTAxSWh
svD5X41ZZtyd392FkCTR3BZ9cVIMOnK1RRJQ+1C8N5dSAkGQK3sC2l9xm9nhki7H
vUuOGeRgkyvRjP3JjA6cReMBN4+GQnoNisno08cYyHIar6Gp4pk+6M87OotoTIBJ
GQstira07x7NA0C2OFsJ/pp8lF40oKsmv+Mx0Ta4IlP0S+PHJ96qQP7Gj+6hPBOh
D19LPV3RpImKcUKWOwMlbt40TUO6pV7YcN3ft8e0t1eQRNFg7I9HP+sku1GehRII
YLyi4RKG9BVyboxZ0bsNwXYDfYAq+v4OKDsZGm+9d712LUKpBskqJyeYFO0clUUh
9JheD8vZrh8tgHi1r5NC0Gtn6lvsMMzlg2HfZ3HfRhhYgti4hIE65UJSyh1z3DAV
rJYKZqdDsdbFsZ7CgwuvyEO/uRh3I6/ZuzwVN1zYiCTNe5P/qSLM6RTI50/brgiS
L9J61hRfQ+jcTvdxezJGCkSAjjs2E40Fkdt3vl7qXPLJrBx73rFy7+4UVTd1Z/q8
b2hQGZBm1xYsvvR3nkEtBDbTarOKy8eSz2XLvJuoqHQxId2obtSbyCJ8wiwwCujb
fDoI8BJiWj5DEsHxU3Q34QU28ZlWuSWx5O8sWLFbCn2fmYLDxyrmN99GpIFem3Ww
fRBSW4EELJJB7kb9XzEmE5sRcGkf5qDFR4GgpfuOzwLZ17T/tPpQExzdjAtTKkTJ
kQF+v8zH9+xFNu2vlZvmV3E1os8evEzxd01XCWM6/UIWBjeNqmPi8MirrfWUjmcU
B3Ew7QzsVr8YuWjyeCXyHPRCJjCWTOneJCfqijBk2Z+9HP0LPQLx6j4wRq8qxfcW
qd2SVkdY09fokcWV8fZcSVrd0sfSK709b1q56CoorP329KQc4y4zYb6TY9oqFV74
xNHLwFqFwGcm5q4ag8KeMFva08KMmSJQh3xmES54PjIFSSUli8ousM4H3RpBFFTW
G4XUBJ2HowSlg/XjH4g1Ogph1MsmKjohUEFsQarov8q1CcNsYehdrdO60QdqeRaO
YDH8givfdZEb+PVbYZJ5zzCPblrzSMN7LmBDEeofwPUfQKhFwpeIsu7FtzsHeouR
4cuF3RACSgjZjhF0RHpULxgbiLi12CSxz9dhZ4f1OqIosbYPegJFnWG/koUJ87qO
x3PvCrHymzSLIBBT2T+ysTa9cU+PCRLOPJ/WJkGjQJxYGiTlDksp9kEgbjztLTRJ
RRlgxFagl+Siajf4bOL50ccV0X/P71sy+NGE/BWBtCbSp2MaSgXhna0aOmS03SVU
+J9616soly+N63Ks70yNPlk7sDFzKb4GHU03w8VcPtynQAxpX+QRpj/JBopbyrvE
Y5oUwF6hHXRy4e7zoxUkHpZdWLa+6n+NmDUPCIsk27Iv+xe0iPrjrsf4pgX9kcJO
34mnT1pA79+BgqfCiF/O6KO+yXX5f7J94wXb8LfPSTkYsqU4ObeKFiASGrb2939B
OlB/FE0SVeqEjF2TAk3er5dEYMCmuBjuqDbDqbXauooISmLY1ZVXJZsBzRsrGams
k1yBtyt9vLVf2/1I+bgtoHqxo3dITdKcFlLZEG2ITvPC8MnTi2NcX+aHzWjE2/15
c6iiKpVTIqYiiE/QSI0+V8rFKghLoH77GPqwiwFTPk+cwAp4htTnKbUXpZcPhhpa
wYnDypqqWCP0erZOVTvpchf3lM/3qq5QPMgFpyV3gBM4pKQLp7AfPAQtLRRCFd5r
00JfbGjfSwh7Yg8JUPjYOGt6UezC5RoNLAHYP0tQbH0cSCLhBsXXyr/vpKMYEd0C
q5cjSFNoEObDQUDcHNi67/DRjWOSHXQb2I+Tj/1l7+c85hvrD19ifIeq0dfDnlq2
7qN2JuaouIRWrLJMSVfNyJVutTbL1y+OTnZLQjlUF5pdhuZtY0UY/2yeSYZoraxJ
o03ldls2u64qqvPrmhFLtmRBjTRuyAKVG4Wx4S7tqWes1Oes0zQNKvSbbGqIa+Cc
ZbCCUTjjvt1WwnkjO4G9LYyfuNYn2ixKuptG6mNiyVnQtWYYCbbmO6R6dFJnzM8I
LV9HMiaxQOrwJlc2q+qa114pEPGyHS5dDk7APLKmUCDAtKMQdN7soWSmxdAyuBbo
l3EOSUGMqOKhasnkjIH8reuwTT9TfE5PqM4xvgso58KvQEkaHhkChYR4CiYBYHXT
s1UyqMVibrvUE+B+o5AjwzNX0x2jQaSjIyui2T3ZEHQR9/QVVlVrVMRx5bEtijk2
1WoNyiXBYmRJj8WQA5lUvGtGy6RIxfO9HBMEbKTJAioWFHj+DyrVLnjYtEdXbMaZ
4v4vrWaQM/+jN9XKh5GopGqxHDdwbl8rv+JqVqihVZ5CZURnSHuJ8a2yrBu1Ga5E
LgzhJH1A6gEBCHazcBYuBonnYZqNWYfU4p+H7ul8hXDAQzJFqO1cqSZ8m6BAw638
kEDEuxq+VvtniSMwCLJPZ7qwDYwiTFLj+dJTzvUWji78W4FAhDi9qBt0RPDz58fU
IXdNLgs/C3LnjpUNYtwR46UEfSGvlvC0UhijOTW8hvL4E+YRgFHVe2KcymwyQQuu
F1GGmLViqkzHtGJqdxybjqvcByQaR2uYtd0c2CXyxrI1ZoMWqDzsC3L1aWndu7tW
xS86IKHsXnDfBEUPxb4ubmCVDM4xwFru+j/4bWsl/YdAAtjVxuge5ByZLflpIj9X
1q275Nem+h75r0SmOc+Nw5/2FxxUKM9tHNOPZXwotKtPUSi4IVLBUm+W3dvVtKG+
ERYRfUbQv+078Nfv6fo5m5oZ2PfDzjyy2y0+eyWkcWz0/AEV2w3OPW1JKg1rPWvO
zzrUeqhZnEcH46Q6ghP+vX3eErYsx05PT9YlO+qyjlmWIMH4dAahMeIsI1+pHT5h
2Yp+Is0nlaI13r+V1Za/UceDYCLSlTj6eUhv68eDC3yF3pJemPDL5DZaJzFISh9N
01dWzlB26nkmf31BM2QSpKqCgPw5uq8RFOZ7mnsyuVzsvIWKPIKPKfmxYKjyPUT0
qWJHJwQZxuTgmld9BW76c78+0PScnJ9cp1WasR5Me1M0nqF/pAxC9wGG5aHM4dSI
Bkxidgt2DsP+ixv/2+9KZp3/P5GVaBfZSCyf088j0ONqJD6boV67avM5Mw71ih1E
E8j1XO8u1eHnh1HTRh7sgEptm5Ks9l5CfpWDVsJVTrPBPkCP3AIDkxWewhCl5L6b
tkzsNslE2KD7WAf+Fah7B0SM+srrP/0AeGy0CbLGkhEdCaz8IFwcTxJ4QWJEvBFi
AyTn0RwxtQRso4H1CoRzB3/CrKrqINyVruL2s8FUqs9GZzGmppFvts3XFiRlRGg7
7NtGrZEtnVqov7bmWKsy+Ts9R3Ct+n8cbXNXxZKtyxaFKaTAmMZ8mre6hsMN1B2n
ntmk7fRK2A/DloggSCeTzX/LeSJJlaufJrdpuJ1z3x6SddsCghJPchii8EqCHRB3
RhXJw7w/w0orwiHjRD4h9xqnTut0NSwpGdsClPKtyml+qy4CwB84knpmInaM36ts
lQhqd+vL5delDu7LfwCtjrOb6quLxuD1a6/1v0I/HuS5sfOu55hkaum/CstF17jU
3PrTkbSa7qZp1M9jYxrBhHXKdtnprxgc8N9BgjgUs3rhQZtxSg7B1wUtMXpVptk9
hsHXuM1XguovOSqy2bS5VLhR6odVsnA7sb9hs1Qj2g0f1jGNXJtbJl3yjqWWZXUo
KdFSamHkTXibcWwJWchyMflg64tXOMnjKUgZhrDL4lz4V5pT12ujiKAFHWZLhzN8
wvD3cr+2BfPAIfZ3XxhkFkDQgEfXyYTRc+So+RCn1fcXEIJS8jkY4kVP8QazT5ep
/BTDrieifRhcvgg4TeGCt5ef2MaL0eWyVazJo/MOFHsrcCcZd8muyOSniF7aIhIs
nBsaZw5+FFXIfk7QwFL6VMRgf/FZxKZmeStxnmtyIy0jYzgJYV3ElQhcGevRMKIC
9QXmdBX7+93i6I0t9wN+UAviliqD3+Cj799x8H8DHKkhER1iyVNyJV2ZbFLOf6cC
4FG9c4yhjnYlGpii5u2jpIaszxP7z8wYuUr1choLj2v9J+ga8dIKh/xZrEN7tC/O
rzGE3iewoiMxb6z7vD5fZraO6tXYVpueFg5/t663uoS/jbjq1qpciNQCkiNMtU3n
9PBZ1QwIFrRe0wHfKutRZ4sziRTIw6OEK0l9VbRl+G6ffpWoRrygrzEUM7X5ipuT
zMokEsOWBQF6OFaEDcvZoKzAaUEbXB9AYjc51Ra57X7oD4QyhGwj+yKwTwS2Npkf
LjmjmFtwFvXKukMpztpOfZiEC6aDvvlB4PHMq7RUv+wNGcsouce5IroLuvU9CiZ6
iqbynAMujJoUTnISRMTSsBXl0jnA2ras1D0tuFnkkg3EX5EYz6vkeC+I0By5lLlx
PX6+BLruckFuaZRFK1IYUapxXpuD/CoK37qb8A63A+6j4Ah6fM5BHM1nCGOU/U0+
oNh85glMMNvr3eabJO+TeTR1lpQyzhHyxybUl1kq56DaIlaWMD4+dyfdOfyaRI3B
Dk3QyUeOHFAnptSL8w5WcvVjxpwOzlftkVOg0cjfLavToVXOAlnx9tQh/6i8XjfG
goEq7O7dsuawNMtzr8m+2kocd3SIqdmF55PqVLe821VtGr4Ed0jHoB+pFNi+LbPO
Fhh7oIKwJFPPXNAl4Y3d6wqHbiX5EtQtm6SCq+Fht1X78Ad9H2z1jKPKVpuL1Pmp
UApCBPOVXZ/XaUpqs+/HVL+i+XFnHA0bokiUKodJCZpG2QZ91iHal5bI6NAwaEwR
xA1TgulGnvUnC42oau+w+iUS1NXpOjpalkPCwkB6XPg4NaVe5Z/9BoNEUKNzxXvk
mpFlTmodCflffPJ5895+5L7naJj+/0C2QElVe7WMgQtLtlX1eBXTF5EB9nUKKmPd
KGSTS7pG9RfVGPPD2pdgsroVIHZMwgkPq+kO7mbZJxE9rRBhknYl882LvvAWY8tF
VNa+sw3furlrpt6WuQfgWQFqyU/jTXxB56U6sP4oAzmf8xh7hj39LtVOL6Gfd9Fr
WWLu9HssQoJXSBUXXweyocVBHDD0zbmMngWVBaieHNHf5BDxGYmsnnlAQm//GWGe
DOGEduuERZn63Jut6LOiXsVd90g1HhcyQZ0WI3tM69Bt86U/hUrGXwvcEaIKY3Dd
EzGfkskbkJY5dPNtQvJ3rfcf794dShE+6tmBqBaWNck/KsDN549Wzp29N/7CmRH9
WBymKm1+wra4eb6KRPWkCoSaVyJMPyCRznIKqvW/C5YckRYRluU46DYatlU7LoIo
mdKl666nVyyHRikke2KNfEYwHw/AYWn5NSc5Iokw/OqG0R0rqTQvP6kT4tyGrd2o
balFU2qXI6lWt2BlbSwVtF+CMCnC77xt49rU2KzE4wccUaf5uSaiYZ8EdFVoAw5R
4HDt+j66XpsSlz3S2Mg/Sj+EemGqNPYjuImvP7IWsbaJXv1A5tyLsTQlkaD81og4
8EsFBvYRy99O4N66WT/R7rr2FRDeyc8aRst9hBPUxPNXT2ZgMgBfvAXVi3QRiSKJ
wgqivLjdycEQUyIRurU4g1x+8agdj5AoW55Vs+PdXK7llI5jIX6MMjXhbvIIGGVL
q9t5/IUA0N5Lq0P0uJH5+t6HfVrmZnpNmWRIIzuJDmWPqFlBY0AXcSLwdSXh44xU
bRL3I07btfkwnYJ2rHGlkqSTud3USc+qFCPJ06IMhYw6DjWT5qIszPbovDHd8W57
uPlvq+3+C1llEexJCDRDqaJXmDhSBmzBtyVdicv8d8pF9Ke2tXisD9fzcd0rpNRg
GNMNudKh6NMNN310h6GY9r+m40eY6pcAuWPq+tRrPZsCaEDG65hw28LW9w4nhqoD
3x9A3b2vBx9eayFBcU5J+Rms6vAlxxpeJw74UVf/STUUAalcSJZDixLo8rrGVfdu
MtYGYHJDOOOcytIAzhtmqFph8kYAbQAoLsw7CHkoqCsUhQvADHTJ8G8oGOqVDuZk
wb4iEa7v5WXPrARdRCcPJcgzfmZY/w9x4Uiv1rNHlHV3O/mkgNm6sXEHoGeoDN61
Kvz2D+1jiVtvKpDkADp+MrzYh/MNfero0ImlWqTjNSxr4awXPD6RfMPms4wnkcaq
0pvJ0wsz4XtriWb/T4B0I1mIGOexuHqC19F9/ddqYIU82dT9j1bis2HNODlryZs9
B+OShLzf5dBIwDjZWKbNbVeP0ds9fkBh4MaqqsM9NvC89inRITCrJQi0s4bdDfsp
yRmC3KpvTPi+2/KMmGie96m/Z9XM6wOTbmdgUEGOPxGzcojlH7w/g+70MLPIG+2o
RC9Kk6QPoTftO+1T6uw9mN/T4Mplba1fhqGgbb2rH0TxImjVXP+yNGXQIpPx2xgw
wd/mhlhCF349c5fJ5DMhZBoDM+x/d2tlArMpuJzhe6YyjF/fbDhr+qU1cN6yzd9T
cTXu7gVW85dmUw4WNCaSeXOkhHe84P5eWjAU4RQSfZpqA7p/ttFUka+U5p/BvDfX
JQ7otxSvwmJo/VZNgQ7eOZ47mASa3xt/iCVgyth1hnopQEJjKD9+1rMyr2dGbLOd
jOUP7Ae2u4LRq9shx6DglHIN0gZpfEQBu2NdH3Rt24L5NFk74hKTFStjqPqM8f/C
ZLSrZdzEsK8cSnlvdH3RGVCqUMITPtuXsx6UjC7BimCU8yq84mTenUPcNudlbccl
hJdtskbTKPxTti2OA8Cif9+y155eLF5h669uxCGRjcrJ3iwRYJNdfZiviOef5uvX
tDPpqPJi8WRD+0GtWU5lyIJXf9dBTNKlZS8fdrUCRuwqVZr77u9P7OO7zV3Os/ch
+RH3HmIWPuAjwowgqEe0EoEYJFARPo/BVUvgzfuyZlow8obu/TaFlRfhGCRVnVZe
kj+CNPeFlLfKlU9NDaU6FW2W1W7JapTlN4FlC4CmNxJqnzWMe5CYzuczVN9hFW9g
1Xz5/O4nGi4J4ZNu3ssI5ak+ECEhxipZe/+1vf4CNrT1f99Gff2baxrH0BOl6tnH
EkA8QdxcX+clIBlm+yMETawoTSRD+GcyTyTw1OdBv0g855vPRXTE1Jt/5OH/nhvZ
Y4Oe3GEIRpXOhVtaDMZMWqwwl9gFIcwUYp15fd9WaN+BiL2wMbKH3jOTn/iwtbLH
Uh6zgtL5q3+tdQBSgS57BtAMDqHyJ1fSDbLxVb5+e5K+s7YwkJHL5fRLaZSYlzVr
YZq3Tmo3hMMOdaaxIjHaEdokRew6+hoBQqmce4SUKKeJJfH4/sCIJ+BPmzxnbaYM
L2xXmt9LJw11j29Qww9nM7hKJVgCJnEbE62uxL79M2/gsr5oDXRYbak9MJ3WDzP+
/P209/a9npBB1cWjbpOZ5Z+oBBcQ2qJyL/4VUWAjNs35Hz3u2xZkOo6uhUXaNiim
5FwbYtvByGenJqBl5ixzssL0VjgM4NV2t1m3AqwBZvxTsXBCUjwAPy/eSItBf1jJ
BZo0AS6GtWl7POBtdkXnXzN0hyBiVxcJCfSCbGXlk2w+5LS9mLljLHUbEeJ4Bx/X
Nddpd4qMltyCz1bIfAZvHbA7Raj+4yG24SIuTkGsAyWP3W6XvGzSTYJw7Pp720qO
z/8Oy45ATA1SYZ5AYiZr2EgaK0I7lyO89rrvO5ZslYGMzwFojKY3Wr93y1K7MY+q
DVmIY+Q1/lT4Qt1/4tFYT2bC3tHOEGPq8RRjG3vLK9McwF+hR7zjmrOzOU95oB2j
CCIQT3v1uIxbbGyqYqvNIifP13QlYP+2wNQ2x4lzWJC5qwHCAVyol6hxWKwmu4ix
mRq2k7qzOnmSuUhK+YBc4J+GaAuI/XomDYF51ZzdcY+Bid4FEo2FftOVaoV2wGls
whhXza6m+FRMuT5J40sNq5BhDJ8xYGULtE/r1L6MWra/1VFC6eC/kXCNbggIHeRI
4PEWOMVcn7b7TBMAba+8D5hbPK6wNAVABDL5gDFoKNyBGL6Wjdv6874aYNjrWqnI
ya9wjSflVhPu7gK8dj7j6hZkHmYcVO9tOr3GrSR8Hv6U0KKcKCubhpT80VXwn1v5
8S0h+jZLcz3RwFyz9lGdeLyWrWo6yJyuaByyAZXL2nTGwN/zOp0AZ1MpuZ1iAj/D
Tpf1xRiz0VHVTBSmmsaRF1OO3KqRO4uRri6tSfYsQPahQwizsbB5/DG0X0tTyk8l
r4YO16dOnzoJVsWTdP0d5VXgKoQGEUk+Od5rY0hznubkKvUGcnPoIlMAl38NAcrT
mv7OT2T3dIMrxpFQwzlHbt/9I/xKX/yVI3QHmWXCSYcyMj7YFrtx1xfn/r4+/0gk
kl+9GuJlBr1YLi0xOuj/je8suOIpoxvhgMta4+yv3iMboJ9FlxQ05Ur+/bc9fLcS
2o1Ig0MHm0F2LBgpB7TxdrWp1rsbtprb1qdyn3Lk1v0ExnpOPEtif0C+nLphSb+m
zo8bAWvdaMkSLwR/xqshqpSb8UYI0fFYWih9LACy+02Sbd0ZFBW/I2m34vIbpgon
WDmo2Xljl80nfNbv+fLgG1VPWWFP/ScXwZV+sDTFchMCHkU8rBX1n9yIghQYqJme
10XXUisSnF0nzlHoYvkGUW5YNrTET7349mG10hs68bSEP6qrfmRY/dps7/Nmh8z/
CBpgbB7smq7bIl5QKR83pu3hHMfVauGdSpJhWrkSMVNHDQDy5wCObWve0ZrASfTk
Dh9cTogPZaUbzKTvmv2q4XqOqbs4k2IjkQDR37rLyVszRrt6+F2vH+ODUFZiGH73
9GFU6nj7JURZCFssspXgT88tlFM4TdAtsW0c0mY9g4xIrR0Y4NuZ7BzQFNavwEi+
A1sYHuN6FTGBf2zOjP2NUX3Rem0iO1IuZbqF8c+GsHAjysTrUDPUCiNQjdUpuc3V
axVwP64MqK2ufZH+sLgRmxQaTgTXHeh03bMitYofRHmeFW5gvl2bakERteO4MIPh
I9njk4kTc2rXF4kh6+Wyyb+R8wG+bMKy2iOuhiT3LuysVl0xkjcuqy8wZGb2163g
PaSpa0/V2DUoq28gzqdStvQ5M6w1WQIyT/TqoGiB7hgCW72vVoiDK8h0Eutl//DT
I87YjNGUtKtOercdiZJzC4xCQ/aZPqJADims5FvAkRIXBupVlacZDcgHbU2V0Cn1
NzWNbOBTtFrODSpILBoLr8oy8Wh0laGvqq/JrMC/CQ7O6G+p3bCYmbFtbQboVPaR
1VIL8UFUhjiECFvfsJVcOfldGvVfT1Zp8TaVt5cimPfs0t5C4aJKLLMhzTBtKcfN
TWxkdFAo6XDQjaOeE66ipmYwLXaaaZn2dwcEGPOYh/2On30dN27mEayRFepDXiYt
QmEV3UptSOqHYELOqVjei/zkd/tYH3DwoASpFuQSxqR7uJ+EUveyj+CBVZLbXjJL
9NETLn8RaEmGAEXt0NG8+IQGG9xDb9kSOPNanGwhYwO31Wc4i6/FWwQQ2Sov/buk
U0XhJLA15JIdbPx76yYxpyduW8DErF1Hsmc2g4YexA+jKf2YPMyJMMLV4d2cwZ6k
VOmw3z8/ZXLPs8ZtFIYh2NK/UdrWMsKXwAnsN1EyXSS42VGfBmDMevK/aIQLI2vq
pZ0XjjrvWpvMKZ+xr1Lqmb0RjWIzqMQ2edK50VSAtZo8zDa9P/5AibcenXT68sBe
PHxNKn5SUEBCmnVZzLWma46ANe1KwZW8stnRWmMzJ7AByM+w+7FHtgvblw0fVBsj
IzADzRZRw7TJ8dhpchHfLRRTJSNaO0Ut+pKHFdEXmMjQXO60zHYnxHCMckRRZYKX
W+wHQUl0HPlro6zEjVwEdPVOmZdH8h00zh8QL2WjzLFFzZ3LVktGpB5njS++Y/ZR
tTT8K27CZBNMEiwTGaujCmCOvVp+RKrKRPLueLi5Rw/DWq2h1k9yAQkpCPg7AHhq
8Y/UcPorc1Xei/NQnMj3TAtHfzMJrHtunEh5jMlguoczx4I2g9KhUYI+vNPNJoEP
TsjPeAjm6yh4DBEG7jPYsO3Y6b7NphNV26kURveCUHNOUo2GvKNWMqkHeBpu3C3J
m21KPiupXKWr1JytCHtdqqbL8iwLfW7ZitytkG+bRHqp+rYAhWPVjVl/uOGOLxWa
7tbx6sjd8uHjxbyU5vihkfzA+AvPGbMbL3w5FjjArtUEksZ/2Qw+ORwzdlp8IhYX
/l+2BS74bVLIvL7Nu0Cgxv1NeFAfbhxDY9l1UP5t6UUELtxr8+IyHDy2Gczy/7CK
4wXEYeXnuVCfTla0CVavJIDUG8Osbc9hbnL3qhc3PxbUQ21oOnX23CU1OLPX67xk
yHCoA2FI3pknumyoC4H+d1570RdQyanQ9mRFZkPs2rWPAsWBu+iC5CH/gx1gs6iz
9uxy0nU9ysO1U+cDE+kG7/NbHDa+DY8VP7DUAhjXCb7XdHpJOZ5TcgGJ9sQD1Jli
Y9hRF+XEH5eMz0BerXwujXkoeAPVZO1miYjdvne2PFYzWfGwnudkyfskpJABqMgF
uZr8XUxbvp/l07Oryll1QBMeCgK5JV8B7Hw7tGxjKkseW0cvdhetmllGmVm7sJK7
ApgNscIUl1teTYQwM7lWhUB+puHj+DXPWeJncgRNs8aSpDu5Qa0AnmYR7nPI3FMW
k5zjFVvJWzm66k1Byk7gmgRk53GuzmWkITr2J3WwrFQrV+qy4Wk9I2E9CCfUE1by
7Qyw4JKFa7Fpt28Sg+92g7StJCtLs/+8FfYh0RFna5POB9nhvu/q6yY9eLESc5VR
hCLvZkFfsYqddVUtnxUKYc7jX3lWlTxEtqSCXGA+NkYx77jdA+FI4NbEC6uJDdUP
rb0yT9zHWRbBjzeVA8mV4RKeTnAJaUrGRVH20F1Jq2kM1izG9rx4MnRksRlItUZA
1CilxgaL02T5ewtSQvz69s6Rt5PSyfIz6jXoxz9F+gqSpw3qDOPKyCYJ1iLv1qmw
f+sVIYfdHJxOtKk3Eq0LMgZS/eCdqDiDqYTq5toVE9dPyn4QoOgEXllKUd3YW0e/
0GRw4DjCced6krKdTL87+2n7/OlFRZ1xhCJdj1m2VVQv44TNlJZ35yTfZJSmJsjX
ismRl3C55WtSw8dxrokf91j1gkVABYh59h7hrU8SAs2V2/3S+ggnNzbDDJQIR1d1
VBnVmkGKZuJAD++vzN03pUYqRXGxlmbaVJOglnGNcdjOILpDU+RoIZW4T56/xJLv
tUj1Qqv0Fml9u+qP+KIdYQrafmMr10I4aE3Ga6DErC6yZsKLw5lex+bwfw9x+RH3
R7js1+5NiYBQtSNQ6wkPKfFs3QFgR9coS3gk0yUc46cqUs1C8c7tAu85LJfZVN7E
NisVDmmxPDw3DZYL7oNokEsG7YyVlPJHe9h5gT4YGBb6QbCDTU4jDVOZYb6oEjGA
z4E6pbUNK8HzgkFHC2jD8R50epbpnHcTsxYgSbSiiOb0G4BjQZz4rio6IAGBjcrS
k33hMEfxepFeaxBm5m3qpZlMyhgWjKRuvDM3Tn9WSD/zSwejD3j2cQwu6OlfvXBT
b2uj7wfTCbWigTzhNfrPb5lWqvtLaNA2TC6U1TQ1y+RRcmY0vRVg97vzYWzJmTNu
LIDsNP1bir5p1SPI+VMkXpW6vI1XUadMLolgFE7tInpVtmQ7Y5COkeKHN+fRKC0a
o8zvOoR8qxMZsFXS/uP1leC6gc6XzZAYPKiOQZeWqLHB1qW5ppgDy6Ur9AVnPGxR
psEPsaEYXGVJ2J1o7a0KtmuKNhR0ZAl7CKB/TRKuQ+V678ZMIpiNTsoF3FmrQmP7
jWsyD2QRXLh2mBufYYiesP1YGhefhaXuhOtg/hlrX8lHy+dkzY5P3pcrHeSQRWQT
aFjxAptqd1p3CfqhXNXmkocoXeplmqYBq/11EQ2AuwTY69g+ZgDtxToGl0FNSUtz
BodqgH5bwtvu25eIDMp2HqPzIYJ11/zltp18/ReVGveAHvnrkBeooNjBfh7FRU0i
Ci/F/IPDnSjG7VW0fmzfUp6W19Vyev1GRwr/aBo4sdAGhzO0e0/jjHPvLJlDRWoM
g7aWPGDmBcZ93uUJtC6EFHxWObYXUvZEmLyx/9LCjAkXELwrvC167hvWPBxkphaq
tnjmttd0Q7B9/D/YK70pN5sScaaJ3Ob2wSq4SqHjT7QGVCKQyky7+WaA0hJe/oDQ
m1n1sTptzn8fokUOM0jzV0X1Dv+gL9bSAtKT6JPPTTN573Y5hNXz4XohxqJX8eg7
i198v++Hzf+nNnxLsGR883GZ1L+a3R0Bj8HJ5/GQDrjkwDEHAGCV/ZZD4DsyUfLM
rtKNJn79C7thOmJjTSjzla08Zy3l0/fK3Ilw/sfNbQW3/h5SkHjCCgj1ab8KtR1R
Qr3anfvDtiHX6756AyOWAFxvbv3xpf4SZeJwBpdE/7JNNsaUun2uOTMUBBHIvEDx
HWNd3d4c+oNZ3ky9buaqkzwLskRXDdoSybR9JCNUk/sZ2pZhLIkhADjeKsCCMlQ4
S8FhNDHFL9BGrPlG3HS9j/3bj10ExmIeEmCkCCit99al3hKg3fH/CJkbWCuVT1g2
Z4WisP6cNeggBNS+Okoqci1PqbqG9JxiaM4lDHUifVpG50Xc1cbUdSQKNgrWLbHd
OtRGpFfuWzdDrYEQRRo5QJ26twWQa+HbZjtcH564BO28vGeFYQP8566fLrUoh7yc
vQZRla9HA3Faed5f+fIYuk0p+Dj8yKk2uE0J+PuWqB1WtoUsXOth4bQ3qQJznRZO
SREXG6w++4Ys2HTw5ruJi4dhkKHGGklcS9hW4gfEbu+vgQJm9iQ03/T2NW4hs+Z4
3g/wZ40mAW6SZCw0OKX+YvVmAhPwRneArWIi6MibCTOe6gYYgtZ0bq+MZH6UlN+U
figAsNDeUQ7KQ4ZfocdPu4bYKomS/YhN5UzE8/IvPJv5eAO+hx0NOcxxgfnQ5xi9
LYydIzOG5k5hWrqpRV3IRUkRrE1ZdGquX5rc5QHKCv5++Y+UeIPs2+NWnh0XdPKC
6qUSbrhyieX4hZ61lgRFxiIjQzAP3w1LxXy6OEghxOHPeHZPR336pLMvr8A+bE1T
x9Tlmuyai+sa2ne9gBbnj8ZH7M+ez5YYMl16C/UA7CU7/uxHh6XgeJC68iuB5mo8
w4UstUaFMVgGCiDX3INPWs8QRcvWDnEEXaKUSRtjCDBQGpu5s5aGa7Pb54QspFyR
Oawi9+qM5gj7Ocq3UlAlqBMB/+80AIulAB66Hp/nIxgKZn7WIiapPTmrZBCF7H5F
zfzI3iia/I5uMPpWZEALPvQQNwrtv+cJ98XrpQc/GX05+B7IEbVUtuFTHghrQJSy
M1W9Tg1PKf1N5aO8VtmG6IaFnwyp90U8+SoHEv+RfOeBHsV2ZYDnFx30GlaarM8z
PUz/AE9q2YLdfPmqQdSSkCl3Md885+5Gg4SfrbQe5lIY61uDlXaL8OHS6sMAUnJT
Lw9HS+fiq1nZxl7V1r7KxLjwQsLZTMYy9jeBD6NnbdS+ZxCZ07BA+luC8z8hVDr+
95raFU+kQ0kjvFveeh52+OITvinLYeB4Yl0aRVC8nkxoIEwdl0W8bPjdUV5UZGi6
8Uvea8eXzBwCXBgmHQgCjfzbucVikHQpTUco6iuFpTLsRQjBD7JGgI+FxnLdfkZz
3Axun+y2FQb1DOVnEdvZRGRtFo49BMHnGiXgajM7F7ZxWave2R3giLUtP0zPGFxH
XLOnY39CskexBzAdWjf44iqcupDc+MrSNl+yaWKPHz3fpn19cow8JXfgjwxQvHFH
2a5C8fbR7/DdO+GlrnWsOjK0RyVKmmkKdqqqTglTvijoJels4GlkUofY/zCVOsev
PZNFHk/EgxCDW0NHKzHaJ8NFy4BM9+jwDY0/rnddRnh3kRmnGMjzc8d4r0PTDVTt
b14u5hN46pkzFjdIWdx8TlbH3anRLUIP4mmrU6wL1iulyjHdLRNFcNg4ETddG1Eh
gTamYAIMkaROPCNYr7srYRDr5n0pmk20DQdgwRGz/eV+cH1r+q3QAP9FvWkxW1H+
FucGq0JDOBRiZyKClUUqiCj6db/EKrYJpIBiCXMTKYrIroV4seAPdHEQH4nIWHJb
SsH4MOlREjBqs2jC+/R8wgPRbN7KSHUattZp5nQi6mBp+/8pl/Apmpawd5x6tHhn
FbGBsC8JIbzk2HAKy5+BR2D2fdp1XVdemn0C2ga3VI/V3xBdtpXo0v2gLqb6ai/G
M2zG1hXwk7S30r6SV6ldpq2MrsO8OC2kQTlWHmc429uU281xaNdXGKTnf66J7DN9
wpzSmzMytBzbvhU5+eBof2b9sxsE4GySNnRkoyb/hiIa1M+v1wa/PoEDMNU+Q6BW
5aFb0khcAmpWJO1ec8x8rajTipILpexLXJgPLdSugIck4fkYxdnFV3byf1YQzNyc
UYgyGbrsYTF/mh35tFK8inhnYN9Ui2L+JujPXrxQcsg+K+7Uln9AzLXKFrVGp6hI
YvWFmfIUUnOqkJrErpxzkZvy6Sh/dQepg2fhM8RgYMKASRgfcA1ghEjtNXkCaGo4
KTW5TYxs0WivqRewooVWJe5zWcY4M8MLPJvhGrZ2mIexfDmkQQwi0IvBBsLncMq2
dKUVoJpCZW4IqbnkcTWPmmoRsTyvXqVXGgC9bzKMevIWgZHnS6fzc+Yd57zsHPjr
BwJgu9yaRNAIdCz53lEc0cVrCSfrJomjXVlqgM8BNUibUVWJK3MM9dBHydl6tSRv
E3reBG73mL4O0TrohLFGzqM6LCaWDuFm84JxdbKRn6/5PLt6/mBcUG1M1D14NgNj
FGtRh9kzpcR88DBGPZKZgj+pzwM/uavagheuniMgQbP3vC20G/faMTnJVesUSraq
nyR3tEYQPBbKWZM15iUbtdBsI9fenl8BWd1YdyByyQVDodFTqLRQCKxAm00GNUhj
iQqIcHswJWx72K3v0X3GzSq9GWQtcOiZp5ty2sGpmbrBMKOFu7sJ0eDLDAJu05xZ
/r/KEgZQQwEBgNaJBR6Jfb7ZkM6EWB0pxb8tc+E2YGXX0wfZ1/rbXyJS4nzmHhJK
tI7xE/4On/ydJC29TJvHZ7fCKwuOg6ggwZzUeF3FWU/0ldZ/9t+rkk11etp3HM2J
j/Am1RVRjop2o61zYG2iykgygGy13wnKCfx07emsHifRPsQH+lJ4F/qwULklpeCc
pWPWxocyWA/P9qtyWGt+ZR304urcLUdU82iqbaxY3aYmWPJS3iVzSQXgorbc+2c1
i6vnH9Q+OXGQjsErzzFNUGLMbzcGZPjpVXiizdpKc295wnbGPaJUYDkQNXMDJ7B/
8TjlIvsHIX7RIS5+qYPSB69y80jUQrjkyBGDoM7MHJXz/z5/HFOnkGyOT73/6j3p
AJBN554MtuG1jtv7XB1pnnu0x8m9jCOHFg+u/f6BPktfntVyprlfBVtY78kzEHHd
89tQOHFuccca7Azxwxpa+D9m7Bgz0lXUi3LUwqpFn0th51ivXPZV2N6NVEXlNGBK
9DAEwgABMURpUFnDF4jD0GjsW/uZGG5mt6k2PAuMOIIjWo5S/imAACPYPl4mwkce
BcsPjz1Dll8MCAKkojragiip8iFStRSLSrJEvCWkENTqQ9MbRHhOWLy316/Pmqg8
8ynrWF22aK0eq+IyE/O2MeVGIB7g07rhimna1ctd9Me1kyHyNtgzvtSg+gOubeaJ
MjcXjjj8i1akigO4sXbIZv7zeZCAVpyRtd5zvkbdRxWwpkcSFiVgCNj5uFbWVqv+
csI1A5JAacYDkwcFR33lF78gsjZNPBhsg+tYeXVDR+G22vkbc+pFZICz4yWbZct4
T2Ua6tftEQ4bdU82FAppQDF3SUe7zGFbpZJSKHsNbPxjg2fV4R8hsGrZ6MdvDfRH
pdzpdzKNHxlei/tZgcAF/9cDlTEC3XSbLVq4hHgeh6w5yTxE02Y9wRS2lXu7O5NY
VCigLZj/aoOe3AoTIpccgnWipvMjxvlcSfKWj56GJHe8zhIbB4ysHS4qj+lrZe2W
7bA9a9WhFFhj8JmqXNpx71FvTmfDeDy3NSwQbcUpS/2rMOtjlqu9sHdTK0lmc3D/
kDKYPdeNvPEnqIelv/CtKS7wNQcdC9/SDuFH9pqgTOGrfGaWMg//+tI2U/TB+IVC
hbCBDl5NZk6lc8nDiii2DzsSNtS1ZqSNUH73H0xBf7pKY4qJ31fJbGucTXDPQ7Hk
NjMexJdwVfcL2YKemYScw9KU+0iYfDw9YfXDbZiTFmrOteHxERmV2ic5KQNnPPFn
U1sMWbjxZ624OgdUmWcioGe27VbUL4mmOX7zg/70LX4JrgKw6YSCkxvvTA1MCO1s
wdZwcRAhieMeulU+TP+Pl1Fip6nrt2dYTH8oA2NcvCwS/cSMH13pH88nRqoLPK9A
VD+tOSES3OvDF6JELGUqpXVK58vxgx3uXgcc5jlhlNZbDRm34kh2DkPpEhYuNy36
GGeAiVgyRo+akTyASXxR8FZQRQQPvdmJTbWycNMH78XvKw2/FNq8gGQE07RcdXN+
UdwLDAuzkbUQA20M4u04I47y+ikyJbLFCDnUzNsl56sfDCw1qcs/7URZ/3q9fEtc
EECtIzKcnHpxVlSpOl2ArSGPt75fvJMie+rgZTkXdXxoSgxFZ7NfRJmm++NFH1bs
g6UvCKOtMlO72+SukOII3yMZIiL/USxKsBjZ2EM5XU6twcbRTitzkdHoiN9XRwyq
T7k77nPB4V4Z03UOACHndClYGAx8QD1+O9Z9kTL5Z6cwtpfplQ8GHNOUDo56+Fc0
1q/S1n8eNYzekSbcY9Uc9enkqIJIlkgRfCqUYQ9p40WosU291XcyFXc2WKSIKsxd
XeuX0vB2G7ETBCM0c5uEO22PmuGK29iQRYgFNaAR1oDSBhhHxmiQZc1uh17dY33H
QmO24i4BzHO0KwNLoaCAG+ERgkSHjLJcSt4QhN/lntt8/O9GgvW89U3g4p0BjJFs
0CJo+KBzK9gaHS5/Cu5xjmdXcUQFx9QZeKoc6e3d0HQDPvYp/nTmp5F17PbTPwOL
kaU9Kk1qpxlVpwmdRoin91oRv2TjKwNaizz2ktBwxTmFQNDWlsST0PN/Qu6ODk4s
Yf4QjrgHQfT8V9tCnqOOwVyr+ZBd3AApbEXzf0yj1MFlf1ZAxw32xHYShQjS6xCL
XKdrzR+lLFfcQwPbdrB5GlVUJxXBGG+ctVqda73DWYqeyWaEtrMhZtHAlOVqDQGz
lq71KKmSFFfQOducKOB6gHyZ9xJqaYpdGoz8bx5CNQ9XHtR5NLqe/23JajSKVd9b
LoEJMwxYpNvKHtPIIL+EQd8QJmAnHPh1qJBKlqyCrGuZ/pnQsSoNQ86svHy3/nuf
aYLZ8tpxt4h7inCcSB7+J8q/KJvoWxlF2VwDs8imncfIZwEE2ImYa9TmJYm9Lrxx
FmLNseE4iQ2zbMPi3OHHaxCKxnf944ERY96YxMXbr9iUTORsCeCXcP+SYx9D4GDe
oOYyAuimVLsoKNSrPI0wxbZrLwM1KNEFlIQbkswY3km8NBAoga3D8qnfOE8yWZ6N
Mv1LGihPp6VpcQDPThUAWUK7b5LXGTJ+DVjrW8gHAysPnSPmHF8W51cfaJg9wtkV
hV5loxtqgWzovGz+ZOlWcYGatHpg44dkaJ8wU0hrHUYTwxIoi5TpOZuTks5rpNYR
5Vcb+zeENKTwBh032uR8TprArAQPbQkWTIdzR3S2YWh/SoNYhu/IIKab86Gbn3BD
8eXuPyEJlkwbJ2fNF0hpkGzmTcFGaNuegtwZrB23FjtojAnDYqOW78yLnAX6fv63
b2GQZPARqsiZxeljCSdyobin3lTs1/TtAc1e24diQKy18IClePrVYu3LvlALyBFs
WB/uUnjWsB3sFKy/z7Life/dOHelu/d8A4Px+Bk5EGV+/VGKoMMaOLkfjvCQ6joO
QeDeYk5l/7y+2UktecIRESIYAMjiqMtySk44UDCHc3tGO93JfiXa0loYMQ7qVyKe
ykZSghdZJPhfbrO+kzRY51Zw4m3NVYQJAFf3mZ4LPh2I4/wsCf1E2lXJwiTaV9Vv
W2p0MvyqrITjQ0KDC/V/i0OWIrVdTR+p9L9I9lPzwQRoRuDhVdYb9+BVFIn0pZtV
ZqQsDDgTZ26Nb7vFdEUg1L34ck2+6vyfR1G5F0FNwATJCxj1OEPOGXXS6+NDCIPW
IY7I7WwNFk+akOj0cqVNhSnpNMtf4Y7rC73GAclM9f0LYY3GgwxX2nJKTFvlcUAZ
r9jgvPqUXIECfDNQN+FZBWSc+gsvC8GZ0/NofojACwktBoqksr927w1MBSATapoR
v34P5fKJVchbeVYD0EreE/qgWeVegRksVMqsThvQABnjW6dejVqkS5PuAhONbRkL
YNEpWzIG0ITE/QT/uHQLnBJKeT3y/ia62Y/AlEE0DjSmSthfEPhJ5+nSXixLPPmp
+FypEL9AeDyZND1e4Bso2mcr84rwkWnFg6LUuZpzyoFsGu/4ridai/ga3F3RC43F
dp/miByVj+2eNVeERJ+mP891UFF0EtxxROis1sR0zFHuL/X7xcWtwsCml2Dn3yaX
by8puEVGZWjyM1C3HJ6kdgAjC5rSezWL80/gGmhzBOXfBzoGV+uz8SK4kdOrnFCq
e6tEgKrnHUM4D0cnrFmAf7YitgeqSXhNc+24M6OfC/eEy7d0CXKDpKrBY3jb101c
HoLBJt7tOf5B95HcJ1hzZssVoutD6K8MVPyeh2hSTVSfqUGhWmVWMZXS/bvayAQj
YtrVQWozugvNimbue1ovgKJ81VJTgAmVQnVQwwBx7pz29A2yijs2vzs2ptFVWw11
+Qd1nYCmoFT+frxoD8mOYmM7rC5ttuYXCPVu+DqudygDdGkN78Nb0jWnzzrd9Jof
o8+uJZJlpn7ytIMzYL8gO/kU0RQRlGd4GrPMNm/aOYCiRHtjzBB7AH5oVqwB8HqA
bNgCPk4tnns6N5DnmofYEw9VpLe2EyG/186K46AJdurEFmuQDUTQeXqz49q3mJft
jWaTxRoPdLTQELlwWTGDNOaucyGcSN7RZdFn/Y16NsipuPVUwL+XDS+cI5x134We
aPBM0XGEgQ34DqD+H4wd9k3DTMbc4+RJRge96EqWeJe/9NHL77R5h/lFmt2SuWHz
f2AtdSzkxZ4dlOjSxbrLm3/AEoRVDgMXqCfLqug2f0J+4FM/Cvuthi3SP6asSP4i
egy7EtZDl1tMgJmrDQQDXkbS0cOAGwQsah7ufG4hVAhtm2XXi8f9YK5KWVXEdG7M
P/UipQtazW60Y/BoiCfNv1pnQmQxdhkSW9uLBVMQhha8UQtUCFMp44o8Rck2WJv0
cNZJjy2/sA2YDpBBkcyJ5uqDeSAOW+U6hAfHvoOI3gVN4BgbePv5euATMdbE2i3M
x13XXQAPIlClo+MdUw/UPkICt88olk3XVOrMBTtvetY=
`pragma protect end_protected

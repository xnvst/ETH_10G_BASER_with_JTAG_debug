��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO��j1��X��;�-���c�qEhg��
������.���c�lυ�kBW�V��j"�3�UF�(OpKcD��х�KL�cZ�.�8&�i�����p9W$4�%��u3b5���N�J?�r�
�X���}H�E�A؄��ӹA�� ̡G�N@�ވ��neu��c?U�K�+�!���롲X�s�Ztqe��Gю���o��m�!�i��9P�Wf@����l2X�-��5�68a��X"��o�������KԘCnyj�^9�Pl��k��oD���YA�
��}�X7WU[5�g;N p��g�;4��g���/�?7��.�����'����w�̀��yd�����n��O2#��2Z�~B�σ� ��F�k� -gK�'������JK�}��X�q[p�,RE5\����aY����E0���U��*0�W Y�#����zXaNw��)�z{�/��u�Y�{9�TԷ�1fi�}�Q��wrW��
nQ��Ll ���X�]���wa��os�$��@���.)1�!���>A�S\.���p�UwwLS��/��-������ֿEm$Pj!�w�|�0���q��1B���Ad��
 g!�M���4s�xRN��G�bk�"�oi�c�;xr�ѕ�Ok^#I��Y$�䷑0N��{|��5�h�c9m��-r�3���}y&���K����?��c7�J"�YCo�:�=�*�7o���2/<�~ݥ�!,��D����<ڼ��S_����dʖ�H6����?E�EpF���/� У����m|�)����I�܃<s$��������rA1�L������ͬ��*��H䍛Q�����ˇ	���e*s��u� rl*��_������z����@�D���V=�#�lFT����Ę�U��GJ��>��>��`��>�঄��չnE��T�l�K����}]Fe[�H�W�������P���������gW��2�V_�x��;Qb�~��� @���]S��ό�7�_���&���Z��(��M���WT��h��~�a����t�=�FC��"��	��y��g�q�@Rw�GƬ�cܫu��Ϙ�+qmğûv0D���9;�+���:[4��j��[�G��;Z�v2����t�\���(R��� G��"�:�����Fj@�����e��=(������3�!��y�� ��R"�%	~[	ؾO���D�/|K�1�(j>[ȉ��&i���{��0V\~��4��2d3�E4.q�g�R@��3�Ƞ�`�1f��D��Gs[�m&���I��5�'�0�`<!���5���	푛���&���GGJ��8�a�?@%�"usch``�®n�>�ww[E��,f���0�0����6E��M2��if�O���!1G.��_K�5��㻰��~A�b7�ƏfB
��b��wi���7ⶌS�I�%��5��s۫čy4_�cRCi�����q�_�
dX��>�i��5�C���~�Ϊ��ǰ$��������D�|�����F���4lD҆��m^�$qFIr�^���K��R�=J�aQˍ@
,�^����$��*i*վ���V������m�������_���櫚��8{ZLU���}_�R} ���iA�*��*��<�
i_>V*�\�h����m�$3��8�����7_y�p# ���^����&�63��Fϫ�����V��Ρ b�E��}���$�V�S��p��``_$�m�D�SO�o��N��G[������ou��ϑw�2�wӶ[r���R?���|�˞S��}q�S肻Fxs0p`���堸a����-G��L�X���Ń����'�{��s�UY+�,�K���?���+��k�p>�Q�Jñ&t�����+�d���R#�mD���Bx�xH�*��Lvyq��ϙ�����2��I�w��xa,8I��%�s�a��	{�r�G}�?���d'o#ί�Ǫ���Di����U�!*�����`���ܞ TO���a�w�(��˼�2�d]������݀7�.WWǇח3���#�"�]�����V��.{L�	vŧ�4�� ��"W�`����Z�3%;�ObZ;&1\���i��5��=r��\!agW̸����XK����^�飵�!��h�����*jvL4^���?��k��/�0�pã��E�t��d���~6�J��CF��FI�U�Ao�)�VRJb�7"���O���?h�?���o`-ٚ�O��"cFF���qߖY�ԅ5���*=_����#*�k�I���-�Bb4Z]X9(ߎ�5(1��*��{l3��m�Qp����G�;=EmqNH�s�Ә0�A�xx�5ZT���eqZ񛠑����s$HA �}���-cH�{���E�M������F6��Z �gxu\"�b-�U?��ń��0��ef'�WW�u9��Ӟ�BT��X�.�W�1�������1ڻA8�N���%�P�ï]����=�y����FhST�>"R�"��y_fDj�b`r����!���sgq\-�~�5^�8�o�!e�qj�q[B\:i%�4��{��Ҏ�G2a�b�>�w`؊�X��[��3M*�Rb�GͻX�zX��!���/48�Ľ��"�κR�X�Z�t���D����^�.��<�t�
�1H)8�K��&��W�+����K;w�c��s�[�"��wu�^6%`o�R���4��Ȓ�j���,+�� i�}�
����Z�>P�8L����"�n����G*�-��G�-�va�9����F��S,��|u8�植M;�;�U> sޭ�ƺ��A�!�"U�D� �i�t����-L�4c��������贻q��3�';�M��Sʺnݠ�<͢�OB']����%qWj�qT�,���Ŗ�ϸ�q����j�P�����·Vh,��-�@��y�;�Vh����� ��Y�u�Q+�Y'��:늛���myQU��Ka��n�޳���J�E/ѩ�&��q�8o]�!�ң,�� WKZ13���O&�Ϫ�s{R/x�i���� ���ڼ���8f�5#r;H�nYͨ����0�<ܥ	59cM������2u��-@�B�$),o��5y.�Ar�`��r�c(�d�43�W!m�qj.@�/�Sa��M1����1��6���p�7���c:��:�TsRXs��)�C�x�Z�SE��)e��Da��:^Q��ulhGh�\��b(d�,6�GȑO�ƁP-�7T>nZ$f��/��xD�9u��"b˪e�f��ú�6^ΜG�]<F|Q#���S�ADm ��=׶�;�$©��N��
���uF��h�VV�h�߆�g�x���=��=��Z�<��qߗc�x�������t�;�k�*�νo/����L��-gw�����T�6��?���?9,ϥ!$�����Z���<h�%ڈ��������k���ڂD�&�oR���a���X����;���~t��]Y �K[�ȉ��e�����#v$wS�d�J�#l��Ғ�W���|���X�D��Xy���d��ũrE���.~O�=�����[m�8\d��A[&���9�M�w����OY[��K��l����1��{�z?�itX:��1�&�~�Ca41�bh*[��2��$�d�#�gy>�q��4m�gr�����f�Z��.�۴54���[�S��W.#�*<��E#��F�*U|���g���=~D�Ӹ�i��Jg�%��C5z��'��᧬�G��~?ӝnRiA�n�,^!!�3�%�����+� j�Rz�ԁ8|^��`R��	�rҽb՝��R"�n�))т1&l��+vhr`�Z ��L	!�6t:iH��amQ�n�$w��T�W$���������9u��<�Iޞ!�uz��c�.ؐ2f#X4�ߴH,*�@S@���K�O�Gz�Wz��U�e^��M��Χ���~�5���D�)&����	����v�eևԨ��L��[7��|"L�������^�DG�h\��^/�v1�gኰɓg�@D�qI��V�8�
�ʛ��=����b	�^�_QTke.��=��3C���ή莲�Ô�d�VeC��詚�A ݁�X��|��@��G�&�e?��=���A
���f���~�F� 3�<�୻��^��Wd"��a���vӃC� �'�lcy�լɪ���=��֏��&����
��-�!`KA�sN����n̨��)~�4�VJ���M� �u�N�⍽ہV��ÝV���d��?�9N�h��6��n=��]R
���W�Fy�)W���	�N�18�7�0/g乴t���&�J��>���)���Xsb8�����L��ׅ`�q��δ�@�=��3?Q f�[g$�ac�� ���Sp�z��M�X������6�֚=J�1�&�G��=��ƺׇ�9��kյ��L^�|�j�����k�Ԓ�s�FFI�+��[D���i]�f��Y�/'�P�����i�N3.\�I�FT��"ȼ�>s!�_Q�B���6m�0ÏX�τ��si�ڥh5FD*�F峴�e6f���n,�t�{��~�F���|�^���Β���d���O�[�ht�JK�e��c�?s$��X���"����ئ`��y�Y�?��_�[$�L��s�7d|���6�ZߛO6��/�������������8V���h������B�V�0rncs@�>8�|�?�X����|Urt��呫F�[�Z[o���Nk��2{p�4��@�����dB&���5I	�]-��ׂ��$%U!s�7��03Y�x7g��ܕ�;7�@u������Zq;����|q�eꕚ��V��\�2џ�{D1���$y�k�j�}������΄�V�K���G���V�Ӄ`����!��D�{��7�%��|�w	�h�''�I �fe�8S���=��Ӥ�lH���.���˕bbW,ޭ���`��B���0d���+x��\+|7X��nK��Z���&��-Y�b���l:��v���q4Ya�6����}ڲ댯�ui8��c$?=���WP$M`京���Y<$$��$����-� Ɔ]D04��ɉ���ǯ��a�yヌr�JfJ�T��ŉ*l���K�6^�B2Mm�D[+oG0��H��M�Y��l�`�P�	�HH��ݺ�#���A�ƈ��D'�f��KM;�M����C1�M�J�lQF�f'W�
�0�5Z���y�uf�m��vu4F��_�0,j&�ƥ�
�(���'0�����؍����m���q���vC#���}��$?�B�#�#7����V�S�^��]c[�������+������B�ѣ�}��:��NC�Le�8m��6�(J�	 <IZ\$ё��=��'�3�S(�mN.fo����a����UuC/����th*�m
�z~ڄ�*L\�%��~e��s�oB�9h��^���!�#)S
���\ol�@G���l̹�o��&@/񣩼P�P#{ ˢׅ��4��R�:���
8�_|�7�3�� �����%���T�(U���{@���bV��w��yƲ�Y����}yKߺq�`�2'5Ae�s"p}Q�a.��Fq�]�L=(5E���@RV���PD�'T)\n��lf�E�=ߔ&0P�� �u�r�t�1k����K�$����� ��1�8�D���PنjE��\���Dˡ����"GA�H��VD�_T.l.�*��Z.�N]�:G>�&�t�s�;2id���v�ĜUFA=JB���k.��a��i������<���G�BN�#�ܯ����<�����@�ǯ�X㌩�³��1�&�#"��K���-O�F���� 
F ���ё^C��tWF�3L���,�'��NL�*�<�u)[B�y�R�����(��f�q�n$�
�lVA2���1t�k�Ȝ]4�	Vpf �2�b�;�ۜ���+�z�D֤�/?K�TU�%G���dR�6'��K�&{L��ѩ|q�ў�f,ĸ�/2��ŝ0�$����K�͊#x��K�|�j.m�#9�z�^(%#��O��d*>�.��c����]�i��@�tF�7�ƴ�7 I�r�7ǘ@.Fd�!}�'C>��
�B������,!I{����Y(�ڝI)�h'*�����.� ���������t�]jt����j2�3?W��Cqģr"�#Gz�!}��$�N��a�N�_��19�?l��g/�R@�c�0�U�ce�P���۰�!�T�}cҸG8-�vq�
W��Sr�۸�s���� �BM"�IO�͠�h�nߓ�	����&�`C,O�q0Q��ۇ@�_O$�*�~v0a:�kl�W!���,�D��в�``�ϓ-7Go��.��ȖOU��gz*���������������������8��#S�]z�}����I�xb�_�knC4�}[{�ꉣ~�B-U�����cKˎ�� 7���GҨ�7�����7�h��J��AZUe���F�jл��Y(7��׶J�V��[\���I<W���p�;�)Y��ډ��N4!ɔ��t�%"��n�m#��s۰օr'���6n~�Gݛ���{�a=��
"�}��y hp97�:W������U�Չ��\k��a�z��y#��������>j\�*�km�X��A���ǔ��z�T.�"2=ҳ
�6�Q�SM���J7�X��ͨ8�Ơ�&mx;�f�9a��[����	�_)�i?�Պcy�33�V0� �6��^��逡}��r��?9$*�	����\`����-k�����غ_Ѡ_�3h��>���لA����3����w@ 1X��
��#������\A�Ƃ����C��vEB3�EfZ3��?�D��35�JD� �U9\B�يG�bO�\UȌ�A
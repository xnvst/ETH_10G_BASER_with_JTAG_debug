��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡j��-��l� �3Wʴ ��ȟs�/�\�Kڰ��n��T%�QjtD`K��R���S*�h
P^i��W��p�7ơ`�I���¸dm�	��E�������NFɋJʟ�k���*���<dj������٬v��ʭ'Q{Kl#�7JJ�\�`��u�4(� ��i�VV���Y����_ɻ�99�"fZw�&\C7j9�~֊�8��+eo�v�y�\-�h"�k�K��(M�8WT�9�۶�������BF��2�ԤO!Kv:�<���+����z9t�H�u�6��U�Nw6����Z��i�9�7Uh�?՚E���A�$K��h@� �`Fž�D�F�4���,^/1�I�d��mʚ[�>Q����۫ʐ|�Pv��JԨ	����4�0~x��Eɮ��PR��d}1�g��aMV}1�+)v9��u2Hl�P!�Q f�ā�!��~�|�W��R��y�d�~�(-y4B�l�ٺ����!/��=�7o��D�������[�%��]+l`{�;kTN��V<��!hح�A�#Yv?;��ד-}��4���vN���⍟����`~y�)�e�9�"��N��jj���\�Na�~�d.���E'rO�f"�$@�������Ic��ph$j' �yD��Y��������%d_�\��2|�m4(�����7�T�[��4��������;:��~�x(�+_�����x�;��'��	m��ch���F'r�����Sjö��M=�l�A�g:vZSC�-��a����1'�)2�`�vp�P�����ħ�aԳ&b�0��a<��RYC���h~�Τ�M����Rp�4c7RI��+�$"������_��mViU[����'�=�(͋[9���[-u��z'h+EGKnH�I��V)"��y�5�sİY�����Ag�hJ��κ�z��#7�O��pW391��R�j��"Z0������� �J����d��<��-�c@���G��Ֆv_�z��o�(c61�i��^e��^5�GY��-�>]���ʙ52�-�;x� Ќ�J�<������gow?3��N�0��������}��,)+E����}�曲-��)	-7kɘ/���d>4n6�&yi�yc��`.=Z��K�&x�/�wT������$��]^�E��:���K������G�G���jQ A����߂������~6�M��9�詉�.is�c��[�������z�I�;�ȃ$s2b6,����J���G�cHđ��AO��'�瑗�v����LLVR�<�'όJrW9�=(���k�΄HLrD�˃)]>p W�)Fe9�<�A���'X���ޓ�2����ͅA�?����pe��ɡ�����U��j.��B����Fn�,xP�
�T���Jl����R�ii�j��1_���w0�^Y�u�����Y��~�:�����દ�?��5x��G`��q�s8|}ﴑ�;Ā�̨�	Tj�ZO6�(@��U5�Yƛ �l�L��n����dX*VCɣ-�R���M�W�s��=�
�-�4xt
^(K�e;�_	<�*T�,��و����9��e�zW�2.�5#���[��C��Bݳ/_e+�2@*�~_��.r��--X��^��8`�����>Ȧ,�y�P���0Z "�	�/�R���>O���q>nĪT��^�s����}�M�݋�q�����ޖ ����z�c��F�I���kAXlo��sb6O �{`�>��j�8�z_�Qq�ty�;_
 �ǉ�^�ئ�8��3ڷ�Y����LfcQ�i���.�󔭸M�	��uj.�s�U%�U��Y E;�F�Wį����m��@���*�����t��)� �:sU��6�Am<����j�Ԣ[�9�y��[(�7DT�P5��b�k�#B���&�ų��em�V�	�_sr7+O9���3|L��}���~����;?��\|��ݎD��я��:�h(�9({=���n��b����kg��bG��f��J�tsS6��^���l,5��8:/	wA@�|�)�U�ߟ��9K�N{qD��L^Q�M��X-��*E�+�̣_BuqHQ}�#�y�F�1){��y."�Frq��f�����p����_��������ťcܮ���7�h�B:��[�d����f�EA�}�'���삯bY�ê�ɨ�X^�6%ZV:C���ײE�J�� ��'��VP/����~��j�w)���(��H�-!�<�&45Ш���פJ�V�=N3���PDC먺n�>��7�[���0�j⫴�_�!cђ��Ȳ��tB��t)"��ֻ�I��En���X`S�;
����&)gK ��q��nww��%:9�����*~%��j-8��E��w��N`}��ȑ��}8iK0��ZYJc��<`�S�^ץ}M[�����_���Jb��<:b��n����" ��M�&�6��VOE����C��4�����ϥeI�Jr�U��j^��@jvn�Id����=_%�rHwT��<З	�{Z�O�J��k[�8p�V��y>��u�M��q�!2��k�D'~��N	S�L��
�J���
UB��E.����w�W,��&�5V���'��^���I������9D�w�J���(���L���
q#�y��� �x,����:��7u(u;~�eYYƖ~� 4��r�NI�CL�9�$<�y���dmW�~�
/�p�[f��� ����׾V��7�s�=��.+��9��[@q�m�2B2��3�����[�A�:m����W`0��,�X���Y�:U ��o�C`�䤧�k�vW���_c	ƽ�ՔY��E\P�ټX@F�����A_2ap&d��V&��X�!�0��d�4�v.��遆c���V�.8��������KK+1�ּ�*}���g T:�=q)'�1G_���Eiό^m�i�t����l*�[z5�3�6���L�/�7�%��y~�=Ǣ�R��[{��l>�N��z֣q��m����.y����*8ahX��$�[q=nyʎ�|�R�et�B�&�#��E˿6�v�d�*���)���0d��V��wh�sDxl��ӓKW@�(Lhf�r����f�qt]��s�Q��E�y]�|:����؀T����ޏ� @2��_��:[��7P��R��|U���+̆{��>���u0�E:�V�c��g����9�O�/ۜ�p���h�A_�R�=~���!�6d�1~S��]>�P
������r�8\n�y��6rKܶk�E5�\��Q�1ye���<p��1���r��]Hw���M��\5�ܦu�wl���|<ܥ?���6
�Jd�
9W�����'<\W��*Wq���*韵)���}�@|:X[���IP3�P�����u�M�-f��cA��>�h���tZ��.�1G�Ye�p�jm���3(�m�i3�����C�/&�qܨ!�q�\��aH&o(����Ei1���ϯ�(�{�_N�8��_�Q'�-������o9��#��[?_�f���,&2���<�m���_�w�g�^[v����u���s�XX,�=���X�D�1�	����b���e,�%ti�_�$`�O��ݮM�F�lѧ��4M�J�K�&-���p�NG�{�=�""�@����6J����^��́���gwA��0a\����2e�0��@?hɛ_�����y�:]{���y`�K�zS���h���!���IH�l@vh�%��ڣ+5�Z�f�]����ӖO��>%��^|�>X���E��9PՊL��^"�!�q�f�l��_TWLg����hI�Χ�,"�é7������[����t�`�"���9���\*�S�Oߚ�ʕM9&����=1��T�B��`J��@�v�"N�r!.�?6?�k�4�� =�W�җ.����PԂ�:ѻ6����Jg���3H�\��-E7�5U�փ��f�ζVK����L�#���Ȟ�x��h�S��E0��g�O>��!T
����C�e�ɿ�R	�ra�bv��˧�i�k�
�����+SHHk}��&Q����'��VV����(ܞh�@]>I���P)n�tO�Y��hZƚ��j������jQ��G�pF&u�%����GI��mS@Ep�� �<�T��7߽�F�0a��	�>5H���2�{�ڵ�<C��dx�b��َ�X�L8M�?T��R=}��d�>?�
U��W���3�!~9�T��!�w�A^+l���G���Q+��ޒ���7=����L�+M�F�
�%�L�m/]p qB��:���A
�L��Wӓ�6�<@H�?�s��wa�#y3q��}z9����s�V��h��	��1�OX���Ǒ�V�����Tp@��Dt��� �{�ޭ��rd���k�QD�m_���ܿO;9a6��j��W�~K���:�P�9V���l����T��n�>�Si������r��o�i`aj��?A[�g���ˋ�D��?o`m�7(�[^�O]�7�xA�t�q�p%D�E{��K7MmG�X9S�����P��I��f��oe�K������k��ɔ��f��ۻv���(wn(�gq�n5pV}�����4���ұz������v�sk��Xl�?�%����ܳzT�{��#Cd��'��$�')�C`���������(�>��Px�;���V��7h4(�Ie��O;t��*]*�����Y�t�_�����DV��Ё�L��7���ᮧC���2enN��'JI�]��(˳X�����n��
������|��w�s-�̋�#��M�B��USJ?T���?��T>%С�MH������SWIݟ&4N+��_S�>d��udtBT:;�밟͍,�6 ������!�����$m:�.�E���F˟tУdҨ�8��ٵ�0Tk�d=Gٞ�Rcu��ت_����F�s�
D���<"���fLt�%��Me�v���!���b}z�m�����+��[1*�ѹU��=�lc�^�T$Κ��
����J�-=�{ϊ�G��ap���=\h|#iL���I�Å8�l��,F]�4Xl�Q,!�b$�@V*�'��Q.X��B���l�'�-�������3��.KD���10L���U��"j�'4Y�(��� l�;?��)3$�JL�$�Xlj+|g4�qV��ɭM�k{	ݟ�G���b5��C���9�c*�ہǤ �?L��hT[Ҽvu�N���g֡�(�*�ć�RR�^��9Â]�����	Ϊ(����v�Sv��1a�ʓe��
+��@$��Q[�7)"0`�ۚt�L��Ȁ��J����tPȔnte���������D #4+�1�8��-d�o�~����նϟ_'����9ɿG�6�9��s\�y��l�Jd��\�Ng��t��2�Zٶ�����c�v�¹�k���%=�Qq����႖�hgH"��"�h��Y����j賟ɗd�.���^�����{�ա����=��-��I��y�P�m�2�"�����Ӎ�˟����H�	���EO�n�͑k(Cb�����l-V�O�ޅ�� �ӟ,u0�	��|��ʎy�t>)6:�����[�^�NUZ�@�
6s�A�?��i縇���$g����&tX
�}P9Q��`�W=l�4�&�0Z�z��O�5}Lͧ8j�#��m
gm2�|[���4sb�Sd��az�^`'.F	L;�K#L�A�z˒�ik+�� ��m��&e���C�{��nZ��|w6�iu�w58X�f`��������#�612����&kP��A+􂕅�5�9o���Չ��$~v=������&�D[H�*���!�v�]r���q]��AFJ�V:�T{|�1�Y1��3]6C���#z5F�Ȗ��<n%��ww�f�� �?o��������`1"�����{��H5W��X�Q15�S�Hq�M�_�뷜��'=/�/��ǲ`�Q}ne���ʾ��� h_B�	�x\��4崡F/����^,�+�H���z�ug����(8a�tK��6�-���O]��8'�謉\�ץS����Y'�9>Z "?H"�p`��DZ4�1�Z��<Ln4��O���md9��[�$�M
��6�����uVە gC8�w*|g��U�9�+n���7�՗`�qH�Op�M��|X����'D
ꆽ$˭~�V<Kc�?��q�j��x�9Y�{���*��'�H���J˓\b�ZK�1�K��k>ߕ��'�s匷��r����@cX;��s� #��WɱP�#��� E�a!"XNK��pY��D�U�a�46?d��:Ζ�^2�ϻ�  �v�sO���e���!(������vd��9�n}8��&�k>�Jȱ�ԏ���B���Q�#�W,�@�ͻ�t��.%?�V6r�+�Ґ�-��Su�>�� ��n�G�v�U��lt8r����"�̜PI�2��pD|��,�븡)�O	K1$S�b|��ӁQ���	��H&K)�V
bߋ���uD��Ė��6�_0$�Z�!8�\N�����J���C:�Kj}�?�����2��γ��r��Kza�pBVT�A#ՁU8�#��+BmS�n�^-,�H�:���i cW���MI��WEnd%���1.L.t�G�r�Y�Q��Y���.�/GI���y���H&|��Z���pn#/�k�|�����=˻i�* K}��^ v����\�wU��g/�dz9mF�:�7���Gr�L��]��R��4&�@,D�DZp��$���m��Ј�dP�F��h��1���9k����q��X0��R6�
���(�m*��G�8�r�*��l)�xI�X�x���:"f������Ǯ�Ђ�E6Q8�7w�T# f�3Y�;Wp�Y���>P��f��⡠��ω��A�l�W_1�H<,1Q�>�H����s�؞�T
�"N�Q��L#��4;�s�$��d��:]���O
ڌ�+�����]�I�n>�g`����ܭwc`�z���|~���4)?����@�N��h�-'����C}� ��M�S�*��(\����8�vmR(��#��C5ߚ~���8��çw�����BмZb����t$�#d��^LN5������[�F��?=-�4��SC1'��j���&��_a��0�A^L_[{l�$[*؍6����� E��8#�ޓಈ�):֘�$
�"�x�2����΀����\��ߠ�'�Wl���˲�P�r�d� !m1�	Ӱ�'ăC���B����T�@|��ȭs�����Igr���!���t'�ˉ{�+DD����a�m&�qf�TK��i���.V��V�Y�Y�B˲\����B!Gq��ZM#rS[�K��y��(�Ƙ��C;�4��mH�;��+�S?���m����E`'p�ZK���G��o��"pv�ԓ|,���n�R����gGw����j|�謤��O�ǧ,�쁚	<?�P�$,�ϴH�Կ���y��xް|��U�Y0�rdk�
S��fV%|�>��An6vz���u+����H�2c ���ķ��88뮟T��״�-�, �e��G5_�0�Pg�'�����kCK�3�et]��,L]bhwZ�sL� �-<��ƐA���;]�����lu�W��[wU��7
�>��H�ͱS. *Ϛ=S�0?"�C�95���t�d����Bd�G�Ф���Š2���I��dVQ`X��N`N�`^��i�vWG�"\ ��B�o�sY5�N�������\��U�.p���8���`����� F+�$��WK�G�F�'��ߵ���S*JaHA�b3�`�Qg�ndQ8��RJrQ��@��)�(�jC8�4Y�Y�^�#;��Xa*~F3��D�Wg��P�.����E�%����Į�����%f�����9[78�����&黱���3�$i��W�\����v����Ǖ���m����-���!�LC�Aei]>�y�������w��O����J~�M��q������*B���'���b�
;%Fp�t�i��E���
�p�ٱ�%�^W�B�xRyC�zNk�'���?�v1{iZ��*Dl3ԧ4�&8X8�Lo����$�<s�_�a}��J�D��MO��K��n�� 뎜��=�Fk�|�㽟���C�K�}��Q"���w�hj`�^8�+�:�@�Z��}τ�k�VuX�ΑN?ć�p�5�	%T(m�c1_�s D%���4M4�=��,�G�����ao�Rk#5���?� ��?�����"�o�:%�bG�A�t��	�C�xQ�v�{�~�����s}A@e=�����,�ur�Cz&�T:H]���P�[-�G@���M��ŷA��z0�t������*�߆#(/o�u$!coNOzg۫��%$�G���_�zgs���??|ل��pYޫ�����3���m�XV�D��>^�\�0C����]�#��cc��� .�c�)!��^k��M���7gl{�)7� K�}>��#����Cڥ�NG��8 '��,.'����G�w�8C�xE�3��/�%�̊���`��cG%'[D�þ�J����+���G��R�D��3s.�e���r������?8ni��i�=a �I��ȶP����z�W]�:�(���_��	z����NL��/��Pu��M��3l�_����� �U��Q�_>+��nʳ�Xh��mwX��&�X�D�Ms�cTud�| o���$Mt�H������V��E�Cz��p�j��3XMH�[��M����c(TE�G`_܄��ڒ�|�ß�h�\K�r�����)�����F|��'��v�@=}�";��y�����W�<Lhql��6���r���P+-��ץ�KH=xIvQҝ�n��/���T��������1Q�ц9�ߊ�^�F����������%������S��n\y�KY�����~�ic-8�Z�з�o��+M�� �ԋ�ޞ����r�͗lj���R���\A�Mhy"�<<�tլ�)F2s��VZ  �T0UG�MN�G��6�}�ۥO��0��9o�+uh�@OZwF
�v%������.NJ���z8�������;<�+O���3O��};��X��?��t�l��� 1.��m�y��:?i��Fܐ~��-�wY^��Lm���,K�F�R��>"�K_�zt�tռ����"n�&��G ��e��o
����_��h'̧���ۡQ���S�G�!����|)_È�d-��(��d�p����H��jd'�ʗ(�JQ��m��t��.��G���K�\�����آ�!�ܯ�>#VŜ��>�A^�X���4$vӚ#yo#�8���Y�LYdI��#
����ʯb�~��@!�;�k���ď��B�'~�����z���.���ט}���fcnAk���Q&���)����I�u�B,�m�A��?���<�6v��-�hE~�sI��k��l}A�R|�P����+�we	~�V�P����?�5U����>��MLWO�Iv
��D�d��Y����Q�CfH x@R��Ig'=9�3���&V@�d�Y���p+TDb����Q�oP�tb/N�'�dR|�;���~omi7�t��� `=��*ȹ�ٔ��&1u�D��ȋ��8��Mn��|��I�b����g�T	��*��s��pݘ��L��H���#rG��ر:9V/�%)~8%�;��O&'��i�#ֈ�xf�$<Q!�'w���5K������L���;�����<���p��^|��^:��NZD % Ni������-�鯻�3�	O��^�����A�G��5����� p�B�OSL�EN���8����&�� ��s��V8%�JG�Wox+���d��Gō��HFro�<J���\f��R�>ub����U��;�O	�'��S+���X]Xѕ̇D�(P��JwRK�d�b厖N����Oxǽ-�j�p���dK�=~���ͮ�/�+�vQ��m��de[u��,D2P�H���=HT���'�aR y�>z��#o8�7�-�P����H�뭎o�����,M��,� �tI2��_��*2�x�[��\��ӊ�Vk%�,��n����k��f]r�F��A�����Z�� /�	�3�4���q�b�<�w�YI�Н���2��fύwr>+���|��,����me.��I�C1W�,�^��N�ܯ�e��u��"x���a
/2��{�rp'�mZ��9� ���]�!�Յ���ƴ��|�&�B����}(=�L5�mI�^����"d
������3rjfܺmG�ui%Rm�D\�eV��P�öO�}=\Q:��_�^2�~���̹C4t��/�v&�������] )[(嫿L%{/ג����� �n8�����u� ��ϐ)'��NόĀ?%�Q�pLZ_l�h5�J?y
0Ϳ�g	oS�
o�}o����	���8L2����t�<�zy���7l`g
o�O��/О�j���cG����cF��`�a�¡�' iSL��c����qx����vLY����,��o� �c�7������X�`q�wVi�;�L�ɰ�V����s3��?��}��Et0,�C'�uOǶ���#�0�ñ��VD��|����t��[�+�g͙��q��f�Khԯ��Z�Abˢ��b��؟.��Br=;��{��pP^�I��u�q��M���V�B�׵ߗԌ*��)��ȞɿQk�.�D�d��d�,�>�$��&���68��oN����wm�L;�7��a��O�&,	2wt�s�l�DCK`~��LhB�3�6�48���~9�?~Ύ7S�s���2��aW�$W5�yL�Ҝ�����k8��v��aqFg킯��z�|O��"Ӝ�+�D!�]�'��g*��� ә�_�s�?��zW���2 uI����ÉV��"��ˇH�o��|3,��=������[�pp[S��n�_i�VJ�$�a�5���OZ�����w�t��O�xMi����뫦�TPtf˼䂡�����Fw���7�F��{�ϥ��٧�T��7!^�V�Ȉ��=��ǌ�����L���$$!l
{4]�'�յ�F�JV�~��.��I����}v������\X5��G��Q��4��]8�1��:��)��͚o"dj̈́O�dך�<q�~v�J�X�=.K�(��������bV�I]�~J�ɀ�{�ى���e9��G��~��RL���>9*6p�rHEи�eX`c"9wv�~���b�o\��95�$���$�I��mڳ����V\���Lī�?1���� V2�a��BBY�]��O�l띁L����)��h���.C�<cI�$�+�G?q����Tr���1#~܂
���䨉�Bf�b�/k1�hAKl-�S�r��'�'D�a�˅����W��D��܏7�\$�2]?.�Cz��z�Qݙ���Do�]sbwn�q���$���b8T.Wӱ�l�zke�n�8X:��B:o_oLb�+�W�e�����A}�P��J�L�����
:�%B5��F�VlgR�~�ʹ�L��7f�.�_�%4���!{h�� ��&=`��T{IE,gyI5Gl��A��
��v+�4�$��~Z���x�Vkz���ȧ�ux!���F㬦��(�=��)�$^l�3륇VS�˽.)�ȼ�����hc��;�W�u�Z�|8Ds�	���|>��a��|�><-k��r"�
�����M-�����g�׼� ���QL��b�B	805{Nwgg��k�I�$�Ws*��+;FEv�&R�at�&;��<vʅW®��Fse��g6�4�藗��f�{�@��Xdk�X�8�#���m�^����cJ����͛��j��D"��9㿇,r�d|�6k�W�!��=>��Cf�.��=m&�9���l�w`��)�0>2=�ժ�~�J�M����>xTGx³���{J��*��n����R�%dz��i1�G��J�at=8���{܁���J�@��_U��#�_�}��U���֙YHK���0���<��X`+�7�Y
O}\��M@��IoEM40����z����*�hG��Ac̆Q:�E#��k��M��A��Lc�0�Nu�i麿K�N+ņ�{B�3�#��E4��+��&1Zb�%|J�?��}�*g�qZ��?}{�^��0� ��a��œ�s?��T�=���|��m���L"��)`<�$�k%�9�����2��V��������Ϯu��	��1�K����M�h�H�c��i]J��g�oجe:�B���c�`8�h]͂��i�����P��cr_RA;�Gߕ�W2F�cr����3��7<�Sӄo~�U���.@�T��3P�t��ÔK�D�5IgN�ɀ���"�����g�Xl�S=��,���=��_ے���b���=��D�
��+��̢:��;,�̡�lF������뙨��������{��CR�Kl���j4w4�|��n*u�F�\�{/�z��d�[������X��e�ѡ�x���_j��L�?��s�ų�n�d4,f�%�a��=A��bѿV��*�9��� �I�R�w2�X�-Q@W�}D��	[eN��~ɔ����X��TG���[�v3a�=Ц����"*��et\Tҵ����DJ<\�m��!YＫ���$�n���˟���C�~�P���#��ݏ���;_C�9Qf�[3��zju�{���S�"2�P���O���`u��#Q��Yh���8�.�I9����@)�{�*w�;E@�l�&�:�OO��RP+Ŝ:�!oP��K6ER�~��R��]�8��_BZ��D��08pJ�:����*��ö���K*����k���@���>�>�o���@ ��ʤ�iV�٨(�iAy�H��H�L�5C~l:�+W�g��h~f���Ӥ����*���εw�D�<���p��d*�
n�:@�9�o�~�I�C+�]J0������F� ��ajh�B���� ����#��f;���݆���),��X��zS�`Y�1x���0�=b
B�@�E��ԝ�"������}�n��b�ځ⪉x*���
3R������b:C�G ]C���Ru�R��;P��8&|�j5���"��� ��<��.�����!u��kj(xL���M�h0�	�%A[��B�Zy�}�ǉ��C������ħ�w�ύ�p+���C�!:�� %	���H�K�ݝ�S��qS��C�d�?�2����חzKvof4Y��c� �%�%j*O��X�4g�a+�3�X�\dM~�����P��������xJ�c�;Z�I�?��_�d)����:�/>��/3��=(+��n c0[�)y䫺Zh�8��y�2r�ǜ�>�U���EW5�,�k�	�Yl��-tLS�<,�o�[��5�1�n�S���8�̢�ls<)"�m<1�a��$\f�
{s�g�h��35�ߑ��"xZO��,	�����)xO��&УšhV�Ʈ��a��Eo_�O��3��|`M��Y��n�����ςc���8I�m�L����f%��"�����w�n`��{���ĭ�ge"%���I8��v8G�J<"��I�8���V�łh��\�7��M
�JV��ɶ+	�P`���0��Ď0v�g$Y;7I�[gEd��/�#��s�Y�Υ��sDYU�13�I�l����-"�`v�r�9�r�e����F(��I�Q~��63p��T9����9{�&�t�5��u��a��K��3��	J�*�1�+@}~/�VR�T��R-���%����4��s�lC�NL�MI��ôGʒ�k�})�`Q�Gb��4�af����)8H>�9�����exTH�_�oZ޾��	g�VV�:$U���N@���Q��P��Q����J�w^Ǵ�\3X�z�{�R��8����-H:�6!ʘ�
�.�.
�H��>w�ȴ�g��Y��	�6�3E�س�G��WQ�	�W}����_�P,�,��ɛ`�4�@Fn��E�%�U�`mj�@>�Ą�QH��j�}�z7��������Ow�.G�?��eA΄�ќ�ܶ�MU�v��3!m�rRš����eM�xuXnt�Պh��Xk;.���R�OMC�a����	]��Z���X�۹:y�?H<��S6����im� �һ�}����j�I�*�O(�X��{p��ecjz<|pA�s��[�Ssh�G��&}�K�o�V���Ι�8�kkUVj,�V� �g���/i�W��.�UZ5��1�V�������Y�'��e8���Y�Wu��HFֽ#�W��5��VWh	���b�LTq(!�
7e���Z{������9�D�Ck 
%1V,��7�C��ؑ��? ?k�wFV���#.���>��BW���a�oH�:��藠���f��u�@�Pm�';�c[w���Xށ<��d3}%�O"Nr0��բ[�� �Gű[���U�h�Q�B��#�w�s��w�a7�:��bR�j"�Y=	T߱�$nJ���(��q"��00�r��� ��%A8O�^/���(WFS���C&	[�:)���1_�
���w> �>I�2�+��Q��>Ĉ�ΈU��]+{�e��?�'��W�
�]��ݒ�"^�ɊJ���5����^$}<xlI��듑!#~��H���Zth+��2�j��@9��7BX\�YH`���V�Ƥj��V���YJ$䩊Y��wɱ��u ����{s�'.~^�,D��^�챸B���	$�/�L�h�=1C��%�[yhc��ra�()����g�1��N�_�w�yD//�k�]q�
��W���ۜ?�_�$O]�;(p$|5�-�σ85:��x��
Zt���f��.���9�.�,�H�D=H7(�Y#O��<��1��j��t`b#��"�e�,'�('��!��z�:.&&$KL�-'�~���@1�;�����|>�z�C,]A=?&T2XJ�Ob�
Y��̎����j|�t�T���j\�րo�3��.&4���:H\<8��^:��/���PW��\�F��I�n�\J?�X8 ��r q�'��$YE�����Ev��-WVl��d�z��$��;��	Mm
;_c��k�^5t���f�']����	�Ṋ�h�4�S�D@���FjUF�s_���;�+�Qe�Hz�(j��X\2�m�0j�����YU��d$Y�1���)��E:j��qX�>wk8H�RK��B{�v��L�>��#�8��(�)Ut�8��{LǹE�)�d�z��)܁�����7=(��>����2��A'^�YA
R�׀��'��Qj0֊�N�^�bz�K�Z�O��|Z�М�n�wļ���B��3��������(� �`iN��Q�&k�cщ4��"p��Q/�P6g>q�@�"��߱�����Xςŋْ!F�b��Q�m�d��"�"ǒ�r\	j�}:�F��g�wk�K�Hje2�M�!Hsc���ʂ�%o�B�jUz7��bٴ���Dp?�����cm�{��-∱�~ W�'��?�����Z�(��u�6�Ex�%tFs�o��oD�ԗ��z�cX,,�FQ����Igc���C��9�9�����ڕ���j����M�keh8ұ�B��bdn^��$��t��7�E�rՐH�u�[V=�S�(�{�S��iU��|q���U4�m��0�1��v��"`��%^Ꚓ�D5̠������;��}8�Pޅ�O̧�??����|RڒP���K룝��5G��2�US�k;���S����Z_�	�N+ũ,��0Qxz�{� �F�����ӥ��	�Y�P&%`+��ɿf�U���~����MNԻ֭?�"sNms�㱖q��%k�4ݺ��߄�Dk]��Sb/�p؂��^��	%�WS�.Xw�m>t1��,3�_�����$���>�D�X�	 ���^�9 &��d��,&[mQ
��7Э�B;^�$���*��3~��>( ֌��=�D������+�YU^�D�?�CvxPV��y��.(L��L�{���?OH���g�A�����im�
;H�qq�4����-ٶ�0��sO G)���i5i��>�����*R�ˤ4�Ԝ��ᾟM/,+qOc��[s���pg��p���h��X�-���F�<j�r'.�,T]��Z�W{[�I;�ϴ�b,��d�s�|��P�]'��޸(�������i��k���X	L�7�ԭ�oJ'�1<=��\�%qg3:���V�8��\aqDyt&�t�3��_�t�� �Y�lc��6c��(
fP�O�E��vU�a�TR������2:���bmvJ�Q��<��ܙQj)G.T����P���c���x0Dp/����2�4y�~��K�y�Z�W�w��7��1�@/�B��\��Q��C5_�rᮧ=q�T@�B�	r���F&����yu�(�}\4P��(�9.ՙO��yd?{U��0J3�a=�^A�B#q$l��˴�L})�G�F6g���<@�2zOI�Ӈ����("���Y 2�}x)�l���a��L��J_׶R׽f�]�(M�d��6��)3t��x�#���O�������E-�+�W��Q�g�֟+
0-�՜豿8� X~��| �Ͽ�2C~�_�{;���	J�k�<�`��Ԩ�v�daDN��%�k.��#G�ɥ64���؊|�Y.H\��Kr��o�.�Ax��V� 8��uy�*{�(x���	R�G�P�v!B5�y��vg���x�J#,4��*W�%��`��s,��I<7����9�zy!�d!��Zǃ�o����_��^�rQ�ǲ�`#�2�~qz����	?����$�5���ʩ���S?�ڢ�Hp	6�Y���N��w�,ہS���P[)�t�Q
)�������*Ǯ�~�l�A�mh���� ���U���C7\�=_`�?���LS>�uU� ��;����k��L�^�[aq����U|I]X�߳oFPb-f|���zjg��a0Y8~�:�g�	�Zj�M�v^ҹuw6D�in�b��#��Q�Es��#�2c2�� ]��������6��oD񨔄/tID�PdnC�{��]}� �����۴�����4!���~D�s�����z���3@7R4 }CM��K�C����G0`�S��\�pY��c����(���	�ւ�TH�Q/TUG�o����Z_B0*��\7�VLeo�@~����A�D��NS2x�)"�� �����C���]�,�.�z�k�f��g�Љ#TMLuBJ+.O>�`�.|��x����3�p�������
	���+4ø�P?�wD����,��];7�Y!<�M��eB؝h�K^���3翘�F�V���e�_�#�֡>�g�ieqxn�!6�fȾ��@�s&��o��Z)�b�=@A�UKȗ�2M��:�gUEJ*����42��Ξ\�l¶��b���GP�S��+�WI*�ɞ�(����ٽ������r��3��4%H�;\�w���U�+�3����S
�qT_����:3��*��/�v���'���w���F��%6꾨�xJ�_	{�Q���E��Ʉ� ��t�<�`� �b�|������������D�����?p���1R-���x�k,~�|J؊�r2kGp�tb�P�7��_�0�2Z���E��n�m�X32n�Œ+}�X��5G�}�H��B�S	MfMb⽥�F��%;�+w��aw�f7O�k�.D���'&,�1��gp�+c�):�޸;��C���9�����)����f��A�B��bg��(�<���������nS'�X^\Y�F~֞�ɨ�_���ۆvջDB��`���@t���x&��cs"���"�٫���e� �6��˒��"t���_��K���oC`�5~�)	���\_��V�HN*LUҔ4����'�a\�������st�
�q��X�`���:3�/��3i�$??��
{��;��|�pp���u��ߝ��-its���20Z-@������<�V�"%�>T��G ����.V�K�q�V������`��D�=�.�A�~̈́��2�y�dl,`�>J�;	FG�P��ߦ�;6��Ť�y��qV�U4D!�i��,�NFk�29��w.�U_���|�b,]|��t�1�x]`�0|$%V?�Јg��0#F��Ŀ5i涐 ��11�JXиc�U|�f��@�k�uc�ɂn��K��ߓ�.0F2��@�q�s�y��	$��y4�ׇ#:�K?�`�#N��dA��?��������-6�H��i�_�Mv3S�c2:�f,�JY��^��b$V+H���i���k��q]�@0'�H�����y��/�������0�L�W>����Z��P�1��M
�u��C:���t<�|W�k�3��u:-��Cz�M�Y�|�*�E� 㭾�ݤ��I;!:r�,�L��o�� .���)&�n�:�N�q���_��d(���TڝKqƳ>q���{sarP�!po�h�:η�l Q��ۉ��*�jqej;�8��5>SחM�A� ����P!��7��Z6�gg�l�V!�Yh�g���]�ܣ����q&�U���ſ�*��sZsڧ���"8��H,;�=��O��8����XuRS������
�k�aj�c�~l����S�׺�k�z�.R;�)\N^�b��ޚD[&��9���e@B��M��n��i��!/�3�=veBtr�>�u��	'��l�`��@����Ѣ��_]̓W	���Gb�� �$�E˄W��.��ȃ:�����v�;{W�|�#�`bѹ��ɤ�~@��0����d���M�T�25��l�H&�l��EG���ǳ�wzR/����ɂ��((z���WK��p�n� }e�����]%^�GZA�i���dd���x���5QS�zA#���������{��o�si��L�V`��GM��X��ծ��[�����+��}$C_��Ǆ	�/ŋC>��diE3w=�R@_R������rx�=�Ўb�{�b0y��3G.Ö�Ge�9c(�������'XX�u�T9�������SP��F��Th�mMXy,w�)&��?$��
��{b�G܈�4U/��3G�;�P�墺zC�_/���~1w��t��!e�2�_[`�l�Y�A����yl
��9Ie��S���_:j���A�sZBAȥ���P^�|J�}��@�Z����a����%q�V�U'8���=P�-r��%6�7	#W�#�;TkEʏ]+��+�r�N=P��������:��c�>������5�2'�h�bU}Oגۼ��%�z�d��Y2�_H��qOĆ̩aì)���u�?�]5��K��'3`����ÔC�OwQ�,�l��,TY������d:Z�2Ad��k-ZM'W�F̎o���p<�1���L0��s�z�z��o�G|H.�9�6���\[-$Sc��FZA���L\?�\6��M�+��7v��l�~!Zs�A��K�|㳴9���/X$��Ȱ��;�E^Jlv 	�VK�I
C)��)�y��q��k����,J¼9�0#��A!^Ze?#���F�Q�J�����ߡ�̪3j�i�Ǝ��	:�d��r���$��e>�5�5H`�P���7��l]���{�f�n7U���CoZ�C�r^�=pL�5�M;⓳,��,-{NK(@�hG@�2��+BR��R�j��k��a \������̼2ȃ�Ռ;8�
�p�����2*���ู����zt�d�H8�׽�ݿ����uk�a�x龊���픨��Ml�(UIX"�ԑ$ה�1���%q�tFK��Oi���2K-�\�b�
�ZA�7:�5�a�h��k�G�臂D�=�G#��md��i��g0�ok��?S�ۅh��� �������;E�e5,,����f�h-��.� ��{"�}�A��X
���Im��yK��tWcm�4Af_8���1!E	̶qj�	�'�hJI)
N��e��/p����G�)���ID��s���C���6&�#�>`�����͑��Rd������b��@�N��h�xLy�V��C����`ޫS�U��>1��/>��Mp@���1�p�8s"�Y��Qs�Į���B�uG
�u����M�E �	��.Ij!􄜃F巬�)ƩƘ	��,r���j�H:(���?�S��G�`���EO�D�{aN>|��5G�"fzi�� ��u���U"Mi7��^�w���{X�)��3#������Ѯ�B�rO�f�����ͩ�f���؎췔�+��c=��8�G��<<��Y�5�)��9��8�ĥ�ݵa�� �%FҐH�>� ����D9�˼�oAĥW����I��(��s8dI�t ����D4!�jãb�U�-kx�c=��Ś�h��7:��?
s%�����.2{��9���9��b��X�b2'8g�.�0����=SPqL �щ�J�n�6�~��T(�����[�kxg>�/�*o?���a�������X-\o3;
Y�4�l ��#�R�;����l���i�#T{ه�� i��A�k�� ;�_De���g'a��U��j_w!��v��֭�ohl�4r���? �}���U�9�(�&ĐE�����P`�o-I��︔��(i�S����d��[�[���谆�EM�z�%8�Rl�,�U��5e� �w���rq�?dCE��琕��s�7Ζb�����B�6�@zS�[|����޲�%�j�@�n#�l���	 ��7�,�`O��+c��bKF�JhK����;J��N�?q:�8��-[�b��!�L��4������f v_�U&�?���dJ�*�!)��[1��J�,��@�m���kRv+ݬ�p�X}���gW�( ��=�dF��03���C��'�s}3 ���z���<*d��j�b���^#����-��E/�<t��޺�"%�yU�_n~��\�`���=���S��H���E����_7�܅�� �^"��_(""��OI	6�ȶ�G�Ld�#�w2S�`Q#��VWl���6����Uݹ HK5�;�m�Ӭ����,S�Gm�N๕i����;`.#�7"9S�'�@R�h�\$��&}���ґ����֚9�G�N�y�Ő	��0�6b"N
:ν�x�n���~���"*�Ǘ�j��|\�e�G_Qu�7��Z=�R�ܓhbbC^�K��(�mG�X�tЪ��ܑH]���������F�8�άi�'� �sHi�ێ�y3�a��qj���@l�sHl����$�
/�Fݡ4< ��!�ƽ��%�^�B���W&$5+���R�%�xA�R2��U�o�[��� �@�S�ǩ9^��D�����TYr|��� Y/��_;��2�gw�\=�ӏ���P�2�L�_N�S��U"���Ll�R&��w�g0
�ܞMH	�D�r*쳁�&</5\��'�ÒP�@��H��b��*Z�g@�6J��N��ԍ�a%�j�Nf͹ɍȴ*�Ӟ�v���C�n"����\Yi���[�Gq��w)o��ڙ�Q�"\xo8w5���g�-cŶz�4{��!����ƂJ�i�X�>��<��6J�9�c�!�M�m�4�o>'�i/g4�t:)���/g!���({�Se8%Ļ奝 �'D�l
��C��f���p���$�xa��,���x�[�r��ŧ8%Qu��J\`�"�i��	:O����i�� �ʠ�Z2g0�2y�|��G�(ع��G�����ؼ
����C�5��_c�w�=�*��~��E��32�g�Q��.��_YZa����C��2�����;W)?�Q��'9l��㨺��p��Jw�Vf���h���{�nk��,yBy �)ѹY��9���Ee>7��G/MY���˶�l����U�R�(����u5Vɒ�z��#ʏ�;5�l\/�A;s���X�Ư��>8�i�4�N ��P�DC��%a�mF@2�UxJ�w!zמ�r+;�'�V��[�EUdwrOJq\�C��G�2y��D��K&C�TT��9�ɶ�&ۑ`/��MZIg9������[��aK����|�S-6�O,��2B�9�I���↹�0�פ�Pe7}
K�T�-�O&ܽ�Vf��Q=�"���>)�ѺڀxX��W|�L��M�Ę�:7sXڬ(ؘ>�n��x6pz�W���4����	�&�b�	��
�Ό��.��H�k�)h
k���N��������v��=l�'J�JI��]4�]����]E6�/pE��\FX���U�M��hф�T����TW%R"���E�[~�T�ﶮ�v�\%���d�]�g`U�~ֱ��ɂn}c��M"���9�b~�ݒ3��s��;҈Tc&���Y��ZM|2�1(�0h6�TpFyǧ�\L7�h����X�\����&{����ӅN��ʵ�#�UEW�9�҉C��F��:���ʙM�G�}�Nd�uhcf쥢��-��+��t��3����B���������0� ?����٢S�Z7.�� jbQ4�on��
p_I�Jƫ�3[A�<�����:�t��E�a�907 �9/�sw�)�T?�|�c�%��e�௿���	�ܣ�U稃����&#��F H3��];�T���]�,.e'�qO|W���$��ۊ�ٍ��x ��DEB�_R���h���E<"�,L���6nZ�@AWS^�=քu����:s�.)3`���Y�1)P;������=w��}+t�$2zC59,+���$؎��:���b*�[�/��XUw��"�<�X+ĺ>�1Q�W$R�"xD2��±��5{Ewx:�IB8���m���$�� �6���3�C��p���Upp�5�0�����#���6e.a����� ~�TJ�'�Oq�3�Ls6@V�T� 
��l��_ {`o�|N1�KJxބ��j�*�`CM�IsK[U��F�j��9�!btʒ�"�{nֵb�I�q� 0���F���k�P[����M��
�{���ђ��'��1_nJ`�X����91�����I������?Rm�LƬWY�k��0'�ˈ����q�ݴD�aCV,#Z��xd��_�`���	~�n������y��U`?�H[�,�?�o��^�\�@�=�:bd�-Q�+v���N�����Baz�����C�z���|6�C�����5z�*��U�	��Tɺ��=��m��\������8�%�KGۑ�D�V�S�hg�`3D��"
����~�>��)w���vt��d^xkS���>Ӏ�������v~���3�����EL�H�� �6no?����Q��{d���	����8�������2q�L��z�7���'��q��w噣��l��+d�G���%�~�P��*啹�<M�P0��ь��n��X�"����Qw�r�H���g�t��Ԋ��[���m��[FҪ��@ג2��jChMrYM��{���D�+3{$�]5�x��Tg8��Lp@��?���?�>�)7F��%dE�ʨ��'m��r�~����ǁ֒�?��4�A��J�tN�+/���P�`��-�mY��"jZ�i��;m�(g���p��WJ˦:l���­��ғ'�b%��?s�}(5\}b��e�g��HD�M��y���Vχ��'�*�m��*O�;�x������b2��JkA4%��M�������A�_���#6�	e1�8�̯̍�� �pz�k�U�dS_�s��^���?�#]���� ��Zg��=�"�lx�m�F/��봵 X�1��u��7�ɨfB��{f�L�^�7EDpeQ�Z�Yl\T7�a��tM��a��惐�cr���:�-��hbs\��ʏ��v�ă��9d���j`U�#*aۺ��s�:~a�}�N��+�p2���6`�^_�2�B�c���7�c��H�c�\\vB��l�7���X��f����Z�� ]V ,}���rotq���Hݜ;7�n
( ���sbAC߼n̳��QlE��;�]�;�)����6MF~���f��T����㸧L��C�+]d�v�?�f^W��VQ�ֿ�@T�%.m�3��qDT�-xU�?�.E�d�ލ�{m0X�U��C�K��um^�_a�/)��"s��rOw 7^t9"���l�|g�M�w�x�����r{��F*3�OD	|SB�B�0q
��|D?~��;���0��&���v��,
H���5&7k�#R"�Lة=��0��/v�r�s��\9���_���A`5���&�rÕ����a��t
E�n���@�5Oj]��&��N�a��)�TEl�;�E6�h2!��P���)�Z��J+�j\�"�^�
�a��@�+�}=RB�A�׸�!N¢'U]��^	�
��1CEL�/���I4�9q�^�������;��l6�xf�`�b�H��,�ѠCT?L�hC�(�����m��ҕ��-D��;CT�=�@�YJ��������xye?�:��X���eUGF�K�h�<�S���D�$Ö����W�ڗL��%������ƬŌ��
d�����N��ã�;�:����������h�5��xrAe�W�,[���>��)��YȁY����E#5Wi>�����Yh���mX���)�����^_E���ہ��UW�Q��0�KSX���#����=�� u���ķ��@���]�Y�����^��mutAg��t��Bh��F���`�%񠬯�Q�E�O����k>z F,{cX���V�q_a�$�I�ëTQL���ʨ�B����I�N���֪�Ȓ>�X���^_n��ӆ]�S���Q�Lj��/�ۈ�P<��-z���}�Q2�F���;�2�_4�,氃����0�r����Eqp�y&mȩ<���ЃC�i��g�$}ɋ�$9�ؓ�
��k��@5�;� 
�Hr����j� ��!�qГ��U�[�y��C"ހ��_����Iq<�N��#��B���u���'���f���E�1�i�d+��3��\۱���wM�S4e��}��Z9�et23�^O��".g��K��<o#��z X��5F��1�^�L *�d2�j>ɟ�p�ц��<����@h�2���� �(��v,%��͇��NF�P�S�En����q��N"�������S�W_��3��P��	�f��z�fW=�%Z����&�������g�0�[I�m���1~5�x�u}ىϔ�ٟ�@7���;ʴ��vG���srDZ�E�s�G/#e��aVR�^�%x5Ot�N��
�Ȏ��UӶ")@uO�������1,[
R�{]bRd�����pİ	��S��ɾ��R��J�Ga����\7��ѻ1x�fl�'�EP+�������ɘ?�f���>G>`�
H��x��]������.�Dr��4ؑ�B�"l�?�V���8����oC�a4��A��Z;�o�7�*��j��@��u�۔ӫ�����j@�%����M��%q�-cl�w^P�mɺ���+�v44(��k/�{�����5*�tcLm1]�g����u��Bܓ|��6?.iӒ^�3�����g`�����DM���>|�B���N�@�ݰP�o���+{���J��0��R�7B�&�#&��t��՟�C&���մIh����~8E{(ͩ�[zV:Uv:�L�]��QwN1��\��S�Y�t��_4�P�#�Iٸo��[1�'\�#+�2�>���$�Mb�#���u	<L��<T�����b�ɋ��S����#IŔ�2L��Х;+jd_.��&>&N�����q�_Syk>߶H~�aɠ�/��C�m\%*���g&e�1�$,J��W��xtz��v�4��l���g�z�6��O�z\�j1�\�+�E4E������]�S�%������7����yq،<����77�N0v���_B��\GP�N�L !�ʱ�7�`�{�hˇ(�G,w��|>�f��ZqX� '57���FA��Y����;lw��=��}��>��8�a���;"��k<��m��k�~�u���M8�\zF�x�W�̨��c�l��_�`K-Cm$��g�i��G�����~q�R��8���>(}g���N�2���*�^#\lĹk�^����6+��8�����Ҩ���S���+�2�t-����U� ؁���Y7"�{����+�w�Ǫ?%��+�m/���I(a'؈�re�GY*	�J��u�yU'�$�y�����<i��ï����󰌵r��m-��6*yY!�7�	�6�_>�C	����zǕ�&�0�G��R�zh
*8EjR5�p
?����ؗ��RZv,�Ro�K��l�$~��%�d��5b�-���w��/@�W|���>�v=�՜W^�{:p?�g���c�m�!5�F�C�����g͘,|uU��&*h8Ov����PM�d\'�b�����[n�v���%�]#����N �``�+K��x^�d+�>ɬrb9��O��D�o����8'e��!f����8��Xqj���K�M���n���'��
�,�NJa���DE��Js���_TTt4�dІ6��� X-L�$�.dKס�ߓl�RUC���.������T۔�Mr�_b^����,Y�v��,�s�cmC��g>pZ޴��n�Շ��؃��.���)�3�*V)E�^b��_9s2l��RH���}��Eĺ�X��t��&$��=���х�p��ʵ2S�o��s�>Tػ$���a5�R�eM�ʨ:Rp&�Q;
�}h���u^��� �ǂ^�v���Tc�pSK ����|�V�]Z!��ڶ�s���m���r8\E�azq3 ]k��J4-���hC�־e4lC���vF}��z���Z������>+�觰yG��4��陱m��]D?|"�H�W{�W��V~`���m"/����{X�ƶ�U4x���������3��c�M���4mQ'ᰃ���y~�w"W���kc|$�����Ĵ���9��߆�v�n�����u�@�R��Fu�����y� �(+�R���O��7R�D��O������>E�ޫ_,�k�k�}����e��"ǩ	����*��nD��������UH�NU��G����o�m�6$b�DҪ���p9ƞ��y�X*�b��7�a
;�dfQ'W�	����6F�/p6��p8��Ν^b>g�l/��(�/g���I��\�<����˙�����_�́=;�j7�S��],�N�XuWmLom��V�iW�̠�k�k�fŻ`RM��լ�-Mo~�J���h�Vn!�#T�֔�f�F��T��._x��/-�܃����'^�BtO9�M����	HzE(�I�c��7TC���	,��m5���~"؁%>���\z_��P���.\��V3�	��z��r!f��p��=n����v���%�i�olH��,o��+�
���=��2�Mr��4�Ü.?���q�h�oV��n��x�F+�%���3ըǬq���6vȾ��cqcGo�\���عP�Q��Q��q�����Xh4U����Y~'�(?��QJT���Z�cޛ�է�����T#���&�)% W;}ʤ�\A4������q��9�G�U?�5�z젔RG�ӌk���	��=S:� �D��}tP$㬂3���ލ ��f1*�_���L��>��v �JH�z.{	kJ��[�΋cO6I1g�#�D��0�Vz��$&�aQ8�R^��[U7�[�"�4��Y$���lz�-���G�4?>@w�#�}����8X������[e��҂���d�N�*��9�^`�cbw�����x�����6/SVґ���԰���fa%�� �;Лt&�7�+{}�[�rw��РЬ�z�)�a7��O�(��U)�ǣ�j��\]�7�I*q�Z �Όt��@_�'8��J04�J>�1!�{�K��+(�\ீ�'�|��9F�����ïU��N�9�m?�h�ӿkJB��|� �Z���03NZ�9B/�f��O����ݐ���Q��^A�����=G�<O3���u���ǋ�Ĵ�j$�]X�J{DB[�D�����L�!A�zu��,6;�y𠌷��D�dP��,χU��:t�i������?�y�bc[�����0]�\J�O����O�B.ޭ���%�eKOrP�'�_W��Sa�p�۳�c4��m�>���Z��tK�۾�d>���;�\�b7P�:��գ�u�g��A?e���G�M�sJ� M�U4����*u�_�I&�dB�%�j�[ZL}��K�g�B�ߌ�ђ����9��l�ٽfh�i��P� �eA������r�G�z�ʇ�ˎ�OZ�{JG^&�K;t���q�~aL�	���ـ�l�_�5Ic�&�ߓ.��e�+b��IBF"gԯ^�����$�y\p6F�W�F��6y�hd,0�������U$}�Lѓ� ����!�Od.Oл5��==���A�M������L`��K��fkԁ^��~]��n����	O�HD�w3�Lt,��L���?��Lhq�Ӳ�C�v-ߙ
[; �Z؝"���ͳͨ�:�n��D��[�,��$��u�_�V��[�Y��Ƶ��1���)��13H���R.f���}���3����4�c�>t&/�
u1��W��A��s"`��R��j��O#������)|D�!3�AkҺ]���<*��.Z��y�(�-�Ń��5��w����������D��*��FJB������O���Ł2G�ϫx��I.�Q4'��I�f݇-^ݽ��_�F6�|���M��H\WT�U��!��TA���f�s
��N������:ֵZH���, uxvpv��ނo��qSḡ���W�Pu߾�\פY�y,�S+ӯ}��
�Ph�H��'G��4Ә��Q���;��
���wPyE���#��w�"F2���8hz�F�s�|y��1�ǆ}�$�RO����&ͽ�i{CI�
��R�g��o�E�v1�v��q��B@�d�7-�+峉��KSg5�
dI��Q�D�����@)��E%!�1���3Ӿ�� �P�j�7������[J+��Eu��e_5&DИxH��ʪH,@�d�ԁ�`�M�4J�*�>�%��H���K�B_zў�($+��:�- ��1@�4��[����0�_�yWG萁dy��-8�ҍ:�� /e7���G�@��<�@����4�a����M�3�i�����g���-U8'1��ǧ)]�<-�8o+�JC�^��g��bB�YKy�ּ�����w��8��,��K;夽�f}�4�DN	���#f|������(E���h��<�>�O�F;�u��64㪑5����ր������q���~���(f�}+��{�>hJ��Vtj��^�і�efeZ���x{��W�������'�u&<�G�����c�'����Wg��GlU'��*e4����E�"���hHD�b�SB!�t�>�/~qP�����ϰQ}��n�Y��>*��N>��i�B� >c�7x��[�yx&\�!��ڳ�(�����{7R�鎫'�=�Q��L	11�ْ�9�&Ol��i�]LWyn�V�ۃU{G���s�8��Y>3c���Y�&d�:��Y���+�L;�j��Y����-'�$6b���
���2ȫ�{#qW���]� ������;�D?WGq4����tC�-}�Vգ04
�xr�?`�o+�������M�9±H�6��~%�э�	�e_m]�}\��i�����ns%�,��?���_n��z7as��RM����ۺG��S0�&].O����'��E|�=�~�bTs����3�m�B?��y��3�E�s�װ w���/�h L�(q[iƝ64��1Ǿ����ո{ ���
@�+��w ��w���������go}�)��)cϾ��v�W��v����P�pO��%��'��$��d�I/D$y+y�R	f��~~f�
Z"�A&lvA1By䣎�&���X1fM����Z��\c��(�R�R̊� :I��T�X��Õ����X���������!���^:�NΆZ�:�v�R��>Go�x��bG��Lb��"�6�G^�[���ZR>g�H���FSΘw�3v�=b�+��}+�._ϱH�V-�e'��_�+H��z4��2C���'�r�!b�J�Ђ{ߢME{_����E���,��Rي���;��I؈�n�hԏU{ЩN4Ͽ�{8�� ���Ÿt�.H��[o�^k�ni�pU���~�<�T^Ul@U�[��@�I�r������-��31(�Hib��}�Sn6��iDŵ� ��S\� x�	���"/��.T`�pܹ\�c��f$Q�B�˨nWݯ��B��w_v��XD��i��g��o��Ӫ��@~���ͦ� �dI'Z`)vnN��E�A���_o�P;$�zp��qإ@�����A��������T�T힭��xl���X��a��E2�PѤ��,̐���9���=��<��
�o�sK�du�i\�B�)��~7G����ʬ�^t��X�&c%�zl'/v�GG�uCc=�a�I���.Â��V�(DF)��`�-����iy�0����$`*o�H��e��+K/S�� }4co��+��7e�Ɖ-�%@kn���H���m�#�p2!�I(Ƙ_��i��]��='�7���,�3�R�����k��ZY.:a�0�ǰd��1��S�	����C:H� W({GQ��#l����#o=��la5�Rō���P�S�?�����Fl(���}���d�����?n����:Q�&j���tt7z���qm����u�&S�bU�᫅�3`��)�-_��4�у�ۂ�!���F��|오�������˯�~�����'��o�牧i�p{YU�D�0>Ch�f��kN�j�z��M���шX4:1U(�D���")��!љ�0϶�
�ģ
�*�l���ck����#�}�L0���%Um�%p��8f�)��m]�%��/���z(��:�^S����>Z�l��#�e�p�����%w��#��ly4�����u	�rn����[x;/h��9=le�_'
�,1:E�{��A�����ht[}Oj&:�`��2���_��F�E2E�0�B����-��i�v����LE|�����M<H������w�5U�2E��m�X7\��A隟Uq��`�d^�ş̒UB�����*B��l&9��B�M�ڥ�t����@��=U�<x/���� �k��X�ho�*�C���T�:��"l�Y���8���m����(�k'����p�s,����̮'!3r�a���M������b2���c�Æ��d�t�L�!An&��U�4��Y�/k��5�H�A�j�U��|q]��j���ϙ�FwZi��Ə���^i{�t��n�l,��@���#"@}�<D�&&Fq���N�sX,���+�nQ���x�(;;�<�h(��!�s�2l�!����e�)p7�
?��6rt���8�Dj#�Ag�挔{��C�b�6�d!�#֔3ۨ`w!c/�<$`�n��W�V�lhMU�2�>ܖ�1{(_�{�"Y�4�rS���KJ�s8�b��C�l���ڼ*��O�*]�����T�g���+=�-* Vfڟ��< �eyԐ�%��T���e�=��h�ך뽈��}�j�|������WO�%Ί;���"@�&6z�C���w=���I���=���bF�b�+�b�Db��߹���iiQ漊���@�+]�-�D��X���:4}�X+���%fho��
L���5g2C�H���o�\��R�1yb�xk�;&ےp�\GS� ��YBzC��m��8�G[k]��U�_P�m���j1�d|s���D;ca-u��w�)wz8�T���;�ؿe��b=��_O�(�"o��]��BZњe�w�<�x� _��#m]�ʶ���D%͌��=}��G4	�7,��!i��s/+^S�|����M��:v����l�j�i̞0�V���fw ��^~*�$�M))���"�u	�0�%�	���l��u��dtsX8�� .�O.o8��$D1=�3U��ʑ��޶��uʁ�o����t�n�n��EEd;�� "����k툻qt�b�e�|��р�F� �vR
L�-L�i7<��Ƌ����/�~yT�GXQ� �ӡm� �����p�]��I�&�=� ���"(���� c�)o��K�T>!5�+��OH�nq�>4�(s�I+!�hQ��k��8�]����C����
Z>���ϤT���?n�Sw��q~�%9�����'}+�miw�H|� ��=����G�xY��
=�.����"�8Fx�,]��Y�~�=����݉m���؋��Λ�?ѐ4�]�H�&�;�d���ίIeI���Y<v�[����/��5V���n.��Q����o����h��k���mx��6�q}��p��Gb�a�W@z�&��#�4����v�7ܻV����R�#:� ��3�����Q�y1`"G�Q'�@I�;jq���SJ�"�-u0�lg������k)�#<c_�h���\��"������RlA-�o�F6�oy!]���ê��g�6a�=dm]�N6�'�� /��v�Ŀ8XV���̹����0�3�E}ɼ�E�滜��kӑ�1$À�s`+_��������m��Ի�@~7:&e�=��;���L� �>����G��Xs�%
ߒ1�1I���fS���5�}�]��:WHh�@�m|��?��P
UB��v�ɶz����h�d��}��u��c�ȶ5��ț�s�k�%�[k�:k�x��=��!%���wGs',c*8���<�%�Չ�0�3��4Ԑ���	@_Y��K�{u���аS+>���ב�=��.����
��S�y������n�c\��-Oשƥ��be�ecJz�*���u��)�����g	�z�z�wq4>�\���*�?�.s@Q��F��?��L1;��5	�8l������ ��{�|���
O���{�!���H�ħ�U�``�߽���~|�.���T\c<Ф*M4�� -W�pr�	�e�ν/3�p�mAH���5���f�
���x�:�E�:J��R8VGE�S����g���@��5�'B��r0��H�u~t�Θs�O%mII��'����ʮ}��_�cC�;7�Z}N�<�D�;�,nC����2Av �~�����_.���7�'���a��MY|�QϦ�1�,�!Ҳ�+��H͉T��T��Z��v�_��	2^��<����ǒ5��[�������:��ع�Xp%&��:S���)z������.�=���
Ћ6���;��c�-�ȡq]\�6�߸l%�s��,�1��`mhSCg`�dx��?<b�g:�����ЃF�l�J�I�w]@=�q�a��Y
������I�*(]�P�#f
⚫���tz�{$j�~y�j�e�K�--d����8U�	ε�L7R�l�-��!Q#����L��]��u�Z�~=�����y�YI	�Y�N"�#{UZ���chFi#�x�C�uX��c�]���2V�n��f�9�	C��B�?o�{��ni�Ĉ��gi��������/`3
�H�+�W(��Ą猜a�60%W�w��Jo�;"�w�T�`����d�{
h�fJc���{���sg���!L�f���s�B��9U�`-������J�~����M��)R��(b��P.`��Zo�����Ej���)�s.�;Q%��{�z@� Ⲿ�Ce���0��ï�9Ř���.!Qۣ���,��i�T���%��X�[�#�uul�8��(�5�l굍������k�6�O� ���x����i3V�r�#B��	�Ŵ�R	۝��ɠ�����DH�$�<�	�Q��	�p���b<�x�>e[RE�2ۀ�5d	dho�"����
�lL���pN?/~*3�*�%���g:�cHA��H����_�v���-?яl�)��Q]�S�����y�?9�ҕ$�ߠ��(q����~�������Խ�ߋ�.)?��_
�A�y�-Xj�pH'���^���ͻU&x�9�ژ�f����8���o㮤|a�}kՆտ,�H�j�1�L��lvKI׭D�~���3�*S-$~����	�ټ&���k���q�6�\eE7��5�괟	M�K��[���|l&� .�f�v�FZ1.�s+I*�_� ����*[f�Z��I޴+��n"������e3���e(猽b�MX�g�u�N^�4��_@�F/:���{43+�y�����,�ʌ�	�Sc4N���g�XQ����;pʝ Պ$qE��n�2r��Q_�lz�$���܊+��܆J�O*$��e�q��\�l8����i@}	�-]��tYB�Qð�M-;����L��������#�5������H7�m��J�a0��Mq�:C�LN�kc�?�a�Կ�e���mWn�.p�Œ�*;�ϰ�x�2)f�.~}[�b�thİ���� @���ؚ��DB{�]B��]�%3Ÿ(h���9k5k ����2b�����M��������.��֫CZU7]���t�.�̭��X��!m����Z ��9�ћIQ�9c�U-^�%��E�Z]Ó��
}�ƃDtO��5�L^arR��G�<0,� ���Nj�+��u��ن����>]�ը��T9�x�O} ����VE����"��Ӥ���Z�M.��zy��3Vf{<؉k�u�	��Ѝ�>BS�yD$��5x�D)�����3� E�|D��E���=���hx�cu���gNH��/��L�_�iFy9ͳ�=.Z�=mrX��G���r9u�r�>�f!���6@*0�aA��q�{�jۥ�_ʐ~���"r��)�y��*'{�|L[@�f����8G��eԜ��)kcQ���st4y��d��:�|�gjq��cQޝ2*��3oU=-cH6�(׮��z�-�(�B���r_�/�~H�ܽ3��e�G#��f�6�%�����43�b�Y�3�W���^���j�<�M�}g8N�/��b0a����!M�>tgc�xi��f�����FCŖs<uX#����Ɨ�"i6xJu������k����6�S[�0��%�=��.i�DAː�<��!c�L�����Y��a�b�4k/����Z?2B��>>���	��j`�+ʼ�{�af����'f��uE�cc7"�Qi��
����1Ic>�o{|ƛw�9���ޭ@M��8��5��={I�^��*a��D�T���*;b��3�I:\L����G#�6�����>4���l):gp��Tt���5-�&7,���1���`k�<[�^��ɍZ�i��E�{�����nx��?�0�pmZ�<a��Fv��"oh�v7$#N��7��2�
A��W|	��lj��A2�~y�7���{��~}�AoFQI~��
?ԃ�2��Õy��{��2=�l�2�ɔ򁹵�V�A�í`�U<�o�+uw70n���y�:�����*���026�W�7��%z�b�z��b!zs��kY��6͍		�)ԃyt��n�es������9�>�`�H�5o��'���P*w��t�
񅿧E�额)hI��;�;�4�;z�4�\�Yo�)��k���b���qeh�Uf����3�����t��A2H�b?ӐpA��U'�b\�!ؙ�"���]~!6���&�FH�25^N�s�	���Ʀ�c�9�n��0�F�HG�8^������b��ZK
<SP�)��T���!��0�|�|쪆�}��ӝ���M���dOx�R��M�,boQ�0�
i��Mj�6�R{�scZ�ۋZ���.Kt���l1�H,�:��0����!�I9�}j4���m]5��
R�7��cy��$���A�sg]�R�D���%�r�["��$Jm�w��-� [�\��$���*��s�F��Ưĳ�b���qЃh_R�CZe�gǈ͆�+��2��˰<�W�_� 12U�s��ЮD����)�m����J���W�8��Dq�IpE�����B�D G�{ ��P��L�G>�g�.�ݰ��9}��Q���������X�>q��\�R$_�P���+�^��h�����H� *og&Rlt��Ii��3�O��u���kc���������% ���h� -2�X�f2�����F���D��p@���g��t�� g��LV4BF�����~:f�j�3���*�7�4�7����u�Hp�L�S��Vׇ#�g;�J����[(��3̢��g�������H����_p�.в?��|����F^�6�%�tE8)�+����?J�+[d0X��
��P�u���F����6�\����PdG3�h�~��_�U�95�K3�A��©ʳ�{�m
=��`8�w���%���1
����Ʀ�l����E����b��nI�M���-���A�����~�<���
Ǥu���s]u��d�)��{�`]���������֥�烃��
g�t�h-5D�����<'�sp�����dGoLE����q�R�x[;1�$��^�aAs�@�ӄ�맯@�]��I7���a�Q�h܉I�3�u<E�sԞ��� $�
jFhj���}�R�i؜|�g��2q���a)�U���I��+#H���38�P'��S�N��.��Tˇ���72�)�?�:�P饈�P.�ҐC���t���꾞�
�*�/C��[���?�QdU{zs�{�`4�|�o�.o98v�#�;�Ӏ�襑��^���b��E���9�ab����5�z��G�
Fw�g�X-[j���	XpԢ�`Ѯ��&����U[V����!IH8��	�R�'���}���:1r�qCY���BmXH����dX��G���!;��14x�+�&�7�H��
� �����(NŠ��nK��¬^�8��޸�&Y9صM:;@&
X�Niz����0�?u��b�*�{����&Wރ&�&��<t�ӆu�@�l$���@�5��ʞ��b=��o�>+��;���x3��M���na#�>,�DO�Z�|h���@]���o�gs���%�ik ��Ih��W�H}��'����#<���Z�DHߊֈ���s�Y�".�Oq�����D:A !���"���;F�����k6�v~�cm�*��n. @����l%���8��;CePz��~�g'�<7�%8��.�#��I�댶���,������A�uo��zs�J��SK��0���N�����,l(���+J���
���w��/��|כֿݸ�	Oz�"{*\��Z��	A`�;�e:"8��VE�Դ�4��/l���Knf��4�!��,Йh�N#�<J�{ajv^�F�=j���	l:����Bȓ]Cwoe��A/5�
�Lu@m3�.��[�Щ}��pMٕ5�,����{��NG$|#m�SM�̿D\}.z��JO��ʥ�	�+�v�h	�ѰG�V��ɃV�����lV�$1�������9�9B*���!�y�������:Z��0� r��X��������_K�2S��z����&=#>%�����{�i�}�x��Px����B��v�����D5���󬋚��&�Vx�?�_FwDڛh�:3�{��z3�5j�ѱ�����޸f���O��[�BXq�P� �^x	��;���R��q���5,�����"ũ}9�4�Ko��}�*"���8�5>eH�x�
{���=xp>�?<�F�$5�6H��iߚ2�<>�$Q�ίc0�@��xc*>P��y��}[+u�w����Sv'�bC�Rݫy����w��aU��\� ia�f$S��C1�
�6%���E]Y'�	�ϛ
^~k/�]]��� ^�T�/o��s
g�����}�cj4_<{�L����NB__B!��g熆O4D���q��v|[㑓��� +Xɲ�so�-�e�wN�W�J��]�*�F-)⒯��+��bi�����	����«�E6�]{�Kc'���@��W��,�����-�)?h66�.x�E��9�jN\@���}��?]�Wұ��5��}����]W����T��y��b�o�{{�K����"���W�|��X��8[[t���R4�Vȡ|�rH�<�G� �[�Tf��7/�Z�8���]eɇ>�.� �؁��ۼO�J[:�ٖǪ���kK~B��F��� ����`���*᫒�u]���ۚ��_O��9��E;� (��(�_�"v�ntl3�B���4�9�o�Z���D�yߊ�"�ߩ���(�E��!_Ҡ�v����0��:�=�#��<2
��a�����`�Z�J�c��ԭm�Ԗ;�m��1��@��h�����Op�D�-υV��?�*�W���?�����9.p��|�"�%Z��t
�ؾ�"��)D��=��q̀M��54U9��7�9��O�9�n1\{��f�'����	�D�vG�7U)A!�(U7S���$D��HP�f�ׁ%��/:�m���y��N���ґ�b48yp��j�����/��p�3�_�p4$�Dt�rŏ81F�+�<��@��������0F��O�1�LK�E���v�*l����w}D;��JR3�A�Z&�y��4)��~�,��I9�vR����~=�]L_��ʬ��d�V�r���8�74Ȫ�Lz���}N��>���æ�9����S3�/��;�u:R�Y���{��-����ê%�����x�U��R�S��R@[�tX�wV,�ӑ͏A7m���Lfu�DM޷q�aE�=��q��q�����G2t8/bz�m���ŗ��s�o]Y���c�%��x�ƅs��:t�����fdI��'9ni�)���+��3�7���,�iYYQ���K���]���!�4(7���Z�X�#b߲�#��e�Z��C0k�V��E�g�|����R;b���V����%��2CbEq/�IjX�ڕ�Jq�e���tXT?�҅m8D�٘wy{|����&��(��e���)��CF���/,�񝲤:klS=߈�W<H��P��Fd�i�Y����r%�y��Cȅ�8g��Nk�S�4�E9K�&���>Ê6z�)�\_6��4|�&�uub�'�*�r�aPc-ߠ�M{�`��q�^���%�Wj�n|��*��ސɓq�b��1��!��xt�r��#
@�G�^$?~��k���te�l`��W/����D�W�I�X��=�,��}��[�!ڹ����K�������ȼM�t�jOW��∧`q�����E���z�nҮ���|9Ev ྯ�~C�W�:��$��@$�Ds�e�Ʊ�*6s
�����ع�h.:(c��<U21S�~_��@�V.�֗K�{�i��0זּ��W�� ~jF��Z��[�H��u�@���_��[i� ��V���-M�GM�m�eq���|�hʧ�K��qfʟd*س^i,�
�<;�y$��j	ޅ��J\�P�0�� �eydO���x��|mI�/���S&V\����4����-�L������H}\�9���;VV\�Ğ�Bʽ�� �/|v�1�a	'ծ�v.���:��n�q���@4��s$�P`[4�/b!z�>$��
�LZ8��Gϑ�6q����3.��V�aj�_�+�?����B�Z�Oc�e�@�_�^����$2��P�J������J�GA��e�60��ޭ5�0�Z�"��z!��$=���'��tCm$b Gƕ��YL �=�+��O@S[����>#�S��KD��qK���5�B޷�H9aN5�s���T�a$��, ��������/�L�}PAxVr��ҸT/@p�*3��6�p �C�%OB �r�Z�m�L�AT/�[��?��g�z2�҈4�m'�C��y&��n�\)������r�#��C>xVi�������$P7ƶ9Ⅺ;\���
���K̫*�iMoį�ԍY���8L��:�|6��|�nC>��7�C9Ŗ������P��6D��z�z){�.�#O'������g��L�=f�)�<����JC)��Kx����9'�aK��X#��V����G8`���pw�v�n�!%臿�3�´�A���@>�5��e�������:��sa"�� 8zGp�� ������n�O2LH��l�\��T���E�{��VRF��u��Y 2X~���ʢFB-=��> ^��yRK�}��8�]�m븑uUx�3 �Q�HIfC���Lk����V.�~�"1�*8��9��`��71�J�K�h�M�e���l�ּ���?���_�hX��&�ڒ&j��ΛrOَ�7lF->X�f�Jľ�ӯ�h�m(,��48��&4�( O�
�A%��X�,9�1��=Ԓ3U-�zYx�ȓ^�Xر��fW�NV�Б��Ա����`�������\�1l�T`����ֽ���&Z���ݿ��i{?��2k��M�-����N��azܭ9�X��~ҳιW���֜v���7�cV����SH��h�Lz�[�F��|�c�������"REg�R��Q*�l�\��!5�i
��f~	���C���<sfK�B����F�tTS��1m��c�q�b��>m^�QM��ƽ�
H��6���FRWa��e����� �6`g����J!�s(o�c�����% {��a�c��B�Ͽ|r�۬}j65��wPTe����-��9����(J�f�IW�S�����"w<�,�#wͫ�q�)�7v��㷈����O�	�o}n��p�aG�saK�)�LL����B*>̍W�`�A#zuN�J�,�5G.�(��
� �J&j���Tl��a�J�z�������'Uss5�>���?��V�r�4�u��c�=3���o��|�|V���ǹ�΋����Yv�RVE_���ޢ�D��5W!��`���V�� ��*⛪�C�L�(G����/�m��tՎ�e�1d9V/uٯ_в�ގ�h0�.Lvn�5J��O��B�x��.#��󂻍��.�B�v@K��A���a?nB�����"����6>�=�hN�@�攎��9�,����8 �ր��J��� �$Jkn�P5���� 6�A��	+�C����A�v��j�_ѫCb��K <��m�_�@�I��+�aI%���I�����|���+I��&�w�����c��#lz��$r��l1�i�r,�E@��<Gh0��@��f�ko�k����)ј����	�� ��uE5��|�-�l9ꡮ,�`JR��R��/���	!%�����kjh���Ν5J8���S�6��q����+Oq�ѣߍ7 &��qR's�5����.��_9�wM��2a5�ZrW7�ކ��^O' �Sea��9{�̔gz�8��P�����T����'mR�(���Ms����g�$s?��������D��(��,>�w�"bh�d=�M���s�QZ���������Ϫ���f* mEcO֨D�ُub�n&�y ��E���
�^_���H^���z�?�ʽF�M$"�M� ~a��;�.۸�!����T�\[��M	�L�9��tx$���Y��ө�`A����~��C�ы�R�F\{�^g,��T/�1���e�ci�o�d�k�9d�d!� �-Xw%%�^�%��{�J!U	8�rp	:k!����2�=�ɩ]Y��V����b~_)h�T��UK�Y�%D+X
��A�R��du��Z��l��(-$��(�*Y/z\~���:���\�=˽��h��k�m%:U�����5F7k��r/��to�/�Nɬ�}���irl̝� M ��g��h1v����}h��I*���/q߼���9㒉M�דbzt�X8�5M�?�7~}��s�"EH���~�7���Ӗ*Wh^_���X���DB�"��&�HԪZ���ne��(���"g]�b�|<Qߔ,�1��
4� 	��kB@�(_VY�	0T
�.ԁK:�7\��oBl�C��W ������V���V�0iXO��GY�ll�'�_�a�4���V^v�I�D��5�k�X����S_JB�����m�D^�ߺJ�,���9Oz-�N��R�BNvW��tcm@�4��Y��!з=��o�Z����":���r�c��m}�c�	�I��Kg���c�?�c��`o���84%��#����e��	!p�a��U��4���ܪL�{=�|��� A��!i���0O��I7�)/$����XZi4�D	�����(�)� "��&1���t �����|9�w<��7�(���r�Ʃ�Ty�9�%�U3�?.O�PAIp���u��=�S�$5n�.9%y��$Rp�:bA�;\�+��Ӣ��l�n�;��D�`�<�ջ$.���VK�����p#�Zub���y8�R~��~>��C����A�S��b���35�i��I-L��Վ���J{@�n,�V�������������U� ����P�����/�8����@�Y:���|��66>�{������b��>wW��U��*w����7#���
%oT�!b7�X���S�G@�}�&6k��DU��-��5,T��;'�ڛ��T`FKp�z�5u���dMdlQ��R=��K>�c�ܢj�:<ponR�8ar�x&9*w�[� �9�'��`�P_��RQ3�<3�{d;*Y�O ������+�4�#>�$P��=����kNk3��t����K�3�d7R1��!-~Pㆃɩ1�S�8vrF@pOL>��&h;��q�������$���*��Bf&&�@�`�0~��׾�!eW?��*�6_�DC���\����-�d�]mP:��&X����gl�|Oz6�$n/\m2e�U8K+/&�uK�ĻJ�-��ގtj�j�l��P,w�W�]�E��kg����b������Y�g�ۻw�V��'*�t��qX6ZN��$]ѿD4,����s)<�k�en��P`�fI���5_����l��*t��A�xr|��0����<T�57�Fu㘘���w�=�gt~�]��@Gl
��DQ��O��F��G5�Db��tdNA����E��]A@_��Q��z6�Ǹ�"f�S6�ϩL�i$�o�F��`c�7�t�w��UU�'�{�����7r��KZ�:��P�\�.�Z}�}���%��E��_��)���(pHY����+k�GF3˺�&~0��$�x�W����"'��1YN��44�s�!�n�aOi�J��u%6��RK��v�|�$��u�i�B�E���Z��u:x�7��N���n'C��Pp~-�������n���ڣ���#�:�d�/�+���8Otͦ�:Rn�sr���D�f����	6e݄��5c�<��4�㙢E��|uF�����x���a؞�xMK��J���a�_�F��[=Z��"�̰���{�*��&�������h���ͫ�&�/���?��D��)'�Tm=��Iڇ A��ԗ�u}P�#���X5�;G��	r��qL�~β�ϭ�6��ޚN�<mL�#di��c\��e�ϸ{hy�"#���[�0��,��.Y�؉�O��E�;��1 �7Bv|�^C�u_���X�����U8D,���I���v/T���l��j�����]ϩ؂[A���.�$���,�{���Yfu{k�.�K|A��o��WB�Z�h2,I�iҗ���X+mZ&��
r��h��PO*��M�K��G��OԹ��`aG�ڬP�vG�:�ZK5qr�4NJ@���?+Pi؇��y��T���PA���U����B]	��o���GKgW�f��g]���8!�"���A�����AN3�� ^:��洕�+�h���n��_x��f��r��A���u*�[s�i���;F�����\޳2Ga={��}�~%�	{s�4̘MD�5�8w��C�JRL9?j��y�ea)W�#��3�C�O�?��]�AX��Gv��]k����<�;^c���I��Z�T�O/.w�_=k���Q=M"l��_�\��-p�_��3dH�N$^3�	�@~�7t-�jG!�#��ܽꇞ95���L�����.����a�߂}������C�3����4��uZ�2�
�߃�����ZQU�pVh8�q���S���A�d(��ĵHB?��� ���V��F�\C^ô�2P�3����N�tg�ʂ$����U�2�c"�H|�w�.<�?���n,�&��(Ɋ�4��Om�o,l�O���4��w��$��W���Q�ڌ/�0G�����u�?���;�1�ҟ˓t�o��A>�vk��~�G��Y�����%X��h��6}H�T v���;ߋ�,,١��r�Q]���v|<St�R� ?�o1Ab��\X��K�¨��Y�e�̓�كR ���R��j��-����<���CT�'%g�'PωHQɶ�>��l�-���X�����j'p�5��x����H�M�Q��ģ�\멁�V8��Oj�@�J�K�X�g�5U���+��D[u�&x�Fg�P�8�c��	���J͔k�pb��H���.o��M�&U�<۝\��*��x]�z��6[���@� �QN?ex���N�ղ� ��b�Qt[��,(~#<����i[�$�����@z��u	��
��;�_��bxQk}�=�M�M��ŧ��8v�֑�pu�D9%q0����an���~���#��C7v.�ѓu���u�=PzŜl,�о��a�NU�j��� ��C���Ś�̥��L읯׭֮Is�����H�b�^'���Q��5 ��������N��bm��m&>k��V,tF����/<��o�ڨ��î�@i���I?-	`�pD��,�>���I/Aj�R��A  �.O��Ձk���KkY�w�у?=+�8~<u� ��q�;*��Ke��B�O���2~#������Ɓ9-��z3˟��fʳ�j�az?�u2���t�RRzi����aX�eSN�Lև�B�\aFK��5�s���")y�{|�:ފK����RT�����j�d�>>f��2�l���*{ߐ�2�R�q���͕�)}y�> \���yH�����?���J�[w�x�ስp⢄0�]��C�$�]l�Ũ������
N��Qz��b�R��{�e�>ؘ��fpc�vi�����u��~!������HG��u�X��K�L��q5i�\�ئ�SJ�|�
�a�ۜ�\;�ϸ)�ϕ�?�ȹ�~�
����\�6m�K(��vCr:��R ��$c������/�����b����@hQ��$���2��%�D��H:�p������M$	W	:�,{ �����+����䠭�J�3��2���R?˙SQ����|��5���A����<�(�1põ��msF��#>�Ft��z���x�G�qa���'b�1���/��rf���m�����&�r��c����5�%�K E)p	a�ԈVM��i���#�<h��R�$��2�{y/�_�pg��48v�`���u���d͕�َ��Bݛ�D����js��7���X}�s�aL��n���������-�"fWxZt*��*]�I7���t�����:�����x(��%tIJ1#mc��l[���S��B�"�^��\�mAx	P�ƽ�ց�ԸdM98J҂�����Z�=W�tZ X�%ȣ#=�Z��\(Z�ԝ'�.#�-�F��{�r��� ����BϘpk�[[�:Xss���]P��,?���[;u��I"��� ���u�S�5�CF>�?H�8˲U�7Ӥ=�1@=U�^�ٔ�������[~^�lm$�%�)��%F�2�G�V`���(��P,i�m 5��8�:��G �i�'V*&�A2�U?���%�'��ӳ��3�@H��~?4�QzC+Q�O_�q�X���uq2H"������0��q�\��?yw�,�fd�+q&���j��q;��g/�N�ϿN�Ѕ�$,�Qw��D�8�J�<2�n�K�c���0�¾�9��e�����a��|�y=�LQ?fө��dMS��ԟ!#����Q�#����V�~Y)��K�m=�����]~�h�#� 0;�Y��9�͕��%�E<w������z�W��bM�L�Ht
j���y���2g�8%���U�[5(MU����1��/�1,6�D�C��&J�si���`�WE&J�J �d1���d��L���^���z:2����S��&� >���lb/.�8��Д���(5vg|�? �j�@R�̿C[z��IE��p�T�����{�ڣ:q��ֆ|V	��i��|D E�Q��4���u'5��>���_�����[����O���?ZrwU�����5%�iqE͸~N:f=+yvNL��r��F�]�`�é�6|��kj�^�":`�4��ZR�a�/R'��<!B���\��Z��m�MZ�c,�b/���[��?���K�:�����$�g���]Q�D��ű��[�R�K�&n�%*�F���E��� Q�^BȻOE��c��e�pb� %|�w<]��m�[�0��4�͸�l�;T��FcV9��a,/�v���}\�Kz�O�J�I ���B�@�(�6#<�+�I�f2[i��/����M��sQ�S�2JDŎ�n�� �5��Vo��ф�J�H�D���7��^Q���'����
�Rܠu6%5�/�\�Yb}V��F����/�XM�,刹l;n��PX�WE���d��}���l�ty>8r�\ ڋۡb��y\JrV9 N[ ����+lϢ����/eC>��|�3!������x�U �L��*D��� �S���U�����9���:,�gM������2��BK�����EP��^h���^�L��Au������e��x�~ê�E�a����*~�'�jhL��=��l�5G�����gI5S.�Zf5�s��U��R҅����z�&WC���a�עaԬ�f�����Yia �>��j:0G5N�3�婐���{`��n�y������a����K�?s�4BH�¬�\��l�8wn�	�%�7�0���`�8u+I��詷��{}껬)z�]�~!\��7�I��R(4�f�[��{�s�a���8
!`?��DU>|�8��g����x��$:�3��pVۯ������M����  \��?bm�K̮Wb������e��}@T�o��x�����Ӭ$:af���t�����8��x� Z�*f1��>�>u���'��w�;k:�P�|��>U��8���m�$}&�!�ފH$[��ye�Wxys�{�ȗ�N�Ռvv���ujT�vǈ�oMaP��7�`|NS?N[xw@x�����x��1Cd��k��cr������	�����2��?�}��y�I[E�,q�,ϵ6-�o-�e����?p�UZ�D�� 4�<d$��s,�C������Y�Z��	D~��,��7��7'�ꍕw�W̷��OQ�:���~g<�@p���Pt�X��l>ڬsrl,*/�S��C���}�b0�]��������'���?�����4��:�B5����U�W�LE���&y���CFUa@D���<�e��o4���b�V�\`�o��	��wIZp>����
��z������	����kC���>�vh�K�N^�^��	!�jFAg�&�D37�[E���R?o��Se�ǣ�gd�Ŀ��V���5�kni f�{z�oI��pz~��O;�RvF���b�Y3�p�mGAiܙ���ݽ�NM	��[��]	��SXr�LH��]�{XIx�k���b��T]eJ�	�௤�}�]��!�
����=~6:�%��]̮�"F�]x�!�y���A��gh����2�v�Q�$-@�� ��e�wG!=@�С����b]��DzZ�~&��fS#h�/'{F
b}hq�Z뼏�YZdZ-�!0ǭ�y����ߤ}X-�0u��r@%{,NЎ^ۉǪu���y�|�q��z�[ٗ�O>b;��s��QLP6�\hh�����U�Q��1}��ۆ��l���BIϦRfs��\�	;��7T�1��8���L4�f� �M]�oo}z�L���B��b�$h�q��L����O�S����iEt-k���T�a!�K%��:iNz��"���`A��Gm>a��1��������ņ9�ȵ �%�-�suë�v�oF�j�(����S��żwKU˄�\�D�46kĆC�����66�n[
I�pl����	\�6N|����eѽ�Z��$o,>N�m U7�\�p(Zf�XIƲ(�X �a��$��ĀeY;� _��^��|����y�#�&)�l$�1Z����È�b"&�M��竎�)��j�����X9J�YX�f<:�݌ML����w�4���s8�1��u5P��R��˙�?#��IWt�Yv�o}��;6C�[c��@y��IC�@/i��(Ԭ��q�4�q�-[�=#O1�G�R�X1�o|omu���g�쪦V��p�10�tR��ȇ�A�g��@�g�\�""�Ɨ<��0���P$�vm_Siz ?�O���@�����+y�r+F�Ĕ�j����9F�2��E���G�CFǇN|����A?�����~{���ֿͨ�
ơ�$\F�=�$݄D��+���k�S��9�W���]���'4� ���>��d�������R�7^�-E�uq]��^��������vm����V���W^2A�."��3�ls�v�z��%ࡪ�,����C�"+ϧf��;��:����#���D��R=F�+����������i���L�W�uBM&��+�s� �r��fCUb �49��WM�wp�N��P��7�3l�+9�� Uٿ9��~Zr>ju��f��Q�~,�6�'�m�#��_�B"ڟXf�����r����uw������HޓI�iQm����?�m֌�sgp�BАo�^���e+uW�N���]���cǑ���y*��0D�����LÍ>�7��C)F~�z� �ꮭ�������;V]�\U����Ցn/�u�R��o����`@|���$͸]�W��ĺHCxl��̙Ya>��ֳ��S�~�([|�v�L�$}m�)Bxh��1�8#_f]r�A0�`L[(��V�����p��1��M�Pb����i���	�V��[@[�f�]���KyP~�o{s6�jR���䃊G&�<G�,����}�6|�W����~
]"q��l�J��6�m�a��!b���A2qj��|���_��n�ّL\��8����Gln�8�a�/?ņy������{�z���Ʉ���J$�'%H��[�1N�|W�9%K*^ 7m
�_!��|�U�G��S�Mt���s�����	� ��?�H�`�-���
9ޕ`tu��>L���;c,z^�ϖ?I��s̛>�[��t�Fdp���k��쫶��#��˖H�x�^H4�����t�~��]c�����Xm�>9ELx���:o��i$x��[��Ԯ���Jږ.�w ��ՖU"�w���uթ��w(��9�5�z����n�n2��'ȿ��#��O��je���rH�e��@,^-zK��!}��������v�۞d:���Y�?H��*P��m�qM�C����}K԰�,p���v���C�nri[V����­� Z��ydu]Ń7ϵ �K"V�JbQv�އ�=���O���3��g�2����c�k
P�Ku�΍�{G{y��j4�A U畴����w��@MsX�B8�,�~M2��!>���&�V�|A���T<�Dyʗ�iܛ�V�s����RxU�y��p��h~�?c�Z[y��`��_�W���	�/S8��ձ̅���	5*f���u�����@8�8���0]2@ʇ�]5M	e*fi`�	�4He3���_	�T���}=�����6��V�p�"z�!�;�ظ�!�����,:E��A��cY�o����Z3���J�3�}�D�|��`�BR�f��j�	JR͛.3���{i�k���<����O<q�e���С�2ψ�4��Q�rd$�K<���6^W�[+t~!�n@\Bn�UB�$p��XQ1߿����{����%�����GS�/�B��)v���Jr(^ӺU���&��ޤOj�߶}�
H�^	}6}�x����%}ͭ{U�C�0w�y!�0*�(� �!4��c�Q��ⴏ@�����H���5�j��.>��H�v�%�R��0�zH7�,�zc�����Glu�-vym	<@�����=��%k�S�8�0�f�9���SY���q��TӇ����a��oPQ��3��߬��~԰�>���K=��]~"��&�w��nE+K�dkļ��&���R�kٲ�[<ԙ�6Tw�l�Y�|�~Zb���c�����:��r�{�������Q��v@:�g�������@%������,E�&�����jz��[�$e�F�/ƂyE��Q��[��y�4���;�!h�t.�K�EЊ7���:[G�2Y�;c��n5�0����41��p��bcn��~�D)���Jr��|�����
:R��|��t埉�� �%�Z��Z;�ݶ�֏�F~�=8"����A���:��oF��OV�`7�X�Fhh�B!�]n��P1�-�Iq�&�|[�h���>��R�]�@Z�UV��cs�Uxҷ^j2=��ڃr4�Ѯ�8c��'�ꎥO�M��VF~E��Q�/���O��qS�:(i�H� �o"�&Um+�gM}W�Qi���K��=ht���e�;z�QO��ô�v XJ`7����ݴ��4��=���>x�C_Uj��~Y��#�[��>�[T!M�ɶ�,E�sk�|�te� V:�$�Z�|p����%~Ǉ�/���s��A�K�N�2h�˿��Zk`P���٬�t7T5I|�旼���C�O�mx�F���c巩��x��L�3�D�N��SD3�BS�`��Q1�	����q�l�rT�V��f�&bR��Z+�|Οެ4�(`�(-Kծ��E�����%�.�V0�א��DW;�T���8�z�D
4U����(k�?�T7�:S����~��F�7Glk�@� g��
$:�v�U��	ʓ�=�T��LZ��Ә�A��g
�k��"��ל��]�#�^�P�����iKAnޢ2��X�[���QY)��EѶ���q":������O	���������fP٠��K�9/�Ry#�#b͉w	��j�J!!b?ɉ�8�w}c��B��n�a�a����R��ݛ	÷�P���_N9��E;L�r>��3�� jߞ�]H�ѣJ��?�a�>�V}�}KWЌ��$��?#��5�ӷ(�i/��*��,�_��ѵ�Ǟ����(z�g���蠔�q�i$��tR11��8Y��9i�nA~�J�n��G�8}(NͰ)�$�,ߢ`�.1�3���ڴ͇D#���ǖ���X^ܭ�%4ꮗLb�^v���ڄ��mRG���4��q!mU-�nϤ��:�O~���Р���gU�L=��"�����r�0�J>��g'	,���͑3�ߏv��J�?|����K���	?�`Wqs(ms�Բ;�;$|�j��aTx³��]:`>&��F�҆�/�(i��Ψ�����r�jmcj���qFwl��$��Y�Kn���n�E�d�0��_>���$�6��֖�Pqx���E��j��)R
)!�`��R�upU?�l��az�FN��/���6�H��6A���u9�
�kN��_l�ق8�zO�bT�}y�ߝ3@��� �ʶ�ka�
�T���كLD/����k�����m:�q=FTQu݆'�_��~DWv�p�H�{�ǣ����W�E�PH�7W(������ŵn� ����l�Cu��:
 �	p�EMa.��1-��d���y�H�I�Ń���^�/v~�c�?�D�tM��^5[����Pm��;�B�(V�F�^3ܬ�<@{�)��i��3�'t�+z��J��aT��� ��E�Yw���u�*W��%w����g� }��__��G���� o@Ou��JYsG�D��_+aa��*��
��4���77�7�%y�[b��dW1�������_/�y�{9�G��2�?y��.�ôj�U�l��]����Ȇ��&Tǔ������3k�<.���*���fx�޽��;GC���+C@�ͨD����H?� ��7$��7�9�F���~`���&_2,����m�� ��(�P�:9[��lj�.�bY�������D�������|�$6B
�s��t��2�t0��ڥt�[�|s��c�F=�|(�,�����d.���D������.+ŧ�^��V��ۮ
��_���G��&�!j}�G�=bJ~�G��ʔk(��T:�)C1�W�+\G!��oyն��/��4U���Z��w\[~!F�����j~c|Ù��gD~�	�H�ݔMm%���iUX�8�e�L(�%~�Ⰱ���ce �𹁲Xlb3�mg���p6�����C($��S��(A�R��?�sG^ui���%̺�O'x�6+��J�$�K8؊ߑH',c��Ĉ��є�/�+*�
��|?�U���j�1u����b��U#�9]g�����I�%����fσe<%�9�7��&#�-�n;^P	�	N��)U�����Ei�I<1���ėBr��I�(�"�k��JZU+���]׺�a�Ǥ*�׆��9����a[��I�z*PvA��W�O/�ͩ�fmt?n�`��x|gesS��!
���90���C�����b�R&�����tï![X�;��=Ɨw���n|��S�u����+FO�'�����E�A7��UV<~���k��%�pJ}�����j�ӕA�i�3��}��]��L�Mkc�PDb���� �qNy�^�q`�{JK��[l�����y��*\^�uk3:�܎��7�ɳ���i�҈��S������Pu�s��VS� ̶ݳ�h����,S�Emr�)�0�:�[�B�t�*8:xs����Gl���`����p�a8uӁ��)�6����#�'̔��W�X�b�b���a��dy/��s���Ƥ��=�#e؄8�#�IX��c�����QO���&�>V���wg@E��7�/�,��Q+���n�!�6�Vq]�Mu`r�=�-C����B0���o�XK��X�QR�s�����A�S��2I*.� �f;�O�Y��E����<��\�gՔ$��ڜ�_9f��e��|�Jf��D "��J���m�D5�V'�.�ç� L�N]v<4���⛖l��F8��D%rDjB즵ãڅ���oX��4�Q4���<D��z�s��PrD�Q���!nw(����}��BM��H���x�y�k�H㜥�KTg�Xo��~&VlcR�=^����J~���b�?�bۇ�[��:8�.�X�Yux���^.��a5���Mu�c� .м��_F�
1e /f�ohC�B�JC����uK�/��q���E�<O5���)WqB\{rH�uh��oJs|��ek幉-��ӎ$&SB��X��9�;�[����1��_ߛQ_�E�/~Ƌ������(ׅI���Z����l����E.vW\<d��p�}�<_���z�_���u��Cy?��!1̖��$֮#���7 ��@$��Ӡ"�_�K�w����ީX�Y�G��+���`�2�?�xڲF�D�M=;m���̌�v��Q��ֆ0GQ���z��ϝ"��@2�
���Ne+j/���c�F��MB���C�ɷ?
	��Ւ0b��4N�cХ���o�
�E�~l����bٰ-�������Xg���m%]P�w��rj�0���J�|g�/z�0gRd��S�o�\[�g�~π��`��2~?�y�$��*��xcv����o��|]���Y%K��f�f�i�N��
��!�?�����2r�؃���f4��eܤ�YPC�ʾYd�� �O�x����e9��BA\�)�u�x�"��')���K<�uM��l�����HZ̥~������m����z��YF9�U^�f�G_;��\�m�
Wl�ۖ���b}U��H?,�?���+���}�C�Fi�Fz��D@��n~��b�iXi�4��3gU��a�Z�}����`��1D�9��)�m0�X��z٫���Z�G��vk�}i�F|�X篇8�Y٪)�G �r!�� �rӌO	Ӗ�5bwȁ��z%���\]ס��
zS�j�T��G�V����Eo�-'�)~��4/���I�}���N�\�NCP�G��o�b�d�1���=!�iG	��n-P�q���o��;��я���[�8$VoV�\yU=�z�����C�e��>ˉ�^ۗf�'0�Ȝ��E��~���;��V^a�v��6�
�����N�E�oq,}�`oɏ���=�(�:�2�H�aĎ�P1gw�R�(Ӎa� ���G �F�Sd�EҾ=��0�;���Z�A]_^�!Z/���ġ����/Y�f�T"�.y-�Ux��9Ț9j�/��� C��ݻ���og;ro�-�֘�|Q��C���㰒>������.�`�]�~�­J#���5�i��Ҹ�n��i
	/(s�sH�g/S�{p�橁 j�U0�gQ�>�ڛ%7�b�-5y;ʮ桡z���|x�P�r������Ʀhn&��[$���S:wUQnV&a��*��
�%�ʝ*ҳg��Em�_U�Gs�i�d��8����W��8�\�Ǚ_RF��uvFŅϦ:�AQ����(3�!��N�I��hJt\3��j��EsX����˒%������b��m"k@���@(��8Ń�~�E�����º��xW4w�l��65]�j�2�RY��8�VHl�� ]�;W����_�Λ�^��3)��)x����QT �=f��r��3Љ�g�O���`.�W=��*��m�
�5�7��X����o�K�M��6���;lۛ���i �*R����y�u92}���Q��m��_��sǧ��pl����,vm�y�vF<�Y�D�Ԓ+��e b��g�~�u��ZY Ɋ9)E#���HX
'I���L(���=f��݁�5��J�Ln>���	�6��֧�b�̸՜��rr�%]�wͺ��n� ;��P
F�)����J]OZ�q�˘MD��c�Ӭ�mt��|ʪV��b"7q=��&����'0yM�Jr[?Q@����!
�9�MK�p��!'R�k�B�� 
o� a�x
�=�W�J������!k@��%�3��vbOӱ�D,�g�8��%ۃ%R^���i�V����]s��!�z�_�(�#Z��4L�>�V��N����I���=V�VR:o��8�]��s��L��l���v�]�[D:�V^�񩎭��{�S�z��V{j��[�D����aub��������Ci2�z��jX����j�d��{����P@ x]#|@)�EU�?uf��V���k��ݣ����V"5��%m�������e���SNE�Wă)��w{VXF�M�Gޠ �V�{z�H�ֲ���w1g"�������4?�F���ISP���A��D�9�R���G! S�P-��ۓ`��;(�o���x�$���j �ڢ�,y��@�aac3O�!���[$#`"p����r;O�ѰEv�'�ǲ̩����p~\j�*��F�D��)��^��÷؇f���[x����4j�Jd�A�jY
+�3x�ޑ�9�qYŵÄQ�+�7�3o�$��4qL�2DM[�N�� ����f�P�h*�D�փnu�ή^�,7-%�aajX����-p\����(���Y\gݑI��j������F,F_�ȱ.�ה��T��y����B�`匐���vKR�΅չ�
x��I׬2r��e0%�L�w���7Z̡س�b:�u��%��@���(]B��Hl��A�������cג[X0�3��2�o!�$�QP��X����7p��(�髈���_l��������V������
�C����z�쿦�JpQJ\4�����-�P���f�O8#B����?Ҩ񙊶yPK�)(ğV�!
�Q��ې%����]oc� N��\8�Ӊ�|�!Epw�8�z�/������h�c��V���I��F}�K�H�7�0��ٲ�x�����y� ����³��h%��:�����"����s���'x;���{Z�5��i���T�*K��)V&ԥ:���^+6�J^�
�
�q��I��B����/�����vEt��ê�r�?����cM\���q�����.*�EZ����)��z�:Q9;T#8-d�L��Ot.�5P�o�B���U�C��aJ��C��ϒ�m$?���AK�_��C#��24e���D$@��H0���L�n2Nv'r�~a���vt����v��a����[Ct_�fy)& �`^ٷ݌K�(fWM\��\���2�Ņq8ܯ$��C�2h�3�r?�qy-s9���'0b!��M7��Y�#�1 ��F������9_����D�fBb��H������1���Ða�FhM��	���:��em(	���R�t"}}b�ӏv&�'ݞ�^����*Ʃ��?m[��h��a���с"2�x����X���l�!e�-.Ӏ�3�� �"���;�c�È�]�XB^2�������=���$ �D�?&G L��ptJ	Y��w� ��:�(�#[� y�Ώ7�X�K����F'���$�M(�6nBMv���S�F;�6��èC�K|-C�&$�W!_p�Ύ!ק�[c~��(��[%�C��HXl��6�d�^W��)�ĕ4�m8&-�T'U�9 rT�|J[�t���5���=Mt�QN3����8��30#�GF5)GK��>x��#��}8BŦh*��Ŧ��g���d���C~�WBs'��Qo2��^A��̀J�&��
h'���w���4eOP�aAh���ٴ��%�bW������NƬ�]�x<��4�',���?�*oM��^YJ��!����:���(�>��dDxJk�Z�ă�[�[� ��������vf������I)5�f�0_G#�h{�t/X`Ot�K
2Q��,Z+APA�9���6d��K�yE�h:�õۘLc@�*����%鮵!��V||3��,����P*�ֳo%+�m:R7��J�����"��V=�Q�ϒ���ˤ���L�{��x�H·c�*|C�i��$�k|�s�aP��e���yiF���^I�������E�T����n��B��]%r>�l�\�5�:��
|��]��f%�1���j��i�y�� ��" �I������3��(8\�ԴЗc/��q`|3��8�$ɽ�
����a@X������@�e��w�,xY�-�f^� 霡�;o�0�l� hެ�
hʟ�6�8$L�%X#�����mf���ľ����<��*`���U���r�3X��|�n��m����Z�LAf�1���~)��X�6�nt�> Bt� <���_���J�K��Ѵ6�5��#���2�������U�K/��r=Bx蔂�8 B">C���OI������|f�=迼n -\���R�dU�?�8��%�g���
kBGgÜJ?YS��M"���D��k\#�>-��)���܃� *ʾ�����[vm�y��5���4g��k���w;�:��\̧Րux>S� ��Ʈ��������o����LZP9А��/��|�R�k�S����<���5>�`a)=�x��#�3F��Z�����F��=9˰�Xi��eƿ�	��Nݭ�Q��;A�D(�}5 &��7��aa�8�b�Q�~Ǉ� �e��$2;�O`��
+{4�
w8�����ǂ�(5[d*�H�P#ÆPm9j�'���4e������g}�������f��r�g���Wy0(�T��Rnȯ��T����O#��l�P`@`��:ϓ��iQd�^��[�?k�όڱn+[W��ЋEF��x��3c(t�i.^�(_�6����"��\�/�\"hD�:p	�zk6�Zkr���������3��0�%pW���i�`�'���T�D5&<y�JD��G�Z����i�2����#�uƐ{X w��-�@��_�t�ܒ�2��>J�9�1�dm�	���C���g*	G\�be^�McT��bN�����l�]<���m#q	�X��S�ݣ�T��E;�#���c���~�J�I�)_E���n�G3Jȹ��^���J�|O�ȗ���,�Y����$�r��$�¥̛���u�P������B�+���U�d�+wl���'0@%c/���YNq�����ј�`��Y�q�
�o�f���j��f��7��q�{�YQ�dΏ�v4E���c HA�<3����\h�W�@)�TH�ù�z*��[�f���N�ϴ�Sj�_��b?k�u����5_L��a�w�t]A��Y���/����M��Z`7�z�4����ٲ�م��(�mw���9��D
 ���@f��p�5�U3��P �	'���%�mڝlg�.)�y/g�+>��.�,�/8����ߜ^-u7�L&о3���R���&%
d����T��7E=˒����n�؃-�]��/��7w{�@�P���x�~vlƿA���2[A.�H��QYe�Z#�6ş� *�������� ��셭�Xx5P_Gk�X �ܔ��0��Ӻ��Y7���'�ue�&s��Վ�_�F�c ���zsc��dop�;���(0�p2��&n�&�͇��sO*���%�|�9* Չ66���i�AKWfU����ŀh.31����[idUF���0�kg_z uO�;N��M��X�{��;��O��0I5�!��o~9�ߞ��ʗ�^�KX%&~�����PV��;O1�iBVQ�j�����y�h�m{�Nǧ�D���{өG��Q�0��{��S����- {�Zn�;���\3��M��;��U�X�S�t�f˃��qj[��r��E���z?��EQ�ǜ�ձ K�8��@e���ĺ��L�эS���w��Lw�I��o����\�ҳI��-���mDz3�U���T� $��*�ʘ��H�q!a2Z>�_�o�������*C)������\�!
!]x�#ӳ���t�JUJT�%�Dd�2�!"Nn���߇��\8$�X����k�~�����W��&⢴x������(-YR�+,'�3�>~ۧ�1a�:�ņTbk:%{�e�K�c��UB󻂆F��D��:��DO����Q%�ES��=��#|�q�ݝ��*�4��:{A���rit�ɳ���v,=�]`M]Y���d�)}�\C'9 ��gx��W8��pU^j�초�HVJ���X�u
�3�����g��v�7�?�3B���K��K<_X�@��+y���?8����><�o�6�!�Ѕܲ��D���J̷]�jk� �9P��'�X�R� ��������i�@z��i)�"���%���^1Y-��Y��;Ϧl�,(��rF�����/��a�I���)/w���o^�ے�?�O����'�5�.�tn��2�m��]���r����Uv�~�A;Ns#�u)���)^��xn\ʪ�nܥ�wB��R)�J(�n3,�g�׈*.ԧ�'�3=�Py"C�`�'�e�*!Ӵ^߸�`�A�hvm���9�~;*��X��I����*ѩlU-p3��=|���yT�cGHTя�ZC"�ꧺa #��f� _x�O[�bF0��,�x�z�xw֨Z�3��n)�H7�Lv]�[���f������7������')�.;,O���ڐ~�c���F4|۹�+ṕ�R�C�T2|T~Q�@E��ϵ�]�>jf�V2��,x*&bIC���1���6_�G���]��Tb�C܅k���ħ�S����h�8��7ΰ���>��.�� �]��j)���p�|���p��}�]�V�6Y�Q/����;&�����)�zY��N�=<o�k��mv�����G�M_f&Z��R	�1L���}����H(������Wwp��f�~;?���1v<T�_��r�o �6��]�aH#����R;2#�Ye�ױ������� ��z���5z��|{��n>L��3w-ᅭ����@\?8V�Bd�3�[/��M�C�x�'�郾p�����J��ff"5R��FQ��؟������J3[��ʍ�2
�ʯ,p�6���{��RB?��D0��zh��d�7�,��*c���6*���iޮ��W�qHN;�Bv�@/f������r)ܮp�P��3��|U�����d<��TF�RE�C�u���y6�����=~4����B�)�����"��C�n�?�֜��E~����O���X����(ځ8�%��U�F�p��4&J�@W�xp�!�l�k���,/����LD�-��\ -YB	��g�f8��QE�5�}󧵑W��[3f�J:�m+(�(���s��/Vq�\�Eן/��.q�����K�2@�`+��ʌ��טn�q�<�lY��#2�/ƙ�r"���B�
!6` V�����`#5?���a��R�F���Gy1l=+�D�H��t�aCܤ�����zV�9���նl<>�n�s���:��X�l�D��A��*�F�M�D%3�~�~*m�S{��/��_qh���ItV�S�w��r�ǵ���s^�G���l��<I6.d�gw�V�C������m��f<B�r���v���<(���t�J��9���G�?g�p:%����{`b����+C�;�Lq(v�,�1����M,�aձ��y�8Y����'�˭>V��gL�:W>��9?� /m|��r��u2#8�&�u@f�_7㙂�6��V�q�ED���xNRoG�8Zz�ӝ��DF8
�A=C��%I���~�����öW�TKxY����̙�������A;>��3��?^��:��A���Ec�w�=�qko.�O���F�mo��շ���$r�P�n�ZY۱wY��*z/�>)��<�H~ߔ����@�u�nER&(Wf�x�o�Vc���+�m��h w�i������q��`�!�t�:iJZ~?�)6d����P`��쐱wo�ڛ~�<_���(����i�BM��o�����b��}$K&�zR��K�H:<{R)/��>&A'�6#g|�U��!�AvhwG�]l�^1��hǂ+��3�����M��i/��6��ՊE�ns;"�GH��cx	�qK#���FYpUl�,����c-���c��b�6�u�:��y�����x�?����`\Z�i���W��,B��<;bAA�	�l�����עAr9m=��[�nƻӹ�%sb���
����X�e��y�UQ�0z�F��#�"�C��҇ȏ�����S����A�Sp���6�0$����i3m9��	 ��q����V�_"�DQ�˰� ��T�:�T�hD��G��e���<�=����D-�j���x�Z�{���vc��vy����D��
W�����>������d�]����i?տ�+ޮ��G3��.�=%?���H=�^"�'���>�0�i�)Z�/2�D�2rA@'��2�[D��^�O�Hӡ��5���Z��\���`�����2�����9?e�y���cFH�&G���SB�p�W`�9�M���������öO�")T���h'��{�"�z�7f���)�-5�CF�0�h��W!uUB�9tPA�hU3Q�p����0l5X�H�̣~��e�;��*s��}�.��x�����Wg��57��C�ߒY/�%؂�� C)d<J��]./�'�����Kd��}���^�����W�ٍ�D��UI�4�<�3YVm
���K�}6nL@�P���G?b�w32�Qc�> <�6(��7��3S��t�|.a+ߡ�H��гS�*v|���q�l�%�C.������1�E'��e̦n�^�'�*�!��ń�ԃ��������Orc������	���=�@(ụ.Z�i��r@��k�}�^J����} Ҽ���>����w|�������������Q��2āt�X�6��y0ҏ����hڐ_�m�Y�aM!��`	]���g�Ï?b���0�;��#Gb�N4����o���ю�xY_s�ԍwo�s^��iI!����isp%xC�[pP'�6���c��1:PZ!Y�=wL���}�!��p�pD8���6�%e��IO�㮑_����z��ƅ5��s����E	��y��^=����!��vl*���7:�f��Y9��^��ƪ��p>_P/g'7=PR�sc��mtE!�l���61�t�{���d$�R��{�:Mb�o� ��U\�3�-�9�q#��tf[�kNm[�,��`q&��7���XU�D�Vg~��`��VnN\�i�88uDs��ʈ��ͮ>h՛$��4�M������И ��WAlzh��'��W�2p���7L'�x3gjI��J�d�����گ����7�*.�59�o/�5�ֶt�j`ˡy:�h��*�6W��rQ��kB2p79K�
�Rp'��L�>spt�R�2'��������D���f�R������3�q�v���_���r@W<��C���M� E�q�*���� )K/h'�Z!�Օ�I%��̿��¸��I����%Y%��%#,rL�N � C���!f�~�ef�Eb�M��@55,�y&��T$[�K�����j��]�4��Ef�DUƱXRh|i�Ӳ����R�6�x:�4�:��kDZ�١�޼_�\�̦�T�����'t#���̍�}�J�N�Q�V 4M� ��\�I��J�'��l���Y�C�t�Ձ����R��޷��
=|c0���=�1+M���rB����Rl���M�5gݿ&@��w�Yf��P��(_���*�5Y�����g�M��oM��5�pr+�}H��;M��H�*�T�8�ă���e[r��)iɞ�H�x�^���DjG����w͂_��j�����a�
2���C]��U�>�������sҭ ���ѱ0���ח��{���H���X8��Yz
��2����%n�?TEN�V��i|�^��������k���xZ�e�!W��(�Y��B�S57)u�I�y\C��ƪPD�m������j�p��L�1�ճ�S ���?�����rK 0`uO9�-u��Ӌ�f&)7�,�PoX���
��1�z�xQ
���7Olk�O2���(���E�KZ$�u�pr�pP&�莯8��G"YI����L�}y/I ��`�X�C�w!n��稫�ڐ��[�B�>7j������R/�<���eV��&�DUc �,��i��?ro����O�쬣O�����)�S�q�Q�Okf��G�W?�l�M^�&�Sx�d�-�yA�C'.T��C�:D�e	U�������c�GSđC�Y	6�ItMQAP0keI����$!b���g�h-�2�H����y����^�p�mQ��t��>տ+@n��/Ьj���*֕gP���m���}�&-W��j�{e�O�:%ǲ��n��N��Mw�H�[��j�	A���	'�w�i�!���m��_j���}w�m������[OR��.�O��n�mo\
N��pҖ�4�Iϣ_B��%9��>���4�k���vk�)0��,@,,a�n�(6��ʾA�ლ���K�u�� ,M�[8���k�2i�P;)8��z�q��*���b�M@H�F�ni��?�e�q�YO���e˞"�2�-�8�_��~jX���~L�(�iGB4�t�|�E?>�$<:���5����4�ь��	��$�(�����2Nb��,	H�0��	�Z��K*��`׏uau)���5x{�.;�F�>�7Қ1�?����B��^�p��тƗz� �h݄P*.A�8�?Y�^�PM��f9��̮*�������fl}�'��n�0��NW��1QAgf���3n�mq����ׯgЕ\��2q�6�p�)�,I?\�~Y)�z�w8�m2�Z�9��a������~yfDT�#�����"�T>>��d�Z�E�ZI�-�'>�:�g~n���ƕ^�{֪Ɉ���i&��If�uF�'�G��r�����(����Ʒ���1����8��H���O��c�`�D]q�[1�Ϣ��sQL�Xְ�����<�~�V�v5���G�gh>"y��oF.�P���g���v�9�$������<1Qܻ@su�Θ����
Qsm�Mԍ4�%�UW��9+����8I�����M��s?�ZO���=�!4�/��h9=�[�Dp� Ϲ醀�S�(��]/���_J�>�뎧L�;�kɇ�p_�c���@4�u�P�8�g罀�� wZ������{5��9����(I�9��V���ƗS	������>��ޓ+v{z��D1j���uɏ�\]����'�]�r�J��V*'�_�0�$:����n������}������\�;M"�l�M��G�C��`tk�&H��9�ҋ����T�/!�_M�C:�5p3l'�����{�� C�ͱ�V���f��+c�H�:��q翌��<;s՘��&�����4�ee��_��b��Auq�s��� LV�N�����)fSi��
Y+!���W	`��6;bPO��� D�_��3aj�׍��B��R�N��Td�����5����	�o�?#u�P���U�����m��O/D��t��_?��^]���t��t#\�Jt�$�Q�c�������w��{��CD��u�왥,z���ʠ��g�g��e�����F]�*�Z�= 璒��~6Owh����Vl�LO�ٺ-ʻ��,5��b�ˉ#AQ��31>^#�ۏ�W"Ϋ�
�)�DW|4����N���R�&���뻱O�|	�L��EU�3�\�ᗀ�q�?�>��9~ݕ<�>E��ÒNM0#����g�3^��2�sM�G� ��tt�
�\���%��ܹd݇<�m����Wa4�˼d^Tp����I�J��8�R�LMB�ޜd�R9��Y���&C�&���p��J���RDR�2�H�t�u#��Y���{N��P̠��3\[�%(?�Y��5��Z��хܞaW4>3��<;-���\�#`n���b��P��iˠ�i��9TU�%j!?1<[��BϨ$�͛��{(-��T��vU!ٜ>�����`��cO�C��{��+�k�E��!������1������K�wD��=�^q0>�K�Go �#U���a蛭����(Ơ%b��'��J��\k}6�dy��֯�L��֦�e��nӗ���fܛ��·���P�cf�t�5	Ok�&x�x�nk�\�����{%�r��˺P=����bT%M�V�[/���}j��K}H��߱��փ����ƷPQ�T(H�O}-ZS�ӡ�F���Ia���}D�T�F�,��q'��m�A�����	]�U ����J`����3G��;ƶ�3�m6I�Shqzx��2d�Uc������b1<�����et&r�X�\%4��@i�F�!��N�Wy�x4ġ-�ű���:��~՞_vߩ�-|v Q�C�8Љߖ�T�:4�<������ǂ�=e���TJ�&i͌8iRT�ď;3��ԗ���8�/(8<���)�e揮�t<>�F��]����;�Aܽ��({CU#V��7���(`ȅ/F�ʋ)Z�s��4�/�v*N�L�B��o'�ߘ�C�}�]�]��Hx�S(C��V�g�x�TwY�.�oi7��=�"Z�����o�~;-��=�[�y�9�����8O��3 J�2�'����ߕ���,��DKva)Ы~k����n���A�Ȫ�ڿo��T��������������(!��E/#	�|T��m11S�@�3��]�ݰ5?�HCP����u��V��4���|�~�J;�j�&7���8���[�^���ܸ+��-Q�,�(+O��Jգ�/Yh奎��p�8X��M`KC����[��V,�'�]�٥�{!�B2��j��2�:,�>�*�E��}h�U0��O`����ҳ]���4�������)T���_3�FKqt�X�F�3i*o2�㺕��ψ�WL�J�X(�p&�������m�1�?CLr?N���cNI�?Rf�&[Th}=�|��:h����y������jc�S:A���SS7]C٪�`�]3�8~[h�N~I��I{rJ�a�	�����3���>z�Z+�j8�u��S[���8Q5�j  �ř��\<D��wW�U���k������c*9�|_;�J�����3V��D84
Y�^���K�-�ݼ�o�߅x��="�
��|�C�t����J8�T�ޟ�D�}d����bȊ��s<B��C���E�[|���=����YZ]V\ק �f�M�䙁qM��.�А�.�ޔ����V�c�0������ѣ���V�qRH��`��rnm5�����+&�	��7��Q�ȉ�����5�j��Bf|�'߸o$A�P2��9dݏ+�Z�o��������@�0�?N?���9]��@s��Uۯ	���J۶FR�IWQ��G���wW,%4�M�^��Y�Ul��.΃Y��[.�m+�9�z���h�3C�1��a���V���IQ:�mW�U��w�UVTE�=���Yp-�Uj0'���=C��u��;:��;��y>����p�T��x'����I8��
Q��p�M��91�s��"��&.r�j�͠Ɩ�S��\2�~� ؊O�[5S�?H��Sul��,cvZ5�O}z��� 5�#�[w���N��z+�[�*LfK-���N	 b���xʳ>�$��}Ϸ���7�
G�歈<QW.����;�
+�K6O'a��"�](yH%b ��4��0�	��v�9I�핎6��]/��2J*]�z���L=�H�CQG����m�]�+2����HN��Ż�5f-��D2�F�ׅ����7����r�Y�u�S6Ѫ��:��S�J��{�MI�����T��y��b�p�l"@~�`�58�s�@�7;'m$q�y�F�a����NkHaf�i`A��i$r^�?�������d�y�0�$I��������@t.�e��eԀ�{i��I��(/RaT��o��`c�$J�r`����>��ʟ[��j�'���Ư`S�e%���l~��|G@�}�^�3r>������BB�=�U�ʛ��
�	*��7l!3��t �- U��z|t�b[�G,�A�M�
�i7�qdFvg)g2Fu����>s^܇�+0��|C5GlG��{%�.
�@c���۷x���2�'�Pn���^F@<xc�$e�����!g-��3QOxj��)OzMW����n5���
2��ޑ�%5T����k�ʷ�Y�h��K/��Ij�� ��o'�0d�.G���:�PrpC1fa�5�_x.�$�E���x%�;�BGZ�
�כ�����p�|I����IK_'����[oT�}��Y"{�?�C-�|�P�]�&��%�J=R$H��E�V����H �d8��M��+>T��Tډ�qt\t��@��g�X6Q����KRٱY�9(�zau��8z����:zW�oӝr���4L�n�a��
V^4褄�@��JVzK�X�xt���vl@RxE�`�w��s/i���븽��������XF5UG9�Nп�o3*��G�ī�-d�f��ElX��,*�⓫�hܟ�G�;UK\5���/�_/d4�h�rX*E-=�+)O�:6�9�l�p ����ҍ$�Q���v�Gӥh����Ogz���e��K��r��ǃ8�0�ߏ5ЧK�oX$�}~O��ae��
kW�",(Cl��Y�>�	�㫍{��<��~s1r!z��b�� A[�Y�AG���=����TGh�܌���[���@�Ԙ[jW��h��=Š'��W&���ziB��we���+M��5G��ٴ=��������拢6��d�3U�lP�����^E����������}Ii��t�e�,���q �u��lS�ڱ;���l4���� �Ǝo0��-��I�����05��`n +03��#���_�~ɡ�#ʇx�|ٌ�@G��y?t����R$#*���}vwr���[�b���P�V7��{#<��Aj|��hC�	�@E����eZ�-%�g��8���s�J'3��%��e
��R40/ͳ�z3�tm,�)�1�`��8����ڤ�<�_�kV`ͭ��	RM��X4�Et,3W����ԊYK�\ӉM��;ڍ������Od��hdOi_*Y17"&B�����T7�?aS'!����=��5O����[�B���dGD⭀����»�X��~e��Y�:OeY�k&R3᯽gA�?#\�zQT [�Q�/��º߶��g7SǯF�Tn�7wtR/���P���b��� a����,�E%��o�傐���aL�	�2�>Œ���!����� qs<�*�yU���`F�vWHM"|h�e��B�������I����07�q!�[��a,�r4��f��8�?d^Yf���-���:��:�1t����^A �ş�P���������hl_��|{,m��,Y|<��,�Ɨ��7V���<p$<����l����ϲ��������)�����%��ʌ��>W9̲}m��V\ܬ��,�Ki7x�F�0#��Mk��&�XY~�Ң3�ɥ�����D�L���H�e}�x~�����e�S�(�[*4���'��C�����.!����H��W�Tq)J���Y�(�D�{OԶ��s��{4��d�Jk�$|���0; \��������p�
3�W -�̪`�rD�<R��A;���D�eY�̰�J���;�X!��"�b���jOd@,���d���	A�4	Sg���0u��#:�($�BQ��<I1�����h�;��j�hgK왐�m'�[��T�vjtq.��aU�QH�H���������ͤ�͖|"��mH̝� P�aYw�]/���*�4$�Fڴ��yUk�<�{XT�����O��Xr`�Ŏl�-���3���p�է�d�da{*F'*���:]��w?�35��3%�Okg�}��d�'� �?�Q�;8��y���
��4d?�ڴ�;��vp?���3�x�=��Hg���֗��A�!2����q���Qp)W����&t���1��< �G��O L>���p([�����?p�A�A/v'w��`>;��i�dL�����4��h):'�u8�<T�ߤ4BI�t}��l��(��c�S�����;b5�A)�|(6ܠC^x
Ӗ�r8U˅�]F�-,�jd	�d������=P�/�q�aW��!�u^k���{�w�̺����2ǚ+x:���ٍ��5���	����d�sY�J\Y��6�����V
[ܤ��*@W����$�/�����=~��ܰgRa0;vK$Y�y���Q����O:po��6-{O|J��`�t�҄�[��Z��@|�;1H��R�l/�v@�ڌ���p��n{�y���P&_=� k�?дMֆ�=�	Q3�u�B&���M{�V��!h��۟����B����S9`� ���O$r�+P?��)}m *&B)�y���R?v�"�k�}��3i\s����}��^E�]�B�����,b�Ӽ�ν�P�aa*Q�t.���_�Ou�<��eT�@|5�P�Nrau�u�����ؾ4_����"l{�e�\�N\0���%��-0��]]"z|����^HxH'g�_�T@{nO��?t��J��:W&;Ik�V[�^��� �ƶ��E�d�#��U���+ja�!W������̕���?$rx��) ��((���Ǳ^�	M�����x{)�`Wz��\L���h���俈&(�0{�%_�"�l���4_�5��I׳��8�J �I��إ'�L�ZeǢ�W=i8�j��x�lR���E�A�m�^�r�S�*�c�՛b�j�\��_ۂ2+#w{�Q����dX�:�SJ���s�=����bbe�"��C���\�FUC�z�P4��/ ��V%�Dƴ:I���O�q�{��v�p`OI���X#�)rG����4��2z(���^�6��ς���s����X���.�λ�l�A����!�9�|�������Cc�Y�+:S�C+ĎɎ�݉�q�H��D��oR�6��()�*�:M{:���@�B�_o�$'p�N,�uj�:@������"��G�����Y-8Uzb�����$���l�)��j�j�ac�dǠ���G��}P�����o^e�
�_���9����#بk֝�h��M�L��O��r�c�q��a��9���Q �y��<�����VB��OĞ�x�J�z�:�$]R7�\�Ǐ:���޿ ��e���p�ؿ	��5���F��f�/�(�'��d-������U���YKA�!3�-�8�(2�W�p�Y
䀔����Gp��>I��M1�<R���� @�l�������G<W���9���uT��������r���/�o-6�Ԭb��!䡺*�@�Ё�.�	({,����_>�&f��i6�߷W׋�y��y �4�U��k9� �bx,χS*`X���ܾ�OCrឃ�"�O	 T��WN���|?�q5���k8R���9t��������k��#�S�NY;jT ���V*Ds�VN&m0u���j�*A�ŉe�X�𗝻�A$��PW��)�y:D��#�����������h�K�4u�9W�膊��/K�[�m/~��ȥn���(�SZ��*~��y�z�`L.����]�\�{\���?�ؑ&!�N�^�ĉ���J�#�Le�z E>ͯi�Ξ���5�^���#��ekyT�X3Ʈx&14>���/c�[r�!�f�X�m��:e�$)�����B�9/�F��*d�RW]B�_��b,8��bF�e����ĉy�� P��[�kt���kz��̻�P%������*��?z��
iq�*{I%nÖ�NmUo�� H��!Ç����4������ږ26�iC����U.�5�cqZ����a�$u-7��.�^�/���7��K�/T"���; ��v��+�� V4�͕ҒU�W-�oO��n�Z�p]U��Y��rKHv��&�IU����S=Ԯ.��х���*H��	�Z�+��a&j
��4۽�]��Ն�y ���58��5�K���L��R�?�U{hC(B;�̛����`	�N<>OJ�P����mc�'�L��:K��2�/���4��嫅�疬����ϹL�l|��J��/�h5��G��#�՛���%ju�ۈQ{ۨ���"m@���0��p��h�Ԓ� �3��� 	�p�N��I9���9��A��Ah�2B3��݌Ǔr�_M�	�D����ଌm�dc��P1z��hL�P
��>Y�_����b���p��^�$Q%ѩ<(&�힋��r�"@n��O��ƴ]���_]�WO������N���>��K���k�^>�S�ҿ8|"�)'�Ƨ����K��K�/"��A����]ٍD������-��)�������CT�u`���\]�]�9\`�p���ɭ^�摸��F�U3A?�����d�������z�v� �͎l&.���/��㾘��-ZΥ�?9q>1�o�Q9�)�g���S���4F�ښ��J��+�7NĎ�dج�\}N��)����G�J>_��ئ��y<��)����d�ww*Ʒ��a��gM���z�s�:��EC���<�rԫ�\/�e��MJ\	��P��;�g�H�H�c�U/�)��;o�t}%���Ԛ��ނ�Ψ���S��z��pWomz�}�1Z��=l~r8�=h�۳����}��#G�G9���B�s�l���oZ6�2Hy�~
�������^`o�G�ǛR��T��;�W^?�Bc�2�%[1������O�}!Y3S�����
Rp"��+>��-��	������]q�\��C����N�pJ�i���Ǚ{��|�( j����/k���]8 �Ն�i��;}��S�0��Cx �H�C p�)P>�]�M�-�cW+@�d���l�uV�xI[\�gK���g���^�Iuxa �m���_2e�.;�/q���}9�L�ÿ��T*E���<^�X�X4�|�6�T��1��i�8OL�d����P8K���]��l����]Ms3�O���;Q�~Ƞ	Q���	$a@g��/��X
��ɪ��uZGaߙ�O�XKn8����틉�]�S��qD�f
2{d+�߄z��)acv��T�����n}�}鍢E"���`&P��24TfS�2h�.��M�W��/�N
�N)�S�6�_ՇyTMN��*6h��)�ޥ\�(&��
y.@����k7D���F�"RLAh�N�ڰ�5�&|�&��/Gi�����
�)�f������ϥ<�?/�l%�}������/���C���ܡT��r�:d���t�B7�|	q�ˢֵA��[�'��\�Q��w(��ە�f}�7��LJ���U� /�����n�IC'��x9�ޤ��	��Hv�O��� z+2��%��و�J�tlɝ,~4�&�h�"RL�J�7�.ّck�� ��K�7$ձ�"pzq3;\ժ��tI�7Ûu���6���i�S�X
�e�KÆ�"���p鳅(J����n+���V<f�&wdTT�c��4�["�<���Y7��ԭK�N����a��Zo�$�����X�
-���\���9�Et|j�_].�.O4��c���k�����I<�`5t(TP�+�8O��j]��W�3��=����Mݘ$�������R8b��i��[S�@D|*;Dbً*V\33�&`��fs�Yq~�s�=���b�!��ڊDi\J?���S�g���s�}��NX���*��cW��Yb��]��7_>R�5Y%QÙ��<.�<��$�K&f�$8CB隠�Ó�D8���+un&Se��5溷|�7%}����Rq�-uرl�_��Ď�L29o�LQ�#�[�9WLGBZ������^/ͱ�\���:0Qӓ'e�N�4��$��Xy�p��9��\�z�攚ni���<Ҋ�b����x���=վ,p�|�O�NM}Vh�$��l�\b�
σN �-T�#�o�jn��yYT��Z8��'���vM���Q8�� ���'��C�` #ȃ��2nQ����eD���S;כ��yU5CՍ<%�N�#-|��nE\pmBfK�kc��͞�n �ѯ���k���൹&V�<`OD%kPk���{QYB�-�1��h�E_�'��F�K�b���s��٤9�x��֍�ݚ:��"��4o>��]�UrD�{σ�
�Z�� ѶW���K<h���\/*̧������U�l��|u�:$��;c�,�<��Du�ޮ"��W���f��d"����sҀ�$F%|��m�u|�N���Lw )~�]�:ٔg�
ی^�$S�����R��Ͱ�� ��V*Z�/`Ei�fFn�oDAf=./Hs�H�(ǉ��}$�0���o�ԥ�U!4{�*��d�F�[�HO��1݄�g��q�y��Ju��b��H���U"sR[��]�� z��3mTL��V�8ݿ�)��Q7QԮ�bh��x��,�'���Gmf��>�H��\ K:��;��^�zk2�GJ)�In�V;�Q�'�L��!t�e²r� ��??������s����1Ik�쑯*�g3��6,B������X2�G�pE:���˓��`�Q0|$z?m�]I�6�eL�3�v�V�����O����G���#j��yoC�k$6����a¬�@������yDv\{u�V5?\" ɗݢ��:Z2|�w�1�r6�ܔ�����a�䑥��6�6�涙J[
\����D��cR�3z��^�������$W0�dڄ�i|��lL�2+eӥ��r�
D�3�\�epz����?�������Bp2n��ڈ�y�b����\��2�ǹ�]�G���A_9�/�!1~����A[�⾊�ѫ�J	�=B	6��uw�����HrKh�|:~og�����zf,�Sטu��aB�C���E��� Gfw�F։i��Υ�s0�a�S	'�O�ͪX�m\��k>�u\[7�U�x	:�K-ɟ��ҁ�����Oՙ�@�V"��" �?���˥��Fj6�Ù���F7�?H�%Y��Yh�$DkS��=H��w��S���la��'V-[$9��j�K��u�sr�GTq���~������h��8��8RO�����I@�#YCX�a�'�m��wO(�6�<�9���n���j(��;u��.w�p�@��/N az��m��lC=�ʙ2'�4�݊
Ѭ�����2I��|W;2��B�#ʃh����֋�#�iν%@�7��U'�+�$Ҧl�?�莓͖�j7������Gw(�U�`x��vEg�#���m��uU��2��Rb��s`&��wo�k��D�E0;o�����[�Nd@��Ў�+�冮+xR���0.�z�Cd_�m���)Rf��p�Q��d˨2]ڋ^2\��['�y�G�5Yl ���3����
3�f�~x�<Fw�D�Nvm�0�%%���e�dE��������4�6�T].��+�(�{�[Rv��j�	8וv9�����!&Iۉ�����nmt�>�-�`k
��T$$��g@[v�W���pD�(�&J���-*�PMP��E�B\�7���W��txS�pE7!��`�+��[��_�Z�at�F�"[dt�N��n�T�}f�R����	a����3���e֨��n����Y�����8�7���*в��Q�B����So'��E��ܒ9	n�ذI8����M����6���6$�gI�p������^�ϖ��=����r�?C�ZA$'��G�"�rY�rf����r����ݥ�j�O�t���x��ǀ`e[�t�� 1��m��(��Zdxz+��м�i/���[YT�Ӊ:�)�2�cV\�-��$���Wl�Q����KTӏ딁��I�5��R������#�S1CPƀOfT@�m�!����(����XД�*�B�c}�>����GuC�κQo��P)XB�ѫn��r�I	?E�9���2U�'H���$��[I��(�}'�b�-fi��)�i������Yx(�u���Z�v6�g=m���Wv�����$n8�����K���b�������[�(�[��y&b��h��6��j�Z��3��*�eE#��K;�#)�7���2�[����s W���OF��Y�,�������ɑ�-B���$�[�L�{�M�n�)�H�Ճ=�|����ztԼŚ_��_O"�>l,��;�8w�Z�O������4�z���~�޴�Ug�t��X1�t��_��l6�@qHE�-�h���D���V]U G� C����%D�Q2L6�M#�`�B;��n�����Ƒ�X���%�zz
�rʇ�m�P�6�e8�MP�B�umP�G��T"�/�s���\S�]
���<�K;+��n���ݡ<����6�|.�wYQ��bu�,3/F޼`˲X�����l&{m-��8M��걷e!�����H��ِ�r���84$��6��H/^����Gჹ�� b�K�M^�P���!��b*L�{�x�m���m��6��ɮs�-��#ƙx�Y,XP޽3p���S���ڀ�(VH�H�;�	=��f53�d�봧s|W��NtoZ��Q��_�KJ걺e'K��173*u1e�0Z��Vm�n)j�Fx#�V`����e n�`*�{�ۛ4Q����2v]:h��J���(:�m-R��D��+ĥ)��7I�͜$X��.Q��.��3\M�[(��]'����ִ�Y?J�T������jU�5m��y+F[%��c�K	~�3}�{M䞓"��\W�>+:�齪�?��5Cg����� �NO�.�3���<�� k	Wǯ
Lr�4Eq��<D���X���ZT�b��ZȥvS���
�hf��U�?L(�z��7���i�{G�sk%s<�x�ݿŎ�J/&/X�b���*�*�����Ό+N�z��VG�b�Z�!˘j��1�<4�11�HT��ܰ])��&k����?�A����ZVz,�<�����̆;��p|2>\�H�S3��/9����I<C��;���R���}� �0��ߌW\�4��q�p����H��_z�7�2v�_n��½K�� ?to�F�ÒEҡ���o4&�҈����c�N�Z���qn�3�]��]P	����a'r�Cpd��.�)�{�{��?�4�� xF^��Z7#�'h��w��g�󌓒f�s�W_/����g�k`�'>�ee����j�A���#���O��<v|���o�ܤ~ݖ�`�ՄxCT)�`�m�;r4r��������E ��������o��GQFt��xi��_�׎�T�j��5���_����}�V���������@��G���m��7͠�K���=�t�o��j�7޵�&R��B&��Z_��Z�9M�'���[2S��s�^qIn�?��H�/�/sӦ���$,@Ԁ7å�~}7��X���j�aJ����H�XV ��=c�1]����m�`0~�
�j�/�b��
Ѳcc���7�P#7����<�!3}��5��۾�j4��Vx�[�J4������\��ڃ�W���/��
l�Jg;X��a��w�������{H�~����xw�O��粷M��VP���X��9cL2!wCS9�o`�5�Y�T��N�����I�ׂ.1�i���S"�9�g�MEH�ʆ!�d/H{a%����o�!"�
��d�;� �����
�"I[Ep��n+�W�킃�hk��؀
se9UF!v��va���E�~�_g�W_}]e�N]l�����V&P17�V�խ�D�F�C@�j��S��q/p!�;��#K���������4G��i�H#��ߟT旞
5��;���!��O�������M�(��S*�e���hq���#����������l_3.q
���~4�=Β���;�27B�a�h=6��yso�H�2�o�l�,��u%�ۻGB��\��N�_�'����R���T�G�E⧣���~*�-��3�F,t�8�m#�ή{�8*��	�uz�:`�^�#dJ�"F� d,�*m��X�"r��]��Ug^8T'���M�5J�)@zOdC����a�~��yd����Q��Vn�ϼ�;�'fv�Zw�mf�q��l�}w?`�d�FNKY� ���(��ק�j�Y�����IwJup����uMl�NDt�M�D/��q�؄:f�_�h�(~�s��!LS�Ɍ3����Iޓ�Ha
��>ihH��[���I���K]Fu ���!�d�J�_Q8��r���%�o6�������?��Q:jKᔷuY��*)�J����.�Цj)�I�!uŕ"12�ٝnZ�2����Ē��p	���]^h����*֬(/������,�0׎�&������aJ�����0��XshO��7w?�tHJ�nw��f��8H�}N�H�G㐈,f$����NO��?���"ȹ4~�/Y?�|ێ�jl�M'�@�+����Zu)4��Pk�4}���_ܭa�����OSv<mE#8�-H��l������B2�+T/)L�+Mw[C?�HI,��P���� <iz!�g���kX|VSJ�_$mh�����]��vU��h~w�ٳ<�/Rx�9n�.�'sYOU?� t;�8\���-����q�c�Z�(���ϵXH���/��I�ݛ��Q����8����N�abc��Ck���եZ��"X=y��K
n����n5���͜[�1��MjI�U����{v��^����1M#�Q���g�����9�j��~ٟQD��:���R�5j!@6S��Jds.�c�"�ɪ��v�s0�[��פ��/��6 ���W��Ż�HW���bO9W�ʟ:7#������#��5�b�Ռ�J�K��1�^h�H-1;0�
۠²]E�1�x|T�X7��urN�B������Ȝ��u��B~�s��e��_˔Սi|N���N�� Ҳu�&]�H|t� �G*�$ջ���)1CY�+�M	\ �7����)y�%���(ەJc�QE���jYL�1r���@v����S/A�ī�bm^�5��H�(,�0�/r1�$�?'�$$*�$��dk�mc��mSǾ.�ٶ��Y�me=��8H�)�
݂b��"9��q���M��7���"��������5�TcR��8�mw�&k���tp똜�X�?�������<;ռ8R�P���EҬ�YJ���Z��S�����RYd�7&J%��Y>y=��?��f-��\�~�Z�Y*#LXvխ❗ďp�H8+�tX����y����)T���i�N_�S����NpdyW��@ѷe�N6 ;�.�`c5���(U=1�"�))T�c$���rkP_�h b�c���s�ODZ��B��]z_h�\R?l�^:��]�:%�KV�`}

L�5��FE�o'��s3R��w�T����Oq�(�������WR#r�x��p�����F�V�2�j��//W�:�����+kl�(�/�L���f
��5�;��s��B��T�7�}o�~�Eug�s`��0l��@/҄W��l}�w�ځ8XD�Ζ$Q(��TC�by� �a2�M��f.��k�<�� ��r�]��T��r��Y���h#�m������M�f���!�d�n�!��B��R���n�-�<S|phg������G���# �:�M� x!TMR(�`�ѿa��������	�kE��m��|F"��ε����Z <�V��x��yG��k�)(6a�h�VD4�JHg�¬-�z�K"�h���9q>L��O|�?tb�2"f�h4���E2�:���Ży}��e�78q}Q4���(O�����k%�7���OˎԼ�@�=�x'A�4�H>�/�C�Z|AA�6u������!oM͠BQ)������ �T>�����΃�Ynn"��R$��29XK�yE�[Sf��|�e��'<d�sَj&}�ÿoK��������/�j�}u���^@I��w����t��RXk˪}n\�5�N�X��M���o"�%��B�c�G�S6�櫮�� �5�2���b��t����/"s���>,�%���Ry�-���f.�Pk�5�~���X�G�+(ɇ��Y['Q��'�"K�\ �����ݳE%�U��K״v�N&u�"� ��],�T��c��oo�s�]h�o1[�BCf�)�>TP�V��-z�lx�a&yV>�~���cfYm��F���&p�PC��|����|�S3Q�����^�~J�=>"��3���5��v��I�c�� �,�Ĵ�D���zA���x��oD�5^�F?-��ʕf-��	q���~���%<E|���)� �B�E@'�w�tD6
 @ �jzX �D*��j���X{3ϒ����<zU�-�̎x�o���C�ߺŦ?j-�]�ژ99+N��@.���/�8p����w��H%�$N����Q���*��T��u46�6� ��I�J��)�[�=5z#��5�é"x����dUg�\��q���^���C�b�=�n�VC�Q�h��!<�qϛ;�v�����1�.�.݄��Nf�\9��R��!�J�OE�W:B9D�8���C��N�j�wdB���7��V��������$N�rPQ���WQ�k�
�F���Xx����h�F���������-mD2��0��	�3���4r(t�ԁQḅe3��G�{��f���u���j�l[dh�g�~�W�k���*&lp��F-2LiY�� #�X�X �vYo��(�}�4��Jy����1����Fy��'Z1�<3n/$�T�֬ w��Po]�[�d~�G
�����C��à͈���i�A��Fz�<��:�q�L�������1��t�L���<��M�/������!����$�B�ȑ��%H����S/A�8���.��P�%����|Q[S�s(>��jߌ����[@�fL�5k��hR�|<�~̞}�1���H�E8l� 4/v��V)I���\F�ԀWV%�/��}nV�y��q?��Co�����]n����x~^(�Ĥ&�'������g�5b��D~��&4 |�����w"���ͪ5t�k'��Ŗ����26��-!U��TCvBu�y�&(ŕw���6��ȥ���� �Ҝ���zG��h��r�Ib*�r�����a��^U�R�v�NK��;���{pD��BU��Woo�[�3�����k�2�^
x/E������RKDW���a��k�7�>��K6�G8=E��ɏV��� 9�3d�1oY�u���	��P����5u��FE�g :e�B�dR&)"���I���w��~������EV�i���w����eTr���*�J�,j�I0kX����e0����ϸp(�N/|S�sy������ݔ I�j:�æ,l���9���*������ȹ��W\��g�y��1>�^�ܽ�t����R��I�h�^�����dש�FwO��pIoM��h�=���	i�r0��,�H�g�(�/��;�&qKm�Y��k�-vI���a H�~ω�c���s�ᑘ&�dV��Y�H�2?����	�brN`#�BNԨ��I�����/��7�W�Y�0��~/J uɊzz�T������s���#�$�*�37�Ϛ,�%6���j��4�3`��z5��Oa����1�6K�o�k^MrPM����¼|`�FX~��.�$��"���sUW���Ch�a����]��	{}P���a�`�4��Ƅ�!�����!4��J/�m�(?n�>��.K ��Qte\8�}��I=�D���ѮNlE��{h��}�fnC��%�K�-ZD�F�16D��N`��j���~�"DI��J�^������옃!f��L�^�MG�X����tR��X�k,j嚚�f���t:!I��
�`Y�W4��lm�����.�U&�6{� �'Nn��������c�*'	eC弴�1Sح����gd��Q��q�v�FR�[�\3,��Js�"�@V8G���"��u�:�6s}�G��9mZ���_�
��]GX��r�94f��{U�:TA&�nR����H[�5�
����!��v������^�x;��� t��1J��OG�L�}a7=��y\,oEtT7[�		�֌l�>(d�CK��տ��v�����/��cL�3�$܄
�.�O���Qb�`�Т\:�^b��r��,Y�~�/ِf�ş�|��kx�3�1D�
��[@W�rۄ�����J�����6��T���RnS�C���a��Сti�ܴ���D~��tN�	x��^���δqUTXH�ꆆ�M'q�fO10^����n���}�A�B�CYa�"�34V��14�e�C�J�I±յ'�W������7�	^G�����ԖRp��\߳�q�Z"��%<��M�k���dԷ6j��$��TQ�;w��&��)���`-��p���ȏ���V��,���'�
��w��u���x�jl�po��Ψ@�/�j�i*��݊i�f\�Qx\�r4ݸ��+-1����g�vc%]��C�9��ޤm��,����p��zB��C����v-��}�x�%+Ù�1[�{�ܣ)@ѐ��H�+��#�Ӵ,%�fݦ>7��;�)�qBƽeftV�G
�7�o3?&7
u`S��muo��h�m`q�������|E�M�]3�'��Mv����c��I��$��-�S�+�/�sVl��Z=8	,���_�<�:�k� ����=N��E�+��מlv����vz!�%h�B�6�q���̫��]ٳO�sH�4K$�����O�n��
����r���6��m�M�P�Kc������&�V����D9[)��;��Ӈ�5׉q���+����FjG+SPųEb�����]�Yut�=.����e+$��	��="��q궹�IR�� ��]��.��� T��Mdl[��ǹ��X�2OQhg�:�E�9� �S��`�M�]
.=$��b�o��t=�37���Pʹ��6nR����@��?��G�d�z��X�>KO�XCܜg(��P�B%i��\����@P�],�xϨ*�|ڏIe�]J1]����}O��N��s6 ��$�kC��U_��%[}r����K��d'�ZxQU�`�1z v�f��E�]�Y�tC.�O���~���ոC�y�3��	5e�K'��%�m!, Mm���&��$�5C�rmOe��(��"����~CTeV"�|!���z�8r��%ԎÿPY�ס��a�M�[�k�B��J8�G��	٨�|_)��Ì�OdG�2�@��5)0�����wct�/3�e���V�]��PYČ�W	z�a����B�񘢪��f��h�m��q�_n,� �9��Uէyc�e�C�V������]�e6�M��Mr3��W\㋣����Ž����&:j�� n�o�>�7v�5,��4��eZ�j��'� �u>Z�ӽ�h��x:�.�e<�BC��%��g�A$L��J�T�o�B�����N�,ߵ
�2 ��.GN!(,Lq��K��_~D�D"re�:\+��Q#	{��X	��Nh9:d@��n �i=������~��z4�������8ք��	��@��M�;���i�Z6�7�:�k��>��)��� Z��0�Zr3�>#�aE�-�S�/���p�١��@ P(=�v+P�=#4��1߿,��m��ÐK�XT���n2W
;�%������6l$�Q��&l����L��3xouM�t�Ը���f-`��H��s�M�rH�A���A$:��Ub"n WtS�P	Ը����t��=��P��kZ�<���id����N\E��+�n��Z�
��А��X4�]>�ޓ�2��I�%\��ݾ�f�G�Z�B�N`��ҿYT/ս�P_�L)����}��}帖���3��3��U��X��^\���]�������xfdYmVL�F3D��S��62_?��`9t�L�;�67ǃ688O�;#�C�x�x~�i~<���`�c#�Ж����,?X\��w��qN;l�=:6$��L۠^fۂu���\Il��ڲ �[�lS+;h��.�~#bd,W��J3��WpW�w,��/U�-�x�f&a*R<k�����ݕ�?.���bQ�~����JJ�p������r�4�2��9lo(������4!yi|��\�����4,�� �>�0]�ͳԆ�F���^��5��i;A��pl�G<��a��|�����䒸�ԅ[�e����fAb��� �&yR�2OK�an,�BXµ���sV�^��f�2J�k~Z���Qd:Eq۲ �D��>�@���"]5��]����pP�~)�;`<|��dY𘖨��ݟ\� �$[�Î'k�`ʨi1A=��~5� }���tT�S��C�%_��S�T�Q=�15G���O�Ə��eTF�>_��y��'P'zޞ���m,�֛�	.���?�=��u�bERp���U�l�{{�T����5x!I2g���fȲ�{�6��߬�S��S�d�4_/ܦp�F�@�&#�HW�r/#ݘ�g�ϗC]e@2�T��Gzv��lH��%��a:��ȡD�B�)ξ��zu,-�+VO]��v�!�b���|0s�P ��@�����@�ZԆ��tY�n�`�>�Y��oo�Dq>�codU`��[R�8������Z�˦���mJ��R�n3`���[!�d9u�̖��>&�Ĥ)Z�n�~�S�c�1b�F�}���f��C��]qxXɁ~e��(�2=��w�zq�� � *��D�]�Y���}|����S���xw��b���Ѡ�>F���VM'���x!F8VU�����v�s��6��K܆a�d��?qD�� DԐ^��-��ϐh���H��-��������ˋ^�eG�"eK�\�9��y
�dCS3��G�؅�q����|���jX	� �b���QE[�ξ�7YY�o�1���]{10�	ɠ�=-'&�)(�L��69ouG[q'��+�ݧ��N=�����S�]�DǮ�'D�S3/��:d���g9�=T���e#p�t+�o��I�E�ktۃ\�+�䎝5��C	�����T���cU(�"ҽ2<��ߏ	��*����S��<0�%!�X+��N_V���^kÿo����\@��^��ZV�N�זvx&dl����yy~Q^���S']�t
������
l��*�q �������L��D����!4�޻l��x���Kv̂Yd �g@](M�$#1fUg!��ŀ��ȃ)bM+��1*�	G����;-���uN�B�IH�&>�k#��>�0e�� y��7�=���К�u�(��Z]=�r_�Κ�w��J&8H���hb qr\���PP�9�F5"p���h<�K��п厔���S��P䐻Q�Wm���4�푷�/߻�r��UGmr�ښpLF��N�Т�+G�����a!��P(�\��b� vm���1��5�_*8����;��1�21~=���9��+Y{��u7r�NL�+�Ϟ��㍓� �
ĢTo���F�
�׿�^�7�����+�U0w}z ��ҎZ&�Yq�P��
!i�L�W��
��cQ��\���\	�$"���'~>�x�&��^���5�
// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
FvbmDTa434+HSLaxyHmvIY2hHeLm21Gba0qL6C3YVE9z2TSOxV0GAsY5lM2JXjZ+xpVD8BjqfNJO
ofZd4gwKd0BI0LCwQvfC2x2yKthQfZEoPR5w7PIK5a7bWXZrgoLDtY0+CI/he9roeH5oN4bMBb35
17250WvXJdgiNQvbt1vaSh2im+QT90ipjIaV3oyZ35i5uxQbs2VOYOXoj8QU7AI2aIPQFOM3UoOP
vz3ORTF3POqVOSchOn09tNS8pKf6s4DRRSStZZD3j5R7JIPpnqR8Oa+ZWL38qc6vguTOpX+HUO/4
pPqykXDQXiabAHJMd7P8yrCXQXoTM76LBxavXg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
67fpxZoV5r7ubl9KzFKFmft2mkElYOsszY6snFQVdzooRMDx66DWmbhIf93dzS3gnqBJuAUyQTvx
AM5d4er51BGOHmiyNlpSfVXQEHBpYdd1e1pvke/j8byCe1ot+MLuMJaAaTRiAoZhHMfnBnkIZ8Rw
ssE2SfyT0jBDhQsmlZuOuu+//3I0/CgWyWXF9/I7Nqv7Qd0LUHkRuEc3MboqQ+RPLOAP2XkvR37V
8JP+CBxK8jOgnaGPQi3Qu2VfZ+W5muWSXqGhFSVIUddMhTDsr8WULZijlkt4Oz6EcDrQzFiFBwxY
vr4Yie1tqAbt6FBr+KAPlWkLfLqScRRRGAKumI4a+IfMw+OEkX9NsImK3Zjx3Z16Zrcup3hK5V0A
UMF/wj2YEUo8OwuWnQ8KIZ038XwDe0Gc9SnKVw9+EXG3maAFooMdZgoB1hUn2Axp1BE+KGwxIa0a
L6EjBeBRegGVT2kAEk/k7cG6vVckNjav5v4e68y/yqP/85YCZ6aXdPbQTKI1Ch5BD+7vN0iwd52f
tnYcs0Nbytcap3/lCu6/ZN3PIOWR0EY936qObDft9DBC4Q9FQrkpEfOllgWGRo2Lpr6oD/xf2FoJ
fT+o3qVpqcDZ7Nd6+VJhtrtsXPZtbkweBxYSSs2Y9+x0XhkhUibO/dRcavW8vbaSZ7E1hBjVj5OE
kPyQLwo8sXxW7ubpS690t5Qy4M9jPSDnh6+tK1DSw+okrfvYXJf+idFnXQ+0qtlG3JHqtO+gVwyv
+toOPT83HiCxd7zrMLStUSSKTjlQByRGh0Qy+dKO3tCpkNx8Vd5kZLo34j0zLkw0vrBP7g2U7Qk1
2iDY2gKT6fUhrGD9+Dvxqjabeq+jlZ/qB3Z1x2QDo/LOcarnryfTkizhZKO3NgBH1mBtc+CJClYS
6VMYhwe9kBxrdqnb9llrdkQsMpDpWpT0LHpNc6klIMci6PHXR8S0ltIbVvplfJerBtAkeLQ1nd6/
pDY51/7MFmu4/YeQzcL/fxFhJoDBB3MGWYOycQKrgOmEgEAnRGW0FtlTKG34Q9srwlXUZt+LtBOi
wjSOIapTn03Ut1lfgJFN59TJPgGUM7UG2lqJLNoXTQEwXxU3o7iTUawQ1bQlD2i8WqCC1hiMDy0l
miPVe4vu98RmTJm0HTRwpnYLaKZV/8e3AMAs5PzOwHU0xUk8KifEzBKCOAthahtGbhBDzs8hLOXl
y5FU9l/tkZit+G1XWq5QXBmDxta5fcgPLjOInOYicUexZbwgStAfhucqonWsyIPpYJCIOHKhI5Wy
cZchSk5U47Rco+OXzFmeQCBj0kWs/MGLb7baeJ7K9fpYwzzn3ojo0L8ttXCaVRtvYad9xCaqntH+
xRX12k7DHdYWIvanjmQ1D4XKurS6J0armKoNZ87IB5DJ3Zs/15g7tZ23oonWBnINYbe/dJFsuO8t
ZyC+Val8sfvnEicsIi+8++dr8Z46DlDP9cxDNG+I2+MfB0+gCHlzbyeOYJcIlKEJ0wM+vsdHt/mz
67J9y6HuDb5e6YqRZOVYfvo3djz5jt3od2MhiCH267jOuOG+PdNGlvrYJt2HBnAcsyUOpcYKUqha
Rq/FP1dMhbgftzsD0zIzQYiAaVmauXoj7zT5ppmCOigbpUY0D0z/0hnpuZHrhcoa9vTOedjPvcep
dmCzBwcPpzs/KKKzw7k7QStsuzPxXMc35G7IGQI6NrtBuHEGWP5SS+akWVMhUmVv3GQmwxdnZL/E
F46oIT1uamgoa15YuBoqResL25cnbjjjkumRW2pY86wtryIeNRj7AcvOjyH9J5vpuGrddmzAl40W
jjHLhAhpMvoNQWv0knlBctqvCrWXwFNbbza1kJ1Eg8K5mjqvqZ8+Ra9S1r/MAqbl+U3tX/KokE4t
JXLFuy+p8AQRAfDnlretlqtYZjPlZxuWBe4yM0UOxFIo1CRXsOt89PBbN1HisUbcW4TNQzsBvdvA
JRTFjIAaCY1jpTtfDWNwC7GvBZ8XhNRXSIN+K6uS/9CbKaI39Uao2ARLDsYR/eOhN1yVE1lNlfsL
UAOg9jhBBP/7YvJm5IU3T5zO4RR/zsJgljs7Rl1na/yLWwS9CrPSy7kepuTWRhVyFdfM39NOsRTs
XsBoq7n33nZPmZZ4DkwXgonHg3i3ZG2FP5XVKK+f7opvWRNm4My4ArLntIMf3EAxbns4ymc5O7DM
2Gm3s6YM4RrgDbgmfsbBRgw8sufVk8NEvQmRI4WGsi5LW4q+JxoLUR6Dj+IiFW038QydBPTZWEkN
68KUmNCuBlZp8JCotg3tuZwUUVvjoIXL/aennA2d1sGSoN7N+YN4a5ED4qKOYtWHgiKQU/Kbn8m4
srbgxhMYBDZ4KnCQSmHaY4GcMxcA/Bg3lWQTrOEll7E/7rBD4LXbMtTzrhjMwykK5WFUKTGkjiqA
m3GZbmvcy2C8+BikS56TIt0LATwToju1vRmY39/NdsFf6E9wQ4msh7JRG65sn2dnI/LP0Gql6RyS
wOizmnhMUOK3Q/DgsUwKNtlU7dvOgiMPIIRLr0Ky0sGaw1cccdp08yDBtZ1D3K3lNs0+wDlQeAmm
ldlQe2u2kcK4YXdgkT5S9OR66shSIo8hUJ7ouDt3PB6Zki39ZzpfZbb8OWPhGYov5a1ZlsbSb54x
3xq+mtwcfDU0/hjeo24YNZbHnlgznHCbKzOmBZge2vS55OZs8MldaHffU3XcBUmHNQp7UYVNvG+M
OFPfWQzS2YGG0Nk2tx0xa6xC99ZKS9aL6/UZPteFS3BuHUhZ3oSd4LCGjxsVcMaG2H4ZXAQrb+6F
vZSHmYB1nBC+5EyPfgF0uJUFpGIowdc/W/HVCgp4+nySAxYG+EkJulQ9gMf2/fkd64Z0vqd4omog
AEiSoeswU5hp/otocYB7+lWKq47PtAfbScjk5txwutE4BWA3A0HmNK/3mHXjpG7t4PDqCchcztrF
ljoBPOoeLX2k+at8QESO2WiY+Ny6LiUsNwDVL0Tp3yPLoc6+r76HHLjFpDZ9+w3hG7X/Rj7OLDKv
JMAgORXnqbbNVpy2Hmk1IMCyrto8PGeUoGgAqaBEMc4dOaNq1/A8W4rp0daESYTe4VlYI054W+t5
WIwNXXck+rCo6W+owidISxngPGQjKMJJwLgfcPCKltHdS9/3ZEzIWoZ+cCXTpyMvuLv7774BGtSZ
oFnVAydcJtWJoNIK3+KSLiB4LsQS85QB0xFTcG2bzq9zK5qLGkk5pMbT3D7XycOFZR71uHJPHX61
10rEjnXx/TJXN7MV93MnUYXKEaxVcNeAgRQQsEXnlovoIIvtnYFEja+3saeJuB72lY49BLbr5yAC
Own+LkWEA07oYTcU6gUC0cwp9a64vwJqaZlTgZ7QRio0Jh1Jy/UgyN7LLlE+T9i4MjttV4LLARkc
LQ3scM/bE9/NAnwRamVETpS01NXYPoZn2qgv0q/5IROLLOO3lTKXp14NlbZ2FS5WN5IxEr6s3HUE
CzvFAcrh2QtY/258SghrLbiJBj9k2bH3i69MeiIv4+A9oQr4qBNGE5NTFuxjxHbA8ZE78z8KgjaP
jVsg9wXHrOm+9pAo88SdbZiqWteHZG5I9hqjI91l3alWTGaHOv8zowXbIILdMhvkYWZgfB9RR9os
I5FURNf3ceUH9egXPwe8cMBbU2sg15J22RQ3/to1BQ8n/BJSR76WAROzLM7mq2BjpqdqIalqxa/e
iUOhOqZjG+50Uy3J+dTi9qC+QKoj3D5RfwFVPu3/WSg2UJJYzIk5gq8k4RS2msHUpHgk/GRtoPgD
xQt00yZjMNe5aDa6FoH/Vwy4d99rA7pZU4yuybgVPHBQcT456IRmaXtqzXXA37CwL2oX0h6IXNnA
5LnBSueVZ621wLclMKPYZ87HJh5MhQzJMOB/Nroeb88FDju6fSwt8F6F08JQbyqxok5L1oTE5Fo0
daoAs2Z9iQiCM5HtqjzsT/8wnSbOSGZ5xCf+Eem3skM9ZeGppQehohvdvucHggmrFyVNriOVaFh8
2NJcR8efj9FWu14LJeAoSk+qP1xlDGg4VnxW15Z+2Wgzbt9ICEemqxfP1h1cFj+XrGx416MvR3ZZ
9hRc+6IU8c7vjNRBhsX8eHdgtMscZ6lALdYzEBv08v43/pTMPeE5zJiPj0/t97OxnNotGrbnxRkr
H3dfnAz9L+SOKQoZvG+fyc0H+D2iT5x3OSVqJnDtaxLTPAhaD1sVYWciH/1y4AMPTPRvDCShhnMr
xEWTt8oqO5X20P7gpUC4pqcA1VSiarJNepkTp70JLRl46W9nskrgBthe1wkCMBP8hg1NmKe7NjVR
QHMry0Nztf6tTq6Yzy57b5FgrwUWSMXU0KdhOyN9dt2+U/P2phONWjnwqIezHxTBdnrWHUPrPdfp
I03siiS4oGheMAiDZzSEuWfGpIAntes6nR384jAzAd0rWTgaJPJMy2djAz051nnaVoGsa3oXV+1P
tHXvVaNxWcb9aAN1wZ3qjHLdiGQGXefwNbHxKk2PI6k1NZY3UaCZ2NGHP+NrLkl0+s8SgJXt1pp7
u6LWtt6KFRMVqPSpnMNReehMaEFNo1ucMJWBcQrcPkeJ3uJ/dBFEjhClu5EkxcUIgQ5zCHgaD7At
pvcDunNsUe1BFsTbkYvpN2QCDrJPrgPjknqxtT4kHGaVcO0KAAIS7dS0nRzc/9gRAyJRWxBMRz5n
3vJRXOdYluSGMiLCdQNHEmEUhJgBFCiVhiE1wgC9aG0N6zvxgiWjTPG4rDxIszQ4nBW8N1YF4QIS
o+Y96SfNmzaFNu8+AabXKHSiWSAvfV0QSBlD7Y/p1PaFP4dHqpkbs0D2i8SbHJdmznM+BzzId/4s
nIeE+Nex1U0ylDNE2OD9lU1mH1+6cUpSkIe/WGGBBBskiKWrlQh6wMrPE9wgPhtpJb/dB6rHNKNJ
gH+9PoAVArhSnhGOWRDBvHhqU8II9KYwWrnh14/fDwvdFpM0LY6jJcB+jvsRUMc8hkLVHJCjlurr
ZPm8QWOT72RpaVtHmf1/jdBSX/TNVCX4y3Ze+IQeJ4XNO1Agw3v5woMxULvgJlcmjq+4+X9ysPF/
Mm5pfQZWHpEGZDibR07K+mwhZW395I2ux78xRBAki1v784jrITjDw5rvEsr2P9+EFxUe2bOWt3kN
5zhmhYiu7uIh8lDJGKKMwjCBbYuo6qcXWCR3abJSpmpJ0/cTzPZw20UJCrEBE30CQZ7ZINdg1D0Z
0tqdgah55ej/nLNurgG/b7dQDrhXvI2bih26hcEivJDzFCNXWrDPAW/Hufcv5TJGz88gkcInqAdF
rKxQRUobF0axa+ZrEf6cgVbTbv/EpLqR5KQEdYzaOX+O4P51/6lpBBCK3hksxQ/tOt71a5THgOSs
YaNRcU3LyGaRdipBauALyuZ2FyS6EwI4rTFGuM5g0PBkT76xVTqJTRcUmfDweUNNzciNnyXpDGrt
Fei0cAw5Cj3BHNStc4sjPbsLZ45FOeoN5JCVsU9wbQKwkFxkxbHE5jCY/QuqUufEgcIdEozhr97g
9XFLx+VNw5iyRoI92VOvU09vW+0iBbyaC64xTPqr/0us9jU8APoKq5rWb191WazLAWE3g7RcKCjO
dwkrS+rov2ciVTVvklUgQsOBnkX59xu6c//4VOnVt1jv/FvltASG0LqqX3mCA+TL2Jx+FP4LMc2B
VURIMXUu/RuwZVuB0pPSx0DPEuTqzl3zF9bwq0CEfdjFXKJhZhHEzYLrnNjJgAvuOwffzUcZZObo
plZ284YhSe0myofozMlSvbbpGn1AEf3DkZl79skrQM5tc6HJaqZyH+2qcgnHRJdtxrIHogBaeWnl
n99NtAHtNEn372KCF5W2ewmR28VZt19EbPQmUCmaGtTl5fQXTpsLE697uxnBI07xauTGgCLpmIwy
q6IaYL6FfRfp4B9gMT2f1hO+LKoIC8kKFpoPtCZ6hyz1NYNDFlI9leGBbJS+5OTzlNm5My7A5Vn6
wDb07LltA3lvtWgYtAIeYmRsMo1u6jwSJxRwkNxy4g+Ir8hvu9FaIsyfmDzWc4EUn7cPhq6+tfDH
CPuLmK/dg+vCYFwCPl+mNgtJ/11s2Cqilxhi94VdN90px5IfK7KRAV86Sn5OaLNR+APnUNpJHsK6
Iz0i6nB0rDsOb7P8Bdu0Sx3xKujqxQo4siUtjOS93jShOxquazCh7lmpskruri4wAX/yIgjEGT4H
XTCHGCHM+IaeXrpLQE91f2AIYZiDINFGItrin2XRZiywnqDrk8Dzv+bPA6Ukv3ayJPItRQtaIwSb
uFwuB2OrhK+iVuCLCNvToBsj8ywJGqO0Q3yaI72iw2YX0XEuNpInF+3XG0MdG4KnLgPmoPQuzneE
zzDXz2M0jEBCsNk/ptkjI9H5QaPfGgRVfIhu7CZlguP70tgIeO3Jn6jAJEpUMqXxrmfdKnMix+ZY
aQYIdc4vhBTKybsKCuVGoByWhdzQiUiQ0+npuMudSpMRrzLlC3p0LBJwOuemAIEyL9jDt/Ra7+uz
jCAyjaLeKxUZ20725izYZtiYh7IaqgVQSdJHEI1nW3oIG6QvtEu8m8VUXtzyNHLPrMLSPrItPMHF
VmWqPXwbdP8nTdJZf86Z6tl8I7OJcBkxNO/5Y6lFQ5wmFUSz8ORYLh1gDcOJZdbpUlJ+r++ZjuSP
s2BsJV/46Wpzb8OlavbhOuphLiiVPPTAaFQEC2KC1ELmp/4KP2ybZHhpP6ew6WrF23vI1OQ2oPI7
NAINn1V3NgAajah7bc+hAr+RZdgE7Nhv5UfpNwqVgi6THDlomD22P/+aIwe16NQWxFAqGlx8S1MZ
V8CImy41Ur1eHRPLh6IqEX/w45SyDUb8BUVr71wTggoWmV9o6Zox+LmR3fNmUZBIRDRcJRkTmVBO
DOKpspS9jCUbaK73oGvVIzaoD/umwplI9K+sprjWTZMdZTtXqBATJQtuCA59N3qt51GpU/+wGs+8
G2bYeQlS44nFZvGlcwjvPlKhGQ7cyEv7dmzjH5lAWyxc7ApgAQhP9vYTRq5dFYnPU6ZRnERim6rF
2zO+C0+WrFd0Rbh3C13R14YvkjgAV1mxXvNIwtz+lionvcPk7ETqQsgMC2UQV2C4PgOoTMRFQkoe
fpVg6yHK68UyeBv1n/PHHUHbc7mqe5l6Km/7Su7+4BPzFwGJx3M5Jz4wb94ItL6E2RxksaQG/587
XWbAW3RGtYvhKu0E+axG5NqiMpuwKM88X/MZ0EukBdS+5PDdi/Nf9UcMhtWYWao3yuCCiBoIYpek
Y5zKcoujC6xSRpmEI4tUDdzH7CFNcCTFHeQxN4K4hGUzopF6a+6ZpbvrtA54DgOgdQ/uZ5hQLne9
oWpcVVkRojjbE8a6u1lhldDC1ysGIaqXfq3Z5i5P68It87e7z+WDlBXmhFM3WdGORHkk2kuzDV9X
KTUUxBP5QC3j7YDYntfTnbEksPJ79hCreUmEoQKTcBu6hS/te6lLL+7qqeR1qYlD29uq4RoUpGUh
OI1gOgWAU28K8JUkoXDOWijUS0r2zJryItS6GZxGj0GfnNulS7Ty7koqRCe6CO2CyBxc3HZvu3tw
nCCkvy13TgeZEIKLj3koZk0Jea94ZImpD3bB0dVLYJRVjp+D7VRBaV0+az9nFYUf2y3c2FMBg4Ky
/2Cr+riX0irHYWS0mtnTyoIHA8uFrMWZGzHk9soyR4acKNzSP6DB1C56OrIhqUvBMiROkC9zTFZc
78NKd8+TW7TXUAjVMgXYi0Cdw+N6SOov82bSS2yIQ2u1znOlEiTM2TFNjZS/og6lFx4iwzh1n9jB
dr+5WFXz+LtUesdoo8hgDxtG8PJjAKtdh17zSbtseN+bn0+aHBbyc7iNKIY61ZEAXzUqHoWbx7Zw
uM9T0nOM0KIy/LLkp2fNAfe2cE0bb3XxMfAWs7UK4EnzE5HqTP3iZuW1FJXy1SFBd+o4QFsEv/us
BM/rsyieW6b3M5dWTfP4MxbJr8GAwauiNOO2UsqAaJfvn8y/d9Khe10Pe1rjyW8965eQrp2R4atc
P42vW+6ma1G384DEEMQt7S3PeICo5OuGsceAveE+oLAfiK5oLSgpmyxuX5V0MlilybBvLCnSmVUo
/s36fcouUM3ywaQoLuE5hb9VIwZdlWoagvdNkiCJsBSqHw3pfzPKoWQYfFn/jqjiRDQG5+/gq3ZZ
qA6YVdN36I4xZb4SjGuoVLaU1GCNBI/T7dvyRjG7EJ1aDahRG4Q3C2O6UAL8wtswHS76poELDtNl
Cv6nQt7f8wDGG4gvL/OzASa92rQ//BAmwZRa0aTKXAfM9lOAXofSiYaKbpVc2s8Lfw7oTTEZodb5
p3r7WyELWZVxzHwHoqUjOsDHbCb7x7MEc/yD0nnz608NLSp9lE2S/Vwc9hV7KNMbh5kYQaHIbz8E
OcW8KsvpiBUB3wv6qU1aiUy/cId/IDfyJPcD4ayYkqlF4Y6ErPbv7YGrrDD652aVtjcY74ETw7Ib
FwPr7jHIFjjcBQQuie2r++qTVM3Xr8G5r6vUNrPfp5Po8VfrzM/OwqCaTOGLr/EijCbcMaIMVt1w
QNB0yfThoOOu7eCMMvBzkK4TKMHTphEapvoHN56v8gelCQ3wUWTNKx134AjpNjiarfSyg0Gg7Zek
SIPTmLCGDJw/BanOoGzwFj7hniOrAYnbRQXSr9Wu7QiRbDx+a+W1wbcYjfjXpWmLCev08218RKJz
UuQtbTPQrppeOXMagOtZNclfvnLyVoV+NRIbF6wrIugaxOcf0AC9LiVIrb4tp3QdIcDzsYfiGaDj
r4/rEfRzo9cI9bOViEHpEuexz50s4GVFl7n1FfINr9glzQ0ov6Ea46uqEqpovjZ2DTL3FkCor8It
a0599TJk2POFiDpn+3uMUuTTYDPADBb2/SlW7RVPfp/ptADFz/mpWRXuC+UFAi96zm/CPByPjYEN
EPmhKdzJQBZooXc7aYHnqNEJEeAKvENaJ1hU/3nArk0gQ6eanb71xODZyY8p4LzKFTudSfUFWZPW
5snWPE6HFlJQUwjRf8HcA1LrlHwuZVV+34hV1/ryI1UTneU1PTb2+l3nFtmLpdQHQfSqdvCi4zK6
2/2hT1Mi8hzhSet6szZ9XwbvmCaGmrDV7CRw3p1xmZnbWK4ybgsAurGIqzhX6BF4j4wljmZR7Bi8
Y3RsDVdDrAMWTe4dGho/mykYXnSQk+N7DKaNS2jVUiju6BqicqEPsYoJ9npS86QGYLstgkw0Hqjq
jKvhdfgR2heOvVzjVX7MIyO9ACP9K6r3Rbdr/ddIBGUAVWWvQojAJ8O99t+onO34QwEnDgb2YLs5
LVuKrbFbFzOIqaJFmGoBCB9KL2xEhcmsmB20IFtvoDWZNp5/eWiE2fpJt0eCZgEUaRsTmyxyok3h
xO7WmP7WBiwiI5QRZrWUcjbCq53zPIRNpkK0biT2D5UbyY9a4NohzMRS5UI/dJtHASsHP8hDqjoQ
hufzUcsnW1J2iiVDETPO8DxIxVlsVZ9HyOwZzgbSf4QCMXN9e121xRHL4niVK9bVQW+GeB9FeVO2
4uwiSo+32I7xGY11qo/rIRd/+GyQjDXAWg1T5/WHfVxlx/Q5RZxF72rheXAs/5auLnYoDTmqn5oG
A3tCrqHUWWQjhYS2aBD8tMeAX7rGyw+mYUCcQwXyXBbhSmCIIXEbH4rZy0mEQYUzbVnNPzh1ox/0
p8rgJXp2xBqHKLuvYlpC9mONnhoEPh2+cQ2iAcHBB0D7W3rFnGaG6jqfW8Q3L45xIcmjMfSwJbda
xAQogS4zYY8yaz8ehe2GZQbCd50pq4Nzg5lNn3hjKQQip6FXzlC2Zw9xEpbbYlRW9KW6JPPca0il
miXTFyvG2BiJ99977T0KcDPXi97Mhi9C5iBximmXYBTWO2bKyA3X1Uc64iWJWrXH+gDx38hUpU+E
TYuzcELdO41SzmdkUzJW12XoQHYXt3RNhI2ST113nP2BHN395v2iAZGuaz1w0TKMVr6JsQZ54o9e
ARwgaQmvWHHZUnbdva2hIJwKRHLSZvhoRKwsiKn+cSHYvGpS3PFw6zfu5QdIS5mNDoxCNFmHJ6Zf
+s0u/vg/r+JGIIMezHMEBSYGhjGzPqg7vzgeH47bP0BIWdFJtKkk2uTI6YdjAyz/vZ4AHjP/11+X
g4hFlcRkUhF0B2kFIME8Rn47r5D+SoW6DFs0gIvdecpfwD7j3VVY9goN3vTNtproYsy7I9LVcb6i
ahZq0VvJypoMU8fXMtcVeqLtDeFokXImijEWIkZNUNU6w0NTeomEJujeg5cciqXSqx1I/rYfNw1f
SciNFG4BYttnvfe9W1LbQdO+Iv1oVMNkC94uxlms6J6Gs4Ggz2egoaskXfzw2qeuq5k/H1hgRmVD
yRQ5BsYE6AXYNp4ZRDu/P3+TvthlqRUapedEXcMykKyqLal4xUnjVJhNQJ7MElNioKa+ipmZB8Ys
ZmOwJWenUI9JcvpDdxG8FkbKHiW498/4NzLp3/XZQHMqqZIi1sEt60frrFukGHlzFl8I8tp4SBEM
4E2ToC0I3kz5BF8yhPmefoUQth5u3eq9epFekzDgOCljYh6im/xYkK1O91Wf+ESyr6HaKKa0WLM1
eTG9Qx2+rXv1d7ayfdoeuzFrFQ5qW75mESO4OsIRUro8wnLcN5cffZPu/JV9bS6MUowuM4bt05Ll
PyKtQ+5YujRfzZjd2oNHfG8yAuOL/Cu7wXmC2XtcMDALkvB7NAOLopfdd0dalPDLWADN+zllLGje
88H2nxOut22toFCxo/LoAZOpIpNVNiXgWgxmiqOvtRE4mKAohlGIkRCPgiMaFWHLIMNftD3M1UWP
cn6AcnCM+dI+WYnqmjsh3EbyvZWdJCM+7v+R1XCAd0adSDvBqeBbU7DKEUgGSXHJKnEscJKT9PKy
S+miAQIkJbMUxdWCfoh8aSmgEjes7fNpZHHmOHRvZe06GlTgOMjA7rRdCm7liytAEdyftQ5nrtdG
LsvRDagFLTVLpUmW/uSURbEt6azIosI3Qmxo0/k/gTeAaHb83/wVP4911E7Q70apmxX5HKEs/TkM
2uOF5oWBsbxAqnmpxwRKbUUbHRt4YWCHK0vMQFHtvfimERz5i2vmFT0v3h7Wri++VhthLuSGZUZ5
q5ppzWTZ8p+rF5OXLn8jzYZ6l1iJCwq24aSV4I3ily/+dE0RGXMeJPORfPyG8ltyFEb1cdXKMDNM
HijneLiA7mSn22n0Ulh7f+JwCaK8ae6/yvOpeeN9rimvxVmWMnJDTI+RwhHM4NdS3pvw1XlrKq0L
H58I6oy4JvCpOB7eTHFdFePmFhvT3cOueHBy4vINgHNMajSBthf549/R+10U6ZNi5Sb7IeaHHlSH
1D41WDvknYSbrsCRGhF7KwY57J8qH48FK+jsZPR50gZ0TCXDXGng6ZI/IO7ToDcGtWoVeTkGw9FK
SVAZnZhFjRkZRi5gcB0h47x3VEZvy856JD789YFCB6W+W0a65BrJVsvIKnJCMCCezOfCr9/2SdSN
vV1oWt9dNjNK/q2by8CxkIkLaMbzBXfDNy/Cbb0erkPHbbzjh6ErgATGhFyIPr/TDC3tcogIAmgA
h8Q/cfCiEh92US5RaqisRyflkMeynitlHoXmvq7G9dE4bnUuPZ784V7Y3fGPjHMZg5O22Lx7NNsn
rYNTUL3emMtjgdj144g4bDitGnGtPMtIj9wQa0IaRdJePL/nvMnf2SNaDq1DH14c8GN8E1LMiTZ/
xOpLFUIS+oSMeMFTZyHxKZNCrl+H/VDWYJJMs0Yfrb4a4qzKE7+3vGqSWdob
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:25 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VPVuewdCly1i+oBTCNijxa0K7j2qKXrAYx9IDCNEMVXlzoFQNE5iLEpxjy49tMlK
5JUUWvx/3SYONRRF2X62zy5vkh2f4RnOVzYAu4tEb9ochElUklkGYGa4NanNkZQe
Uum0GzW7oqLjNtLrVJw97phQ146R69Es/TKszBTHW5U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71232)
Mjx5Ztx7NEObA4jfUbbhMotza/ajMxu/n85zoLM2qXwrZvN9y5z+3BLPxnC1z2J2
vctKZHrv8U82FTO8WvgI6a36uXKTBc0tz9+HAF8UTi3xhJEsZQXOczpjkTHTdmQy
MKNAmg0fpm0OSfzi3+j4UYAipSiCAJTRHEe+7hy94H4G0B0wCKOE7r2/E/Ft4Dzz
/pLnLpPwkqQheUlIbk4ufmkUyySBvb3/uKXDRYxoBsxVIxhdXlpKUwv5wVBshG4V
+PeG7mqPq2xibnshNJbRCjmXunwYgps54Ykykog4rSx0d+DW2uexWmbIc6WmQ/4/
oYBDzWUK0hT/OlIu7zigVq5TIfH122r32VjQ886s8vfIPsL4KW6Gt655GXODeGcr
hGD0nZRHWl8vBakmr9Leh69Xgs5X4MiP/SVztZxWclDSzQoBX+H6RSYX9To65cyT
6nuzciuYIOEwctCve9HUjFjWzIsI8UKMbIDvzip6MH6exPP8g+vvUBjQZ2VP8uis
5a1R5ALZcA2jVD8aNgRae2ZJeLNPazdFYyET3Mfwng1My4hzJ6BSGi9gLgGIDmAu
Fnt/fPIfBzRcnI8i7z5lLBScC4vXMlLCE12h6tjqJnlqg8PfvwQNKp8zp8oCBIH2
diCjt/BKVy35ljrxFo8x+9jHk/FCw0MP06eq0ZivxojBSWHRxFQVmAAw+Zty6X3w
5VTumhvorGYW9Pgn6/U5bWC5qdpcki6dAkftWJGmR4nK7qG362euLufG+Fz4B9kS
+KYxyNWQ4e0yWPTdMaDfQJ+IvmegRkUDgEf3S1MPIRZ5bYgNbYmqIIwmGYbJiRjm
xWL+kEp/H8jCqEqoZu7gnJp7K3P4E/hYbx+PsVJBEI5JCgY4vVRH6kDNkuOrOxA/
Vg7L9/a41rV/yD3AjEfy3wW+AwsCtwOmEeFdpkD2FdMbzAm0S8UfDVwrGM3ZaTKV
e1i1mGhJmCSnCM4BXtZ6bPOj5qBf8jKdvJtmzxdW/3zcSEIXVOO9h/0TO0eBj+Pi
25R0iF2rudc1zlcCHcSlxdd4DbXxA4UlMbGk1b3B/pVzAHe8P+AuoreQuOOaZ3P+
PU8afzt5ICcFvIVgFpyc2goD9MEFbHvegVtuXEeVu1jZr0p7JSq4tsYMY+6BWcz9
KQB6CE5E6Tq4iwSK98bsLLCqqwJ2AR74V5ezuA3dc531oBRI1W7kkATDLGvIf0n/
PthopoDrUiYR6XNq8buQ+J4hnUWLddXuAg6wIBviTnzWdmX6BQ9CjVp1yizIDp2C
Hjq44zIKn1rjtEf0PvFKcE+GinoaLFVUwvwdqRSzuqaKUi1olOmL/kzLIKl9vxY2
rH010VN377blh7iXV0hktzL/O8rLnA2IDptmwZUH/+fWkpkZ48455cR9zet/MTY7
VLbImJOFC+cKv9kwmPjm1ytGpqC/bYnSFOX3YU4ebKwq6IVcV67mh2y7/kMDFDeD
IlYdIuneHVGphtVjc1TbVFpr6+76/3vw6VlzSK+JCy2Hky/rwhP/zWV02U4U4ssD
HgRd+CAyo0QATWEXxkXudjZIqHTE69EmjmzWu8GaTo4Gsql/HOXqZW57mP/zKbO2
/RV3bOMvZqhb7A1h+mxPwYYYApYSFbaTu/F2X5Vu1yEQKk6/AGDBau14ZGebjqau
1/lX05KdkGDEryrOi951wKW4Ex/Yi4wdzcwVMfTeuJu1copIkgwautj7zNwGnHmF
TghFiX4ue9I/gpFjgXISS+lcTXepKTELYy90ZsJW9vv/ERn7BJpnEiZPEbBwVqgG
0l6mcNrA1k9QfH/irbq5HszEsmqT32Si8VVpA64ACmHWlTakEIHvNmTMu1RoawMZ
2EFIQIMgLNcgeK8YhXknEvWoCNW7jRlf2KYgPQNDIX0lUeTISOxpjBhr3yLyI5e5
KVjqBAwF8RVgdtPC1hbX7HbagqkAYzxBcrmaC7Xxji5BGz541c0r4IzLh7gtT4jB
OGX3Yp+C3X7tRebiBHzlb/bazxd2KWoCS5HK2FehDEeDjVdXzSl4PbgheAhBx/gc
tVioMLIEpGU2TE94NJw32UwN+i+zXfGko+6ExygfmTzQADFkW8UitXPCvZcyx9DG
tJqxUaqMlH1C67ux2HtbDVAYXXQSh2L9CW4JJFURMJIkIUO1Thv6T/Ceq7uknAQP
tXHrzDng2vi6GvpiswgEL8FcZDDtaYuW+dfNkM1STh5SCv1ljBplxzfpQnTH/KXF
jsPrOPIEc0dpngoJ/uXDyAzWRx+eWRmeCxnHLdUB30vDF27ruwK5lsQgCtDrH1Ez
y81sddbnJY6te1kWSwM5dgauV9N4bCZ/8aRVK4BlHXJdQLfZerfksy0mRfyn1+sG
SoZg7CzYjtzn+2lGsNRfTsiKbB2PLy4UQHnPfJlXvOkVkH0fkeJt+Y+3rIe4VSei
UcpJKEo5szvs+HnK3m9dNKlak+VgWxqxWgIlZPBFWzQJOE7YczLjXGBgO5RYev94
LEK3xGPNm0THeZKnWUCt0/hIqGJCu7k0oY6HtuFf54UzPgZ6/8hJxZ0G+KAuI5MD
lD5gwBBqzW/UH8BlZ7aasOIxz/Kpx+k2nzFD6fIGaLQeSxcq7ioJMxWT8z33+vNl
DnWKzgOPCdS50o+DDHnKB1uPg+xmZ1ViDRVSufnKfEsvKW/xOAX3cKX3INiqzoN5
VnwDdN6SV1G3/Dg+XZvEHhpZ0seDmUrHH3sAxFDelnVfrUS4Yx2ZZqvzi3SwB1ya
g/WGGS75WUjSaSdwCxiQzZYIAL4wbXmXGUcPO40IXuLas3w36H9jVO7KTGDgfRXh
6xf94A/ZF+WbFPTe2q/ejp73aJ7QCzf5oJ7BbdHvcUfKZat0uhiudrfo+bp7wg+P
ZzahSa+1SsFw64Fac+6AMcbBIzHI/HmBgB20k1aK9plaL0qKCWyaeKXf2AxlHL14
F9UdyDFRVbnNaLwLJiOhP3Er2H8POkY3it8pmGsHZjc/WvFxQ8Vw7gWomUXchVWc
ccGXwMMFrVvmBn7Yd1zecLJsvuNh0n4+KKisYOJzHK+45zEGM4xxFWt9PEmqN3/K
aqnl5pA/1lJ2GEE//cqfzlOuVx4zP4Um74Vq7Pab/8RTkcYAZ471CmZzYMGAZEWU
RDdOdZduph0PLqTl7LclUaM0kxNrUi/WSHjO9s8Sn39xQNUGP9BWqQwpOE883i6Q
pzgBI7ShcYMjWP4vA+rh+IaEHtakkTwE7Fa7IpgwPKnXZq93xsTa5jIvj02oVXk1
Zk2hlVefqG+mRG+8UAQs3dWTVZiTlslkZPAEDM5J8+tCzqqtgKe6shNIsBeFKLLC
oAnGACTgDWfbrEddluKGdrr7KvmYYEaUqWOIjEMQCUw2xgj7TmU7E/ZUGHiXEpNq
Nqkl4pFOqTuo3vwDi/xvPRgOmvQANl06r+axVWVHrbNkgVmezM1VQSp8QgC4qVfo
abSWw8LtjsEEWNzRaHzzt3epva5nkgJ1+iaN1K+oTdtEzQ8NS/Ow7K03djNLRJ23
uFPCi97bgBd0+EVFXPOlQyUQC+cdKaUjfkLohqq5QuH/K6r1VpO/DospdFpiG3Hb
rSSxyvSmsTyS3cA5PqslDFCDuCK9hLI93wRxrmfRNcrqzAR9xpnZVIns31BkW9vC
nFRayQN5AYbyiMkV16HzlUIM2VgL8TJwJ5fOe3Zlw8sda5z4n283iw8B4GmMJAsO
be9OBcUYsUvgrHy0Wxo9v+PitprnugKiHzfSEnBuea3EI6D354NvbY5aQEKK8A+M
CBww3QhB29/t8VDEyOKQFmv3sRpEGlMWThY8ner2xYkiznjaddsFd6pjhSciK64p
uaJNKRYlkywPFXz3QIYNbxMHA6ZEoQa8qyuXgJCSMhkQqcWq2K0KriNVk3CbuhkP
LCS6rWhl9D8BqpbQkg7p4RaVpLCy20QxM+7YXL4fFo1Px52N7MAqnxMjVMhjqb8m
YOQtaemTA/FmELpdYLQHX5WYpoRoISHeR+TM363p/a5uBpZFMiy0aFvo4wHRXIFJ
RE/hD1yJ2y8gzI+JmoBek3yA20odgKxlTBjEie8ZLM0mppW0EqhfryLB1TFNb9ML
xlYrFVUYKd5sy2EAUPT7+JIqi+SNQZzWs6D9+iRWrbvlcLwiSxpmupi9whsYOXMu
J9eRXUMEJHoTyypwCpaP13KNT+UthR3y/rGVQ10BGVrBLsV94LSdHq1ryuV9vfOS
rN2dO88AZPzKIFuCjpLpAM65rIISOGzWcyXgNvu2s8EVr2AcYodonXH3aB20I7Q+
QoPMxLOL3i5WTgKS5EAX/VWYVt51jEvp+YWk/Enap9sO8u+8xDuVN1ZzY6fp5C8V
CI52oe2d/BiQNzlGeFak/2bABRHI5ZHEB5iYW4e1HHKUCFSqSurynfFlaYZ4gDFs
tUpuALnKsTydwkAGGa/hZLGEClZQMs1X18+/hU09emQbOigF+Lo5Aybt83mOuFHc
+khoLV2MRJ01EHcwk3H/hYqpRH89/aX1iTM9S3k8+GvjZlOkWmymB/+8xJscpSTk
Y2bgOFIK94bm801haRt1ZHQ6QlUzcxzelBXLLLlRrkH8xmyHdqRnKPHx2QUgJAoe
jII85Q5Ksf+9DqrUMJlDBU325C36vqCL9mRvP/9iqf7NMFmVmD34t+Zsz++BqTdo
WqxvOEg+nOrV+MD/kpxip0/Pyy9kg+iZEZENuagu99hkR6iCa9nVtwv/05VsIJnr
ZBojslqLk2WZUfqi26/2MAxE8U3Hojm1cTtbc4pOulVtAY9bdHTcpMazJB1/zZEj
WE/poQr2EXYxUrR+1wwaI/5zdIm3V2iLmge+f5jOrk01JwVXS2fZnGpHyfBw4ITf
PneP9BJdVImH9j6f83tjrC967PUI+W1myAumS7SDvqEZAJ0+iIkO/jax7nXOf8ky
RRH8WUIuyS+kBLbYRZ+7SYtmQ4uLmJl6wy8Z9ZDtR6zk/+t52/u4r/24rFOkBH5A
+dUUkA03KYogCUnNiBvL7GpO1WZbs6sBFDp1OmYdBKH7eGJHRg4IF2dUhlJYo9KP
EShtlFVCfzs5aSNSI4yqPlEqHW2f/BYxY9UUzX87SFWkZqQ5V6/VPow7pEgsTjUz
NMDYhsbnKbze5dH6c3TkO3V8UcTxC/A+Ld1MyvospfNW6H9wiXe2LdyGxtRHZzBL
bl9QUKteXV9RZKcZzrOV31dQ5uXBD2HkCP36H7kEvGlTERMXbvs8/vKi4kfTpLwW
TY4/gIpNWwtsG7HCdkgl50lpwizX2+eVEARnN9+E4B4BSs25ak7EVFhIdVJ1gxUV
plHsrC/UgBuHesg4YR8rGdOVvjNsxFvNKMS9fn/oxUU/1E1fC4QXKuw72PlobyLm
49gVVo4DbpXwHl1E1MPV+NGY5X6q/MhMuewFYnVga93l6Qr86kdRaUX2ymdUEnZj
kxFbXFPvkosv5jNxbEhrcCATwFG/NRRXFZ7adZZuCEiLVo4IORbS3J2hGhRUIsaI
8SjgN/ZcvSBCZhjPrdR2ATpuGC5Py0GzooUQQOP0vpZubmvJOX3eVBmspUqwlhf3
Af1qj66JOBTG0Jy2Uvi4kVR7gewnpMO+uJNQa54pMG9itujAT0hKHXFRhhcXjq6g
ewygZeRVC/+z9ye2ioUHcRuLZL0vyBTNK+qIZDGk5eRQzRFe05uCuwIE5lWWy0/X
/NEJm0wOqaZwnzmFXp3qQ96G3uuyA/6ISu3THmFIeH+ucBltevnE06NpleQcYMDu
v5pAirx6+W6fJrCEUXr00MLr8/3wMwwzUMt1AKRlvjXZhuKE1AbvnZXZABdpZfCi
BfxP5V9vq1l/LnAuP5OFJIL6uUVDJ3AuX545LP7u7PpM/3ubKLvOo8O6i1HsoEnP
fMfLRU/CVR01Yo8qxzRYRU4Nl0tap7OXohEGPzq3eYDsnzWImzx30+nt1Vqr/F5+
st/AWq6KdWDGxQ3aO+35/wiG6K/kqBM5beJEOJfjW6IesXu02w4wZhh3uLMkCaXG
jV8VKnd8GRiy+HxoYCvf0sJ9A+ORpYgF2TKrZhixqY5uD38M6Xqui4irJXXf64Qq
Y8Ho6aLQ49z6G/zwDolSHnToPN/pVyc+jHOiN/hXaNrkOqGjHOgCXA0Bg4Fu4JOH
T1GBeVjl9Rhfn4FMi//AXFFyKj8QgPEyS9OM7xanOrIyNUhwUCBRLeseQ06BBkMT
LIROdgSDcIOY/H9UVbR9lJ1WSURnrZetF6nG/n1cleVqqD2xkgFVXrqaZ4UzRpaT
eD8oAVNFjvSHFwAu3UvQqGewbx+lH4BHppY82rpgqqYMf8kOCmf/bnZjsVWqPmiM
Ogr9hk8lC1bsduISZd0aRiu13ctD7ztYtho1pX4mdCasuph/+Xs3/zc3PvRKPwM/
jmApRFuEU+JKf08z+gqE5wy+0dFK91y2lJMmtCQjGYx6XV8I8eViy+bvQzjlUBm9
fqLc5cMNK9DS+GNokdiZN0fBjJKad1f3UShS593TlYTQWJCcUEf0EaExSqsruImI
TH77JJ7+oOtEplo2ueHQqcRQooKpj2JDlxBwl42/PAXmG5BXJ8MxgQLBU/s2ZPUi
NrhU7fq3N4tjPSBZOzcl0ZKFbdjvswaygDRRsMYwZCnrG5Ngl8l8hd/wt4XKaEsi
stDDKk+nu8El7TroUv0VKX9ufUUZBD2hQ9HIjnJP9C+rFE7TF1nuhwHNlPMCOwUR
Gmax33xRJt5V7aLHFAb/tWnzC1A7j9Lpz026oM9hqsFgsVaE5IXBt31VkfR50OqE
aTJTyWLlNc8jKH8eCjw03Ur6xInNO42+zfVKAKdBOTfo2E1j1s6nlyPZV8jJx0sR
S8vO9MWLLuXREcBJ00ExjeQMlBeq7pBfoHza1rHPW7i6RZzwmURspiIivGhEitKA
e7yFviYeoo9W5jzAnLW/K4MDsgZGz/sSyDAaq7TqHvKuYfUHV5/9incbJpLzU2ZX
OTn2/niFd337Mdivkzt8iRWgF79MmVmDCitW+if3Wdr9W8igQ7XQ6KQFBhj/Wpgu
t+bJQ3gxDYX62/n0CHs3WpoKSEJP15lgEmfkQs7C73O4IcggrNGgnSQLDK5o6MdS
FdSq88aRdA6r8L85tLlLa1LhZO80lk+NOgK1jm2Q4Q8NTrJQRsalDTC0DMVpEjGu
1d363n8DIFQwqJeT13FKZeo1Y5SRUkaLJyWcMoNPzVAXYyFJt9GTOgDT8SfUoU3N
ckxkVnF31kF066cf2jcOAeFwhWF21JBXRzoLit3acuBxF8th7WYEgktlCds9qZNS
3w2VQcKKRVw0DN1pnMr8hX2H8rJz54oQu9JkF3SImr5YOOIGD0mzbyV9VrP/3LZY
qC05TfR5Bm0rpLMCc+iXhaU/I8foQ6TnEoKvDa4rt4xL4gvEmZEok+Sof0/fq2Ar
+7socCBcpWwDG0FHErK5nXAJdPQE8xz8YUcpGaaTcrke2fzdXZM2hIJVKmDR8p2Z
H3dSgt7ehyL+UbHUu+p1qAjl9WMWoV14kxGeVfsBjCwDKmjrxO9j19LBCCSMcDLI
NH9lABIsD5NXiDv4briKw37TRIQ3nSZQrNf0AXaeHmGFvu3xBja2+l6uo81cSOmg
GJtkkwhWRo8kxjfHA4hCTYF9ZJhz6qfbg6eMvqHmfthraNd/sfKjBwVsA83eEuY0
Kdu6IO8LInXUfVycUI1eedcks/MuICmaVb0MTpE9ochv0Xvet7KWar8E45aF9soU
ER6QCxFLAYTcZOya/OpDOUqOmcB1NAQ8Zt+RImC+gHaeChLSLZhaE2KBg2vf6Nx+
fsABDmZOAKae70bxnZ8OjsdfHyYEkVjdFJCQzz4wX8wlyLkUdEIN6hmL5d68W2nI
5MhFNriUiCqeqWuH277HqBC/zOQzP7Kj/j2DFhb8GyPPqursqqpEhMn2bBezIqmJ
z3WH51Tnh/IjH8GcliLU+QZR0W15Ogkti1cDjjrT7qyceUPuQKJO7qgLsPsPRMDt
fcZTfr+fDaLW79bfHLSWyVz0C/nC9++/pxTarfTAXmF3JZPea38AsSSBRZztD41K
u4xfrDDefxBbkYqJiXCuLfOylQCCVbgqH7kSJvSHXDJdaSba6j3/fglPTGoV3w5S
PXkOWJphysN9KW5tVR8bxeKd+6REBAj2NhLWPQV01XAL58Q1qwxLyIImHYZ6FNxp
dp9Hx3IlDgWr6Syn12AqcBNtzMQchif+XxZY6AjiMuD3zA0ffTumGtDMhpzt/obk
GsHc/Td7TNSjDum/m45J0uE5B4UGb8Rk0DxngGndWD5ox6c+s7+DoDfyfvW7paQk
J0lv2ug11p0BvKuF2V7Ij2EWfpz5u4fjQyOoQyT3VnMVJ0hVK6Is0qEajAQKXmbS
TOt4pY8xzN5kUYtBue5xPXDeUZ6vOO3Qwop3tCkfc61NHFPOoyALx1Gszn4WRYx8
FPyJD9kLJ2tThQH6J9ezETirBZ3fBsk/xfOi+MOc5MgZpgeSFaXhxNrEeSoDvyvE
QGLtYlNbEv9RNzKdy4p8QEoOhcgmUuAI2Gn58V3DRRlX0FmiR7sXmSWYolizr7bD
HZx5Ilyq+N9yR0p64ns7+yn82Pz6t9ik1OyT98NcQ48kjuY6XYQf3hwun6QohTk/
5w6s2XfgziZc31+eZT/rkoTO/xNqBHEm5cDaLXCw6UuKmohx7pVdA0TLBY1yKiXV
GNpOcCJtLOtpHHeNhp04l12klUUb6RbzAauI/09Dd2qBf9uwdeEYqrvXgucLBQTR
zXn3WCdptyfG+Ikdv9G1Iqjz5NAmRRFpfKIFR7uR78BLaG8uKsWA9AE3jgPvRjeM
G3+QbQRFh1jJKY8Egst7apUiNQVvq2MAqVKj+KzAqDlV4Vd364F+2LBuLgm4qdZ3
3YwEsa1qIEHxbjqSEAwkJymVcz7LKIDTZWbllttT20DAVLm/WSl0OsDxChDZoJKT
FTI8Dr7usXydyMIHBnRFk/8DgS1pFCaDoVgDSiN5ia6acELtnWrD/Dqhykaq3zBx
80+jFxMxRNHIDLYxvcfpOgIS0UiuCd7tLasjPtOK0qc80t7+vzNWQWno5BRf9bST
u4eXR+go6xuB1x8+N03ROt7xGjteURnOB48s+84fQbr1Y50NrjJa1ubWoOKlOr2P
NzNl/SNt2olbO9vHsBeFzrTBK8+OT106k4XUuNzvyL7CVfgeU/790IdLMigD/NbO
1cpoQdn6lxejslNAceX0Mn5Pj+0x0ee2EU13wVtPBJUL/5f5CfcpcUaiR/Nl3TnY
s1QPoLZrctvYThG5NAsbZ4uKGvq3MjYyOvu/7DUU7G0wVv27ngBHHpQABdDabUmG
dukd6Imfq0rSS+vbNAVJve7CvkypbC+AQ4S/BCGvI8HN1NO2Ab2G0SrQRXP4MHVt
TnVnepgX1pc6ZVQjxQndrE+QLgJOSJyJuw80xhwmp+/iSsQuOHig/rfYZfPOlWdH
0WtvSgvV7g99UTrawZ7Q+M3vx0k8d+EGslMhCAirxSNn1tiNFCpGq1XrpgCmGS1z
jUQ7UZnnRfj4ZjLPT893m7sx1kQGf97R26Vzfz5wfXqK7XI2BBzoUN1ka9Hhr0J/
MEZejL9DKctsVmAX/Et61tJHYOnxk0NeZ5HrUM9uXG+lxPdPOtAQp5/aLIgi9iNs
JJDrqIDrhlDnFj5CPu90K0Z6GMWCjs3PevRPaikHO/a0i+sklg5vSghEHopO3Ysx
cWEsk8QYdZ66RKnpE7n7ELTuS4OnLewhO2eGOeLGoAYTsmbgluvGthcUkcNlCCC2
NMfmdzS/IHXnPDhdiVqcbn5zv00lQwtOFmOyrHbz+5II/ZzRjmrUrjdzxXtNLYpA
5TjG2+2UQsC1OiOlwTJFWi63YGHoXdl+h2XQ64iHTbbZdlDFGZscV4vKgPtJimz3
sto2pkv7ddvQklYQ0WG4sP7+AIwKOFrnPH81VLK2grAaSH6jRS2HqHWlGy6p4caF
ss/I1Z2RhzHCaKf/k5yvT2oU2VxHQbAGaNdCmFyKcPi6gVZV/7XUAeQkIj7LbZQ6
NX5gJHxrXcnaH1n1meZlGLD7eV5FR9mdQvnZ7Z7MM+WH6DgA5z6c8H4M2ZmxAQow
+lGPqVZrXL6L7eCoedAlN7zVorGYI/nV47msB1lMpFut72WMUj8BW6VkoSktwUNU
Htf8mvCjqzvyWH5sKkh0P7Azrl3U2lzJlR+nUphF8Q7+eMKXbgMPlkRqEzKbDJEh
VYEzJcWo2UxFtewbpwH5BMogrsT1VYmI2hFazudGwrnePQMjLK/DfhtYVTZPtqXD
Nf50DcTQt1VaeWpBPwA0MKvF/nGkzmdeam2ivAJ3RpZWqXHGz5zzjbEsKDWpOaQS
KLJt5R4wiuG6h3oMj4C45SszGJ5HT3T04heEyX1HkdlR5BoKxpJh4klVjc0wsn4u
8hjDvacPUlV4WX/RkqX9kpHmudgSvv18GK8aZpUNzi7ym0IgNiaG19AMERSvB7dl
1nvfnba1D0BJLjq+BdJJC72cCteqXLUPNHRBMu8aHeP9ScGpYX5UVw2+8spj29Kn
CK3DEHXQlXxCFTiBBAvhzykqIEkrtoPENo/zcqdmFjLp2nxc5fGxi8jLFvvbb9kE
ydKQkZLnxb+XRoL3Q+YbV8HxYCZqBXORqamMQw39Hh14AM3YBttKHkl+uWl7K59f
9f+ByJv+nuZTFc/YHvzNPadLqqHwisjjNpgyQocIJ9P4cAL0y4JSOO6+RXH1RJ64
AMYyn9v54SmvtDh6FC//werjM3NfisWU0zlIWxIsKsOHh61y3R7eQ8GcGNb2QpTn
j3ghW0gNRWlBkVgPgJK3E0iK0+4lMpSXYP7GNBbVjtGhVaYSyeFXEhOyqysxLEAh
CtDGAR9hl4xjNKbkeRKjTXy42ifG3EnoUSKiIFzHr/Xbq74A/ZhRl4urB6vFcZbE
m1za4vec332pklrMDECXQXMu2zBmLiLj2SJB3xhNE4fsBoXerfdydCKqZ4tdsI6f
rXTrrHV2bUKfC9Mp6rra97LdtZaqBoOyDnAqKNZ2pBfg5xvZ5LJ2xJNEZN3W6fT9
RfELMo/OI32cPyWauFpNmqPATMDjhojEBkI5qrRnIB9DM5zHlseqCCHg8uDHE9xP
eXscwGY78sxsfUHvGywYfOqLspUJcdKirqpEap9iYmzLVmqgl85Dy9urgX2y8zOW
HD/ub4dXabeklds0Js4Hc6gk8RoH/xghxWkr/hPRLp02Hokf+7GxxvCMf69yEzhj
xFUGu//1nPY9H3vQSpmmoJOw7v9VrKvdIEaNC1ANIZ1va9zg4EsTMAE09RsOiOnz
Wek0nmiNxast/yoxTL7Q59PNJbPpmlTlit6BCVZ4AaOC1QotEWVmvUOEs/RP48vW
8tO39GP1B7dEl1rjtUUWph9KnwZZteI8bn9vyFC6vIh4CmMz1RWVg95bAknCj6Di
0kMnilULSZNa3DwjOi8N3SKk0lOSet7r+X8keYepm70R3zB1kKMxq341fciDPcTM
FVTRmNk3oPEhVMP3wSNWPyEWd7wkGiDSB8+0CJqFqMFL8jhRDL5F+e+SiKO32nZ5
axmLvpfd1WpHoPAi08WO9mFAZswkJkTfnq3z3lNZobPccLhZucLrkuPqU0Mc483E
W0d9rH/N5/1jIAthhi2HvZ/PdJLWHFHKTIHu6mNdZs4ap1LkfBJLJH5N5dSuRbVI
zyuA3hoZ/P8cnv2bWrXAcWvAf84UkaDnYf9FWz4slnnKgCTC+0S6VzYRERnBf0Qf
3YIH3pU/drOq4kq8QNVf29xzI4Qva5mv9klM4hHK8LH+5MOITM231rXZvfeWMvX9
DRtKC0+4DKfOpr5zqiPMuDvFQB1379uUjCwJSM/4JW/SzNqzg00XhUqpqYBrO/bk
G/a7LJIh4ulVwdv7MdVwAL+K5GgBopDhzwXAEGBSMoa4M2YObekDaeN4EKfHQDGE
xR28OusrlToSo31uWczgRcXgIkhCBoHvS0ooryWRtEwlc11YX7ockUtp3xRWuQDr
e1ySbyHNiy3hJkjPkfayxfLiGTCuAtkvTxRBKbhOwLRa/PSLrBkxZhflowiuK0mW
lW6vM4+RImweq0Uzm0oTAcpqH7eHDm+Vu7C7O6AwKRhFTLewRO67JIC3X/h2ndKb
CbfeTZTtuPk50vOENm3qjC0H6lBKotPaHbxZKTtUcoQDnbwu+KUj11u6xKIETLaC
LMXwgpP08Ybu/hVm5Tmtw6ss2UmYaaF1sM0N+IMqJa4BDJCcIk1lo8iZsi3L5tnQ
9wQwBfeVuB6NW+8a++bh6CAutL3Exv2SfN+lKNNeHQdLTTvre7x2A2OxQmHnHqCZ
qdOvxgl+3IJ/7+xBPFTNXZz3/7micVl2W5dMgyGgpbi0YhbSKeUqMeh1BE+4WBAD
/5pRfu/ircU2/Jih7ePWKmhrk16quQJAQ80YhSDHWN/M0+M7D5j1ChfYNdYJNMs8
uTFp8dloWzTGsTTC6u24n+jvyVNUAKpucZy0UJhqCQJIjrAfEgsvyiZUHiqd+uaR
vsHmPWT9BSbSmvpbMgjH3yMp0Uv8+PaDxItb/f6iLI3gY+kDjZ4oehzPpWA6Hnii
McwuNryBszraczSmMYpXAZezZDHJK6bHC/SD4a3AgBiQdILIMT4kxSjt2Htl3Zrx
uDZRim8nH4F1EpkTM5QFk7MrPzmGis626Zb7kq4x2k//Per7si9HfnImkKx0k/rx
9KnU8hUYfyO1yu2snmvlusDoMNd+7oEoLWbmIEXSP8cSNJGzkaiTLz8lwgwzC8Le
ZdgZ7xkM0MJfNhI7zSofneOprKKgaJ58va2PlPZF3DIRuz9rjZV7AJBlm4kWX3P6
WjteMFe8zavfGk7RO6QoMB2yTXKRBhjfnuMt+dcKrYynTg++oUXshwTBDHrG5DC6
8JmzAwnvMHCjJ8tGm5U8rT+5+ILtMw83hK3p5blml9iFXOAk8qv8CcFUHpI+Zc79
XFko+crdzGZ2km9Fsm7w6sUK6HerT8AYcvDNg7Z1KMc5/FfvZw2eEUlO0BetyGvN
yJDizQeDiGTSJOG0UJ4EGeRBWOtGhogDiOECeUh/IgFqebCNvFRwy3skzL2oht0f
wd+kriig12RoDL0DfdCS6l2hSv35mxV9kzuq+zzTJKMbaMbnl8yipEk5vKmYcJdn
wy0ztKtODe/IxLBE3SeNe33Z8Ak/uh3GLe/X8Dtc1DC794jEVPanbPTsmy8A+o2Q
8tdEwb9aLhsUiFeLDKA/J8GmpblzwvasCEkCALmPprTmJI0o092T8hXJ+FP4s6+L
gmxUIXVu6PGwXasPZ8oKU8So8nT1GF0wQiaJQODSE/9zBzlcioYNGxPcbIm5Aqvg
0jfXu2FZCGSLPq7UmyM0BC4QbWTzeFi1VGbKRS1oIVi2ffa6VmEXvOguCUqS6t/Z
STeevcQbv06i94R75vqw2sB8KKPtYySj7Fv8HLuFGpBvAHGVZ8jrY5lTg/LomNhe
2sl7EiUQy/+kh2kCe6DrctLo9Lba7uxQDGZAoZYqpld3gFk+WiMHf2TQ1E1pHevu
TP1TySDBnFkXIJElYpDr004Xy+zIlqUUx7QkUj+rU45mA1LVZORs83oBo9imMykF
raObnDOR/vqhZG2ujeJYbVE1qvuOdaaLI4kuQvyz3Z7x0XBq01a2jQbFSsNupzHu
nLdQDsV9pQUDaFiIu0Dg8sEzF69deDIzGY8DdGKKsGzW/FxjP++U/hxmilkKZsky
mKV0SUUYipoz+Fb3U9ZmY9HdDjAQ+MtwM9hr8GHCHUQsDQz7RLfM+DuLg/D5jLUH
5coE2f5sxbwIFXtWJYOxn76CjC03fxhKbmH2fPXVfqtl8+IpnHsxizeGwx16XpwD
ENWwR3XLPVp3dDlW62pQtS870j/fX/7XPt6CtVvEHTk9UQ3kTGHCSrQbPOFIhXrc
ePbfOHm49PFZsv4R3rcy0WBbVVm4W2IlUUaufw2XLVxc3AksMH0bKDUe82TvqxJW
eFalgZLl+5WfKsdJ6m4PNXZSRfFysvaEd8P2cnGHAHFWb141zl3KdF1Aqwg2sqJU
Vf3NbY1gYpsLrdrJzmrEOE8iBAxn6PIEgGWHjgYvMH38VZ0aTZr6fxEUkZ2jAgst
iT5mRvtTT6p6uUgxaIINnksnTcZmiUVGUMgxkd7y0G0VBF+zq9GoRKL4TSHsGHGm
T44vM3LHuM/6Xu8ze19fVMVL4ttDVhIeZ4RD5Hkdzft1ris10U9mWqoQsxz2bfev
pFjXu1cNSt14XDTXdcT+CtrDrFDvw8CBonsT0MS3ev0ITgipvKu0r/0LrOVswZ5l
MdHnzTCe4BQaATTkNLt1yDJJv6ZF17Q5kto9qWmLl/cPS+PqwqIkABVDnC1Xi8uA
8RFUCGVlr70mBCvgxU3Ft1/u/Q3v6KDI1shLnMYq49rIjyAkwnb59NkLm0kPqPCY
UcqW7cpLSNSMhCEcJx6tvmE2Hj8uVD3S9LchZg9YCMRCzg6Suf8KU87JL33bKy31
FEY9Zdue2g3TKfx0Wr1EoKkCcUpScVwUfvlPa1I6E0wtTcPRzg1sMY3TLyccT7Ca
RFYYc6wOkdmw613ybIsyWn+2Tn2eC9zKg9S+JcMevOzbI5SjxWPd51UwzSw12YWV
hSlPqqZxp567uIM4DhMUCSVSa8M60acOGHfirGLjWizTvNXoWOj8o0RsXRB1PvFG
MN+Nic0r8BcrT0zX+Zrr00274thmieZBuVzLy2Cy5ddhEadkdAlot9QmaKcmRGA8
g0XHZQTcZHoFUrHOncGRAayk6qXQPvMUdY6Dbbts9QZPSIt6aNfIgRq+xigPbcK3
XDa253WrHGuYNv6fFpk9tL1NNjmRL5LPjuiI+foB/T9mcSdFmmYBe6ZpkDcTC9we
itFeFCGTJg63Gl4r9bNil/Nbk5Hgv392pKi3OQq7o8bPdxo41k7wDguwOHsyMKjL
xpXYcbxy0jST+o8cK2ooz6kJE5p6nrOUS8Vs1RTKQhHy2h/8DGjtMBLAWJLTsrw0
FuMbD+MpQaF2ZAt8Ujl9+i6viaLdtNtUOSU1HBYKMHOnhexaHIr3xv1rNOXJCgo7
Tu+VOthzSxUUMuyng0E0WUciuEW2vz+ELNTFdZiJz/1B/ERTxl4yYtzo+4CpoxUm
Djb++5JYOcATezDPExmqQ9o3/xIONxNiE33jzel0BECEuvXsdpRx9iBkva9Avw4I
3dLvwI3Noo3jjfBNBU+Am+THp+zfKotinuLIsuuXMJCq81ZT6d4/T1oo8/3ejvNU
sKRAn9y4acLCa6RJ8M4SXSnK2n0sAoc74KtjOUZ/1Wm2PXH3x7X/1AKuWk/nbB7L
Xs3yZYQ/lTIN+zUbwW6QuKM9uHJcH7MJJVhwRCZz9cuMqj+NXNKHdKMBKri80RDn
+6WPjRro40RQ3Edd0nEaB2vBxCGZfEOjnNxr+/i+b5r3Nu/QCoQMTO5sTCUaaRbz
eS+MPAJpgNc26DcYxpnhW6T2q/x2dGD+/9uqmj4uKOEVN/9G5xbh/fRtyd24RmxP
LrEUNfvrWFu1rsQdIpayTNuaw/Eq/7Ep0ac8XPid+KCHSe7wMNesItleaJA9fjyN
mmZCera2ECS71ZqJDjIGopzSSoD8z+F3oDnJ+21VrDIL3Gz/KFvHbB0MZgLevXhq
hcXQfvkyuQICRO1QORwb6oNbMGtlgIO3v48YyClrrJKZS7ofYfZGkvihdVjPvHUA
v/otGp1D8L1Mvky1qKJ1ZA6BL7CT4H5So+oUFY2IRJaylKqMqC15QgQCogi46Fu1
fxEexIG9yq4o9xiMUoFXU/mxGip8DOgt92X824daej4+NYRj4A1XOb5gXFEhCbRQ
fKeWx5WrKkSUbhvfgmJVJKlZ7fqD7XB7Q4WyvmNoU5UB/8NHB6MUOaFVozTw3b+0
QYJLcAmCM2tCKRxplgujMmsj3DHCynwdc4duF8TwPAX9lxgBy8rqY2McplvLpBGj
HMkqVHubqXor0o5pQECYGBiu9/rHSBl5xQhhRbV3lidaBr6TgCONAk6/CGZ4M5zz
v933UzX6CpjFV+b9Mw7tHQ7FxsRzPZ4xkkey2dMXJPRTMAgPJ7yWNbEljn9hqkhT
z10BM77BGlVrFpOKte2vInHa2rbfL0TwUMSRTlWhlpFuy7RZ8VM+a6CrO0In+Y2z
OGZwcy7CHkyN7PdMitS1HubhWf2xdwONaWQ1Flq3fECGrLrMX3vRSMAcglYMaZXx
BlO3pGWc81nFPNA+4ZaGkexNvS8KxkBAQ+5/tc0r9aOPp/q0pWBpieXYZsg1OH+3
HuwdKUfT3Hga1MG9SrGMXY84ezncGoVAlvegV8t3cN6VMdwZoRB4gBnvJQif2R5x
sWYWPalQAfVmNzSMMYii71DuZ7cGPmxkMmvfTV3uXSKp81RyGnlW4oP8aujqglVC
P5GapsAGhxPglZMpookNc0no9f25xT3s9r6RInEcE15pH3P6QjasGAsDy5uWGBM/
8rSA+v7yCgAAvxAUCWZmCKzofXXQzjTWQcouHJjws8bOxCO6xu8RRpWgtT/JXkKy
cPSBmDLA0nyr+zDLA2Ftju4eeQBkQSRM4i/Un7Rnvh+EnI6CHfJ+58PpeQDq7fae
P6/jyPiry1mQVKDXZ7VQzvkLT/n2V1O8cyVzePT1XfGJnaTr+36uH8EX1kVoiIka
tplwaY6XDp70at5ynHvkon3rPLTwhgMobHjGtXrGzHe0I+kGImWmklgv1QQhhcNX
Pzr966gw+4BlHFzZYWY54VwE+a1d04BVbod5Mr+PtcJN6Dwkg1vnLvqd6SCiVQWu
/wntnTb1nE+lYOpNPNoVTAZeeQl4giQb9Iuy+xQnX0J2ooqy8G/oKNN9nre7lFQK
JDbSvu5aYOdk9LR02ZJ5C4wi7GTAZcfEgjvj3unM8gVnJOg+Q61qDorDeBe64wO5
drz2NkLJTklX5JzYaXRj2vpDZ6dWq0mulgZDGyWSeHQSZhl6OTJ2nPA1Ols/QrmR
e9Y3PtvSgxoT0jwPvxtuUMXJMpimM5TWMjGVgBUFlE2mfmCWfzBfdKXN8wbnSGVX
C3d8k/26gvwpjR4ke1sDXMLzajW2qnotjRuRFTPMORrzsNvaBJ+gOKlyDsePUH06
xJCCIU2hv/cZU7BUHAfZI9J9noCXrGoMHJy4ExjGD8whIkH9MJ76pHdTivPZ80jr
7wWPS335GvNCH99SAbjNYya3uYp0PPduco+KIlP4h3ocT2l5MT4fGStoTu4SApiE
crE7cRNsxC4FXHzn8zmxMfeH7HdYu2+a8W+OWnaN5Q/mQoN0J5sJ+MfN3qCWQhUP
ZoOQYKrALzszVbvka5lmvBpe+ww7t8b+88xWLM51THqA35V+nqiDg5y+uqgTm9YO
uHl+jmdGbbf9HIqWfLp2qx1pSKzI3ru7N1G49Jcn+VWjhxuheEuVsOjGTIY4snQV
A4FLDp5m4M/760YUhXuR+TB/1zK4ZTUrO07LYb/YKW3JQMuc4gSYfpff+WiIonR+
yGevZXTWVawwt7iuFVVLVbG1xfOfPcS+m7Tp+ffIO+KgyCSegYrM+TSA+90KIBkO
U8qAnsz9jg1r6LQ3ObXd/nV2pJdXtnroBX3CfJmYkDAJxeur28gRScl1QzNJuQ7n
Yb6LwmAkTXtP3gygYG56HeKHVV1VK5pxmhlfTScrpA2J7wOQNU4Bhgr3Qu6G1Vhh
dJoIuikJDosMGvZEIWmLRU1JsJzAqzgQqzT3usvnINF3zLYllb/EA5YfdCNN5bkP
k6rVgXmJK0p7cu+1jDcp+fOLpmltQ5LdNn9AUrinJS089tJEj2zpdXT1bHod56HE
rFmGzfBM1aM9asNXRswXSnlhCNNKgZ1A/ZxL04WbPtADRPvtfzSzCX3w54FteDHZ
X/0iD6OjHEZoPdQSgHq5XB7TKCquUe3l6eFpwxdanagfjzdp2+AuZDYUvCEW7qic
Q/ojKelzHOCh/myIQ2LRfLhzr9jvkLwohwm7aNcfOMYkTFYxVRCx8Hr7yl2VfrEq
PJ1nX7MlSYK/49xOuLK6hjwsHLBkpgGHdKmcXZ9MobPLZrNq2rhtdNwEwxX5k2cd
TlOvbYSWsYFB/D1G/b1jP8WF4TjoWu6LuM4FrQ+AnV0Qj6PEsthssgi1adB1NrLZ
eRV0HMOhF7W5svBZaiG52ZUw3SG/e4mp1uJIrrSk5gcvAuxe1rj9H7fog7trKKjz
n4uQEkXCcCk9Ndq5s0CWowFtd9lNmYxXc3U8pMhlcApIbYi/rpWJTdl6syRWVAb6
5oDL/XiRvT8drIeA6mT8B0S5CosRvBKAVsIRVZqfpVUUA9hjmnUSVe1E9pYAQ9dz
mOfHSI2oHhobFbegeobK2RbtPjc7nxrUSyAhVeMHem2sS6fuT9QhsRz+DxGpXCnV
lyXR6RxlUGARpGh18wgzxB1EbZ+Z3F2PSYoHZp5fboSiAz90GtPvfujVANV4ZYFY
b4VTUrujY33SsVkK0xuP2FNsnUqW+D3+Qfs1rp0cG1uRb5gcBhoDAKaGXm2+LeXL
i1mxO8VioIHoYu9PX2tKqlIWq6hQVKZR4hEFdFFHFx2Rk4g4aDFFKUHvvxJa4y90
R44d136Z3c+oGxk8iPnzaHpO4E+xcIbDkQDdmzZLkQKSYzGIGkY/QQpa+4LOSWS4
a9uVw5V9gBdm2i2K7+Stkf70ySujW1EF76Igg8gimp+dEPYH8PsLOvVXH1xF/WMZ
EJC5hibYLjcB9olA8jok6IcI5ZTruu7lgyjci/S8ak43KU3E7OkKHcAtf/9aM0dy
+bsbcPVRV3dHLVlDfn7X209wSYnWbzqLIp33le3Ui+wZhC3AtnFATBTr2Sink48S
r7X/9yKwTfkfgwTBaC/6oqeHhPANNIZTtghloymwqV+oFrwJp6yIC0qWF3J9gYpK
5kV6DoPkavFI/WSq8BtWzApJ6g1atg4FoJzGnyJ7Uoe87Diu/MTJaUe2i2asq/Og
Z3uGz+uybyQRlwM3DyA9/TQ6zP75AL+x9OpHtAl4ZwP5Jh6tk0kPK/QFquZU57fr
TgdywPD1OhLGCc9S4monoxX2FmKUKyTNv9xv1wPKspDghPCB8QRFNgIKHs1X08up
C2qGD9JAXGzcBERyenDK8yBoSXK3Q3nOb9ShIWb8f/bkKe1q6DYG/OOovnIMs6Uh
S4cxXGeiT+cG/6jB6Nf6iQ0skOGnJNhX36TlLN7Auw0khBVXAHkVO08dxfdw3EwR
oV3CP9pyTJ407NFXqGEHowKMb9hwGIo1GbmsCHad7th133OhNyZSMuv+eFZ1rRh2
jOZqGlfcsI96aLDjXejulLgdr+4Kf25INplz7MpooXj+VSsPlePljpGAYHx3K+2g
DgKsystDb+F7TqHUH8tDePW/Y4Fo9G5m8ypUGXIX9N++kyxFJOTVnbLq0EDTZnDu
6HXEw7L3m415Oc0Ju0foeQZ08ryHCDjbjzHn8o2IOc6aKxInLW5JOwmMSeFlj+cg
ZOKDnSQV/qqIlA9cphcysOa/a35Hd7PDAtVlc0Fcem3ub0JmcrpzWXM0mGEQyMNi
nBiXfWYW+y36A97xCyXaCgm/goEhgxRfVHgor/gzOnppJiWLIgQPSimKQnc8x1wZ
mr+lDutbOmsKxEmG3fBMZkKQe8T6+uzJzcZiGkeLV08gVXAqfPGTpavLh1SGFcdu
+q+iwnb2vL5HJXKmlWMSOP1Um9tsiy6EWlgQC9Vw8jOFbxAAAlsrPRahmVupiXeu
lQdoleTDH2wKkRx1mmXyWtMRaA8S//RxePqCyFV7oiWINzs2TuJHA0D5ajjNw8qw
qqJd5r0jgTuSVkuNjuceVB4vpaCIbAON7ATdA02s/8q+CSbBO8NyD57RefeZwN9l
A7gt8qiYn7s0d9t0UXNFlpYWnIx/VIvPzqXwaJsrEqGhnLQZVnhMly3ywdrQ/A/L
6p7ErPkIfiPPA4yKrct+VThZMGaaa7zZXF9xYsEuUTl8rj7JMYrYu5ZfgcNPCnZI
npWgwxg3FhltQbrlTxVwwS9o2+WXgfCINpuZLzBIs+6FaeYd+NX1Z5SW5+nuxJks
Z9k5eORzDznS2xTj2r6n5eQHuduuqeZJ85A/icRSZcFuFwF4K4KyV6LnnAFL9La4
bWr34OKOIWxqAELNyYqUOlL5743pcAc9bgEv2ntzTOS2YyTIEPEhCdydcXcOXOwT
UNrQy2N1bIfv9w93s0EI6zdrSa9O8UVMSJ9+TbmXg4d4K1nEhML4eX1d1SwtxMiZ
EKg88yak+rMAYBtae1xqWU3OOjQokJH7Dirf1mTHhY7r9XpeH7wtWC3+zveJp88a
0HN+NNfpTbG+XFJgHsnopp0DzGlPh7hHrtF4TrmET6+vh+31Us+JcbtQpwYagO7f
frmAK/wK3lgu1KScQhU/Fuuu9psNXN1bKfkcSnhMNVvU56CCyh3kd7639jHlLuds
nZguKsJWVMp6CRLGkHTj1CIDfpMZlx2vM2kLGl9U5YgnUdcU/9U0c7VkfE2OmKbm
XrZbxqwKU+YEAtr53TCN8SoAsINDHOdJ66xhXbRJWmuHT+GVaHQBjUWNTlLlRlFJ
k8Y/4Lz3+wGTe39ZkWjQNq8rVVXwbgWa4FM4LJPj1QN/rClVURGmUGFHkFuxl3Xr
ujkY9uuscozEJmQPKc2PIiyOgwnMMbV92Svy7Z+FadSbuGdM6F/YFBk51MJ/sCOw
fykutq/gMdhAvf2HwkM2gV0kTBfH86fYkkgRHV6XCd64qDyevnGynIdig0RQ1xYs
cTnpLi5Elw3UqiMsS1+m9XRrdQaQZ7QXu+ptugjAkp0uFdZ9GQQro4xh2I5SBSUL
3QZMSADK++88SCF+CixJbOLT9Cdit2NN5GZtfCO8relfdDWizCs6yiSEZE/xtrDH
gEduv9Yv4TDfABfuaXTRwVUMXD6HIkKBech6yYIojdbduZOKbY4w8MFIV1t1ac0l
dnh7Ov/P4N5BPBbnvj3CmRKfqHD5rnytkJ4hEHkvPQB5XDZB4yudq1aiBEi5f523
VJO0wKqxBP/yDa+ajHItM96oB1x0PHqvphA++OZS3QLF06C6ZDxuXULlU6snsF+G
umGKCA3nvPGs0x3ZcgYsO+MHfVeCOrWxmAw/L+0D4RW01yvr21iMR/oMcaZo0+sV
Nc9H5q31qgfTEz8jXxtn3Ovhdjc/WN91XVTRs3VD9Q6E9w+jEPf6MWw2XKBtD3U1
ZA+zFCvrG050KUyUcKvJbEzWjI4/Fnj7VBgb+xXouqOWSgJJf/h1txJYTr2nDRgF
hv77/CwIxVjHY5PQ2dlGEO8iMKXsLQswwzzzGzJnp9e4l1FWeJIIiqwadwd2/vQq
00f4tq9mKQM5Klodq/DnTsZmt2c16+aKIOAF8BqBKAj4vNzClWdRj7XHSJYWwn7x
PM5ya1An9ROXJnbZ5bVF1ekpUxI9EbbC9wv6fVCKs7oDNRsXgabE5SXLjXBfQUBG
72i+UOpQqU8dq1irJxWkSlXL/pdzYOfIeVYFLjLKCgvDADX2rC99FBwL5yOcAifb
C4j4aHFO7BzxNUJ3S6Yiqf3j0LkqN3HoPG7Wa/obty13ge6r/MD5XrlFDX3FMrVl
BuLKF74yMjOxs+hVko3YcVMlZXtUeW2EIqjgVICFbmbFawzoXAFedtMhllFkbzV5
lHNGNMpVMTYOFo8J7OmX7QzZXgmcv0BXP4qw8mMktzMcWhBKEGwJA4XSMlHfb0PR
c1Q4b/AfRsSN0okHL/3F4TlGGbaA2CzO2u0dgWs2vhOBZn23mNRp7svi4rY0zCG4
i8u6V/gQgufkpsS1/aFV78xQnANKnDP8K0nlK8zIJl6+ednS/QiKuExtR4o/ZnWU
PREpt1F5kYLnXFqPLC9ioXlnFqWP6SUM6LDVLRtUA+3FqgaTievvZcj38+D6VN8U
hhDXHasHoEKAuhfL9CW/UI3UrCwq/GjpI/GIOtm5ZkK9vewFTi9RCo9/VkI0h75q
yQs3qbaG/mxAxdTN6Hfrin9vMnaQgAwyUm16fFmlsy28JxocnUgWU3hJhrKpYQiW
6LSAgXFOSUI08FeQFVNOEbnGq+IsPq/eofFqf7hBKWZDJdPu7wLEDiGb6iXKGnep
DK/Pc5bWZ9qSw4ksu6KwhL2C8xdUwkaszUJBIqwZfQhkSBBNJtg/nSzyaPD9EXCx
Pj0appCrGr0QxVlKXYccNbK8MXw3cUNgGqEqKRYbxWswRsHctXBbMUkrH5F803jd
SLGLmi4zkRJ6/7SWY/u4gFxIpMSX/tS6UZUkGZQpmQUZ7Hzafk+BO/4sHkmbktLd
CRmYIcmgOVevt80ySRKPDzUM2JYf2k6sHXpAvcPhgbxDlnV1gOuFWALpPYoYsLuh
549jOdwCPeWaiz7V4rJcHgDOWm05CAwRPZx3BUb4kuyNZ8nQZVG2L7b1JAw1VwmO
XZ6U267NHtEs1/lsr/pk1cYSn3q1Xes4Th6m3oNM2cAZxko7snwZrFwzRWN2SPnd
Iv2JWjo7sJYbkK/VLrRvO1GKqW/vso9hDAg3dxW0/E3eAOdd6q3cc5QkY3//+X4Q
RhZu2cwKJmZipVFaPRBG7OMcVoUl4XfZcrBh/BOjji4hQqXDqulIPI9YjXhnWUt0
epUPMtSmMhuQrxUz5V5nyLHoJFjMHGqoFUEIs0uauf2Sni9NvkAZgZBlKBorUywp
zrLM9xRJD0T7QQgUen7o/sz+cdemUwQrtKmakaKhCKvkMyJgjoVUrPmeymAHj3dS
zfAZ7nb4nB8wJp3o1tt8KH2hkP67aR4EhA1nk64pj1yqd5DdudHXVcjkyT0gFufO
AET2XdYqxFJ9H2JHZkTgXK4MT5v7aUe08il8HCetOWjMiX8JDWXfksmtC+GsFPCt
qayFfxR2nv/9kn3gA+n3FcmYBBceeKmY5LNvZK18+UoC43jjtBa6I3QGz+Fihnax
XRcYEO8031jAooCs417btNXN/L9xeGjMZzJgwmjtVsy6Huj1NmdGX3WKmT79Yor6
nDl8b+NyMuFFO1CWEtIHJoZ4QKuEF2pdgmswWpHjVFgKsIqpFbnboW9YBhGNmbXV
iCuz0RY2Zb79KdNsUoF8cjhAInp/Jvj81RrCVpH4yM4s9PXjfjJXo/LuNqenQWCm
25oCLSs/e5m/B0uzwu7oofTXpaiqfr4mY2OS9PGHZRVH9KAhBlbeOWQ5swg9DWGp
vAKkTykXjSiSYIb0HUTq5VtPtVbDWHuJ/g/sJkmHKNVeNT5CSpXwCceq2UasTSc+
erVF0Oag5os2ZpBAyCDHXnYr81YM/Ie2AyDP/hYcU6nSIZelg/P5kUAfqa5eS9Dn
XkbcGek+NzxKTK57zkNDu8sMEy0puGVvjr2pq7OCikqamkXywTqt2aeG5ggOYwMS
ChNCpq1QJoLuG5NAqGS8ySuPmolD8lz0GZARYAma5LJYPdMUTUS7BfV8DKgazNAA
HRjE/uKCFVwr86mr73X71liBdvB5+vYikSj1AI8oV6F2KpwZUD5kLtig1CdZ/tan
7FxHewq+N569zdFjPPmjdQBrbrgi6DQD53Vp4+VBAhL73C63n2jTRzAwcJE5GO5R
f+hGeuTQdXxeNvrqqdGothJXgkC+zwOyq/VT+sGU/b5n688dZg7+cFXBc7g5LKfX
nYOr8ZcExxF+48F9NOFjealC3cy7+MYUAT9PN7Z4A7ZuWnBYsvx4FBUBp+tx5q98
9GOGYmCpwh6Fza1runEeiZud/tkwlDCpKgo1/kDnXFIpRokWcj80ARsZuyVoG0NE
qB4buxj/5iGy8SHeTT8ok3+2tbAlipwJPQnbIy637w1rS1RjAMY5GOJC7su6Ko9Z
6HU8+IY5jq7A8eRhtVg6ncVRIScdXX3oH6VymNwqajgx+RB9yAAlJLyHjTQODJ3Z
sVHKKPRkbz0SgRwn8chrv99aE1weMDJlRPzm/LJtDsDEtG0Io69HKSsVdHVW4Q6n
/Lfn6hqRi/eUMbYpsw9/LRX0OaOcAJUeOBwn/WUwScjyHoHD7AOejWB55CQqqYYl
UPqKVG0b+UnZZQV0Dl/7yhL2TUFzuIMO9Dy1mDnj5IPrgiCK+J2Cu+N02HRGpJ/G
wRjSy5RXboGmXDnbK2VU5fo13vJewnQayEkOw2zmN0zXImE6ICyVkfgeCiufEVey
wzvQUc6anrB+aYXqkVopbzPrIqjLWuVqMWou1Wlm1r+nbnGWodPQW0Mjv9Spj3HD
aZCAabf6P94zAyEkAOLMwhFDs3P/JtFKUunrGsWW0YSuZYWd/YDe5tSkuB19gh5f
BpzDrxSG+57VM6NGkFp3+Ng2mgcgt7DeeK1SwauWrVniwVCtcnn9HHwjrYSF975T
+OEcc9grrr7i/JxlawvyzzcG7/cenix5bfnPtBtOnPj0bmDRghIG9QFM7Nj3q0u0
4xR35knEa9s02JjzxeJa5QOLx1MW0OlnCe820ALyatt6Y5ONZnnO8EvxZcNLwjVm
DuFbZ63JVaxAkXBuRFBBxe0XmC6gblpXEu7uHZwqLCW3f8uwnWqxylVLe61iMSwV
2FXpzgl2Og31QgAIyhVJRvwEt+h20DbYh2CDA9CqszheJBAQppnN+HOhraL6aZ+O
u8F+iNiBdPidjoWXBeOTg3wRGiOo9P6TBNia/C9iWt9pZKJcKceq0GYfbpt83CoR
fWjFybw7HfOuZD5HtJOYRZNTKRxrZu52+lLuMjNTv5mngM/sZ4QufEYVt3okHfT+
/N8/B6gDMoCFiwynFnnkzzjQo8LpLzayXfpRTW6l992RnMaMxbiclL8XCwtnO16m
lJSb87Th7ykmqKC9nNWtZ9FDruZqh0/x2TppbmohdYbMNS3Uf4Yyqo51g7R8swjf
2I4Ct7QyH+SWhg59ep+MbqNS20nwwkISasgyThEhHHvJTxLEaaMpFxK/76q9CedS
vkuBJK+6CFvHC6mnsYYf2E2d6feJWKPA1yLTJutRuVgfITBvet/ZEHmsadKIKwu6
fPuW+OJxxEMHEzzDRqA1PBBtfm51tsKweV0pG+aCxhS+ds1A0agdkThLBCBJ+/0c
346YvkptgvBoyzBl9jNk+PllqV+81F/DY6LrfLd92S1sOIfwao5Tp1baUJZbcM9Y
zZbumljmDs679AO9wLRPirTu4cUjBTqc94wVJexTTgXpoKBOWK9CNWoXGYV09usb
gn1A7KtORfN1p51BPE/GkNIjMaOROo11q5r5x7DBeX3900wiFKhscaRq9PePQQsO
mCFfJtE7UVhKxVmjx4OCXJ+sDV3B1zH5pePLq9xCWzT4A+lOzEL0QsxGermllYSC
Ck+QnPHuwi421cANPXosmVEzgWmNf7PfbzWoAC48ddYp01Qye48rQuvzTxjdqlll
5fTGK5fC9ko4hq1FKvSEbwgZ4HA0JpuEKwpIQILubusC21G9MnjxcZn61aXUuqhB
t3q1WEXwefGVajl8d7cTloDSnN8fdK3xDe50kn1wKGiazqoWxYPhjrPPkfkUNEQ2
sRfZZzd6qXpZZhGB6KatYbXbIPOabNl5UJvRaBuNmGNdH5/ERf1s/S3VEinpqQtA
qSx5tU4yAzmmGlucpwKJKr3C0aaSY8qmtxcUIWm6Y6qWthlCmazI3kGYC4f4vwoU
FmOxWjRtL0n8ILPYnR56j9YxgfMnreCyeIq2FpLmalbfg4SjUKXFwsI0mbQjGLji
wiMcJDD4CTavqKd2tjn2PolX3uSJQUSQ/12C+w1kA25b88sYJfn5oEBM9q+deooD
7p3d8oUJLpaG5MFt6YFXc1MK0t0eScZm4hnMkTzL9IawD/br/HluNqGxBi2ORys/
jvFD7dXeVy+s9KZeLBWYXnalRy2AUyaz/PuQ63u7kjJF1oE9zwA+6mMtM7khgllJ
xA4gAfpJwDtMggRGTWUP8O5q6zzCGhNuWVoJh6VTZym+dRnyJxaVlDkIKLjRwyaE
tscS30ylFCTn7pgddAy+0JwAf3ekgPRRFZ96M0JGIbhRkkxFRD1JDAMGygbyDTGw
XHj0ozp854blVQOrdayGW1g/73MKjhEQcSbVt2Ot6MJbdsH9Wz5/j+QGVxQoPkya
5vCydRMUxZXW6ImDoXQIjnahHajOh1a8UIUvEmi6FqYNEgUAgVcPbt2yblXxtVgZ
VdHdpQCdwhYQ6a561wB55AA+Qmjr0szu+IKTVrs9sMUFZ5j6cXoMHv3Oqpli7yvw
w6nqbUhqxKWRhwsqs6xUya1z86wlnFXvDeU9El/Rhl8SqMEE4Eh63N58yLUPl1Cv
r+7vrxpe9mLT30Rm5jIGV3ZmFjweD5Rid6Cn6nye7Sp1lLFZsuzDPY90kusahwfB
5Dyxk6sMVAZgH3Mogrx14KYcBK01At8M4uioyS7xof7fQjiqKMB8zP0BYnu8BFYX
oK7jToZbvdZ5Sxlzmw3+s/FC7Pditf+op4TEjcF3h/96Yskr6olrSOxhsN4BY9Vr
lcwDC/oRe8PDMSqjg6kinXHq/hzYs0O7ZmmebEwk1ZdIy0wV8fzdFTTxbflU6PPv
hP5HYjopxlg//1xBLATXUXJbF6Zwtyv+S7pPI3ODWUbu2A1riXFxPoOjr1wiAxmP
CRtDP6+Xm+MQAZsmGrKhQgDUA1v0JuOyizWYH/SdLZ1L94vRMohmhzo23DPER2YI
/Gj64BRfCg8pf3I7wrrpY4YD5tJOEAIP6f2pxSZK6UGhAnLuc8RV3YIT9bep700i
peUIzSWg34/FFnpwFu4tL3QNMJNEIQpP7F6clIsDvtV4HK6q1ayZBNvpJsHUsZ7k
xv3lTFVTpZ5fZoy/9eQ/2A7jB4UjVt9xQ22AXe991Ry3yn1SXbA6HG3N7WBQNFur
Mz26W1WqqV9ICQIwFlxrCjfrvnG+WZhusd9K7jEGG6KkCOhwv0S1/yKBVD0oL14l
tvTeW3SyCrC73hUrh8QAP82FrVYwZSBEqAUeVXHdJuX+29OunOXCyNuXCCGf2mEN
2pYtL1L0hslWJocV+SBwfo34igcPBorBhTzq6sujjQwsHz46KCE+iOFeK1YG9zk1
/RyHfWJ/PHKzShdLCRB4jGj62fe+XOnb5xa/OvUtyMW7vH1JoGUrGPDQsls8evYf
YJ5bkOahIwAit33rumbraB72YC7Lh6RxsOBPbBAbJxC6368FFykm+4gaMbF59fZ1
3LPpGkPNZoNukCKztIN3suN0w9tGB3GvO8Ql0a81j5p5c6UG9xkxRbe7dacPpuYW
TK5DqYiSc1R3BuIdPhHqtVrprTRbpr7KRE9JSF/UCVclZCvM3X/FWPMiM4xTM4uG
79H1B5O1MxURjj6Jl2Bjh1vABjFZHOXWXFj+CMAUCToltw94bgC6ibEtU2aO40ca
QD91DQrhe3yCh1eFGSel430Hsft3p9hEUvMozlha+PbbhNZPmrCBsA45DAUI4wQH
hzcBjnPc1QcrpGJnawQjk3Z0ZlL6isL5vHeViJitz57cT3rKEHMIisjx4B0I0YNg
IuLPJyKiNeL+a1fL+HFHdQYwDkQ9Pve7NxoLA2zEQ7ye8wcw2ZB/yZgTa3NOiUCV
t68UBBLontUmcWOEsmpv0ZEvAOOXfGe5WWc8q6rQNR7esPRzkQUu+40pddopWEfV
gliy4uk973wOB2eCX6BYPpEzY2NqC7jOEnNhaiVX9mHKgbkGbgY29uPHfH7ouALo
VRajru5ZzigRYEiiTscR2TI9voamuP0e6YaROCaPiihG1vswJMmfG4ockXBW/t2P
x0mbdq9cUwtfmIxuzOAroLJyY6hFvqKvCxEN3SbK53a9Mf3rE7fT0Ro9DQSvaI6c
xNI3RGKFSA/27EnDBEi2yJTwh2LgrmySX0BGQezGPcSHwJFQ+8y/5P2MW7N7zkSI
Hl7yslAyEmPzMDbVQ/+dW6XQ3V9Dtkrre1AvxAhbO8cbfwU39JiY7VZgPgPINzdy
a4xObySRQqAAiRQB5+MJoq2SEANGXPbJH4Iv+sjS8CWdlUDsgx/zjn59IUTVHyDO
lang4w9EKTO5wIV1Vaq3eZzlQmtYtfEkhosec19V81TLlT7TKD8Sd0ea+dqPRQcK
iu6FIsQRXe73cgOmV1XtzVdvH/0YiJuTHTIc3qfV6uL8BSDw3z81l7jxtN4zfrsO
Nk+c8P/R1TlWhAJWiWAYzH2yQk/z9kVXEmpmuwbtHqLnUVxQpFrSi5CXNiqreYod
MryktMZ6wInTEl0/bZ6H2lBXK0N+xcOULewI+ruwHUM0EdL9+qLXe2Wlp1I1l+eC
2yNQfX/yphdhPlZvhlilSy7Qb6DEGl2e5TNGn14QegRw+H5d7Jmq/loFuDMD3z0m
967MI8FWimcEW9zjyImnYeBiNhlQeWIoHk+fy6HE8w3Xm8I4VOSuSVqbM/+gAb7w
3fcvDhhdnzbeokYE6RgBUNWBG1A2gFdjMT4j2DbJB/0UW2Xv9kL+jBcaNaATjB8J
lwtQmpVQ4v8y7K1Cb51y8ImF0JSDBFp51eTYjiA/aGhuE+CQegNfMB13wAc02p4H
ZIX27Z79w3RfLdFSnZYaJGPpMp3Hh8hcDcM0CEYdANJ6odA9m7T9y+KJoXuPo0x7
YfOIy7ibjBNlAPjVM6DdwTyfxfpcZ4Hb+E3l/oau3d5A8aE0wSw8iYUfXrlg1Q3Q
m/iB8R3Csbgz4DIj+kjUgN/2uVVwTmaEtqhEga59sCPP2B4JVaQDvQGftyDDg8ke
i0RvgTHrHZT1H7EWmul8BiSCn63MJXArPxIPn+Blf3dSp6dU3sFijc3nIshkvvnC
8FDZS57PWkdlVZ3CqtqtG3PmeQAiWc4MpIrxkIa2V9nc5I6JoamrJgFli2gwhHYQ
wHjUQYSNgz7tbWwUDVNsa+06CAR1pkjbuKeMD1/rnkVIAL8j3dJM0Ve8X0N2wGsY
22wwO5Bg8Jhr0i+vjZ9G7fbVK62nsQEd9AMgbHtax1QENu10WhNictITaqVG5Ycv
kVtOg9gbh2jBRubrfe/y+/O421NMqiBcL2L2iptWtK7NUKfjzfDtXpqGk/A+7xKs
Ar1rITy9GlAHffhPQNn1ANZYkZSM3PWek8LkRAty0MSQLM3xO/iJrJlnxu4SpsOv
RiDWnmskfPyRvb3ydHUW7IbQSbVaayak2dRLam9br3/lQ1wAypvDjxVXya2QWsqh
2g9vX5b0sDiuxumdRJFcAffcnWnWQdkOqHVnlRDWGVOfQNvNI+DJmvHYsa0r5FW6
c1Y4MrXnRwQXWqBZVs2hel6UR7jvAGXdj4QQo/DIMD/CtxECC6wCyx4q74ibJbxq
FiSyzR5L3jwJgQ4PNb76hfvPvD50rBzL6ISYaQDCn+ZyDeWQ30GxRpt+PuaYu9rg
P/tNXW3Z3GJXoy4MCf0IjZcokzcRGETImS2d7sX404oyrvdJvcbPV+N/xNuByZbe
LWWlTqNRcuYnRlDt+gRP1vXgVmPisFHQ0swtFicbb7/vdnFINrQgW6NEwvk+ToVN
4/E5BP1ymbzYq0h06D5fB3fUouhUxmrqm+FCd9V6uFNOk9ysa6WgX/87ZZN2R8Kk
s6t3fCuMrfimr0bDaqXmSU/WzfN+fOtSxb0I02GbRRPT5IoqUPbXA4HyOnvK7yqP
WG5yPcd9k6sM28p5OkMQi3bUs6fhmm96Zy83sd5oysv8Pfhz9vwThmYQfH53NUBw
EQTqJQ97i/S9hsCSXsSyotflKhjYbNXILwR+RHUHdoM8peFns3nPXsu7MGcijLhu
OBjgMRrKzK37m7K4qwQDAsZGyWBMswuGP3pk/t3OZCr+4dQgjl/1BEeuCAowb5DO
i12NO/5HzekTy+QLQLX302SdTGONIclfGvD++/4hfbiqThWHhqXgeFHZajmS7k7S
TDzg4jueYMcjOlCpQE32IgrrP/mjS5Cm8aFkmnpx9opzWHFB4iLcrj6+vMquIch/
p9pHI6dEkV7v8ainJifrpm59mn+fitP4/ucJM9vMRlaQAKitxlkaQwsRTUC51u1y
D6+1SmvhqVqfZ+GNiLsUVkJRsRh/jLT66nrxwh1gcVPrRQ9uYqilBR+3KRMn69JP
qyBk0GLWXzZv41+PZQDhNqk7lOJQOeMLepJqpqGojpfxHs5vqwQbQEyFb+HLVXyd
UQelw3/Lsu39i3MiuVG0agOSF/D0r61aIZ0uzkXXzLQCARZYl+zhoHwqU6hF29bp
DrZlvWay4d8lji5F1YIkipoLjIkeEQHcuVFjrcwucQT6xf7dg0zEH+S+s/D94i5a
oKUEVYIo/Mt4zs4XH8CQWgQKWXrnz+H2cXwBvW6tMF3mk/xIGwGjxgWQizfv8b+9
eXvct++n+SJDNlkP0BDDBV4gONPkudMPIy+W/2fk/0+Yb9oCg4J0StmOWDoqnrgZ
xYY9owUmN0kzJxw8oO0kOo06hn3Z3OARZBasE80k6VsTHYkxu/m860bAdxHbZd2F
dNSVmJ3TQkXDM/VDrsD/e34LNg54Y0tL+Yr/sOft9zIoD4oPkO4W7L3nT25+aq5z
ynsXf3eCwofdQPU7+bflZdv82x8QhNFMIbHFFtoRPrGmSLmDrximZGvnmiY2kTXF
bASdZCOaRIbuTvzlU26YtfmtPJvJ0Z6xnxEjuc/4QgmR1i/mmeZJ14ukUwIj5l1Z
rBWSfhv5+yOm2rYTATGyi7Wi2SjR0wMn/Ia2z3JtpICW+lbmkgrH87QtFhtZno+c
Ytr4fL6hZWiuoyfnrPcipOVfAYCtMI3ZfdA0zZ/7qdbHE2lgIogk0Hn1wJTyNYag
1vSMXn1Vlzc6jH64FL6LJZDb7laCKgQpSyLG2moHgTEcaWX3RbRVQXoL2atopyjr
1/0TRfYeTNki8Ffa22GRZV52xyYZUTrcCWvhKJtE1qnPRfVo7TQ4cFFGozVsizWJ
4fUnKm0pAnq8JX2dInsW7jMNjTpf1WJLW7ZC/o6faWiWg8MVRpW/bAGRxH1UG2iK
ZsfFYEWwCnAcLEh9r0kv9Ws/Mhhnz0R3rltspNW3aqN57YYIykhv2aoHCfYKBAbn
+UHUzZ7YRkNsClE7aoFg/N0/u73/Dciy596HvfZT5Tx28Ug5Y9K5HzHt4j57E91y
avmHQlPN7WU3ziveiBQif0+FmcM0P0EBwiY52j4xJcfsPmv4cAQxwZlrcHY8aMDO
vFll2/bRbX7Ho3zUNc70g5Ytq7vGiGbkPOo9myVr5yJZhqJCQ+NgvE57mFhSubpp
c/JO9df7z93s6c6LX9kXkfAMimGve10dw8LVmfxzE8yPTzyRQ9E6MXykht12YPfU
Az3W7sDB4hD2X3kKF41QNFyMtoFBpRV8mqAodQF8EF/U8e+GFr1/CfaEM+M5R6Zg
pnyB6RVrQKzou02FxYSByNmYzNBn/kwgNd8TiZpPOYI9YXBg5EVNVYxUjPHQtb0E
LbOrpIlsbO7xPJHVjokOnjZSStHWS+XutQ8G11f1YfF6HZgs4ZavfyTBuI5+1QZf
GkLT+0+lgL2e0GRt7GHEho6ORg9Qk8QkaKqwPRhMDJXxqTO4valI4m2gvBLg2ndF
k4npSC7oEzCLpNpbm1XLuBy9XiJ7CLktGYVvowCeQPdrxnqwialg0B2NW+qtywcJ
LjZ9PjHHZxp+XUAC5h7x82iRg2ttxGQ4D747PyFpH/P5Xm9I8mkqpT3P9Jn0fMGP
2mZdYjomtbL4T8n/s6cuDjgOAFDLcy94Ng5RACGf40opkVF3BaA2Vkuwky6J5gFJ
QDCpbYG/+yrYPn06TBzlXcgrKa/w2nKPCYWw9LwuSjDXxfykjqrmyMDN1AP5NEJc
MN7CLXJL8a8m8TN6PdI7YD7m/+SVA0aUZQsfQAtlIyi8sW1+DTJht7pHMlWQn9Ec
w9CV6XegyQ+4ktuoggMwMeMhGjnBxGpvTsu47ksgte2e+yxyOWX7SElqH5/Acoi8
lhOQZ5FqbHv7jfHar5w9oyFPejClvcrqaoZ//MJJHc7YrHgcGy3I7zGSlUFWulaA
2cDDn967xefgfpP2qOc0tJ3W2LGwamzgTF/1Q4k3KAAVMcQuyx7DFqi9uPDxh/G8
C8orDZ8r2YsanZkGgFCN0smQ62l65AwXVht+OhbBuD4smkxErtBJceqMdSHrQ/Ba
/uqAmrapYHGXTmDgPwRRrG0roQABnrYY+3+iyAjpuxOjgy+BGA8yfepcXhssWcuw
JJKLaZPHvtL6b9Qs1uavO+8lj5BhmPl+fS2lYjFJMvjpyJP8Q9gZsYOEZXGfCUl6
NnGkbwyXtQh7gV6onELqOHIysYu6D4VjBrEtma/ioURlz27j67+3Zpn1JmyJ9wrx
HHFGnbeKZvB3+2tfYQiQNW68EGn28v0JjvTo8S0ypD3e5VrMMbdZSHS6d7u/GwS5
fa0J2CfvsPg/HTl2hU6Xb54H//J01rENX/gCrmoL8YT5x39v9je0UL7MYI1OdCN/
iKzPjOn9bVlxymshhw9HUtDov/Dm8T5Tn1WF2CZT8G3FYgGA9SrTxbmuMk5Xfi1V
JpsrP8yV3cZ6qkEq9zamwiKTyXr0Aopm47AJK++2sik7fPH0LzQBrTNMH6aOr+/x
Vdpv46Ei6El8centuHAyHHMezoE2Zs8W9HoXw3ILW8PLh4vhg5znfVHvVNf7dTs5
aUHf0W6uOtofddmqpqGYvgQN0oopiQS3xX5Tbx7y2cdY0S50ah1RflrIbRb6c2Oj
c4HQiF3qNIs5QSoxovHMZ9clh7WTaSnkqYVdREusM6eFHirrL1jE5QFcztAHKZVK
0/kIF4u6x4hKbam94rLQwoew6HkNnPw7WCy30i7oEw7qkoF1R2gwdELdfKjxRySk
ckqcuTOXvRtBkn3/kBKThMe4jWVj3WAMib6Cy0ZEePeAlaOA++nwYJaCLloAbnSV
WyqJoQjOmKnq6UnhsXRhpEC9LjFaJMOPCyv3KYb0G01e9UW8d7xlRM0RH3vhke8F
geuwuihBM6AByKz+L/TYC+Yvd7eq+0VTdHNuxwQLSUWGrpo7W3SsEx3u6D/5bY5o
NuKtuLSsfzybbmJGAHvAT5GCoB7FpNw3qMaYBROWfmdymhmXdOxyQ5a4b0tDsjDH
av8Al62jG1FDZXjXAAIF4ELFDprNEg8JNUZbfcmbIOpNuHIVHN3Jph0HXT9Z2vvu
U3q5BE3cLoN0/2NxAmHt7QjiQVnFwJ0JmtFRJ5AjrZSyZaQCspjh24T+yGhda55Z
u41bgXqg5JU7lpRWRTx+Ll1zyyzfQc8P4Fh+7N0tTyKmDnNj3MjtgxCX2oRgU2ub
YZSCoMTANVoLYUo1qKvSDsUVJeLjOKVJ0p31G0A995vpHuF/zyx4HWNthlzReD64
tuNozI373mAIU2DTIR4nErhK7EVaBU976SUJuJgwZQBh8IFlAdNRt+cm7UkEj69P
SqT0bkx4gRmpqcKpJn8NRCA/RNFrxVJL/Te0HVDiuBSYHiVIvmAHgmqhgPQRftxK
P3eJB0RLRuKZBI08OStoz6Eyv9XmgDdlF9UCkSkTeeKOn+VTINxwvYaOrCCfGcWm
Nto1TdGfbS+9VzqjcmvloF5CPDcXXF5v1NTt4UqPd+7ejLRNoNpy7OtV3HDEBLnX
DT9fpVaPhmu3OB4ZZnt/6005DGbJOFqpLelh9SACSYDUGySv+yTsqBj+ecZPJ7f0
NULsfRgv0Y+r9PWzZ36ZQuzR6GY2Jg3qICg+nwGW7PYVOkTNGQqU2/U3qD6rjsdI
UMpFOhVB5CV+r+Am/Gm/mF9ZxTkr2edUHv1jbqgb9FtDUKge6j7pNu2oSUlUhUtI
5zLhmiDAUcO3MIqQFjcjw0P4OsCr2o2c4Oeb24aNa3Twlu1AatC6bI37M4DE8zcu
p7hfBw20vWqf5kdXACWxN4QnzNx/xb1drVpBNVtyOJYK3HQnQGcmrxw2teB9R8nJ
t5fwWhFn4Okm45XSQCmRGI1KHgTHimNe+j+YbscQ+TTnjKwsMvJ0DlXLH95luf/9
Yk4+Mh37OT650uwsu4vH6ygPCdjutWyaGCpqehS7SnVsQqEOPU64OgFmqwK8lZsX
iwZOZiipPHX2Yx9c8+Y0PMAxRwB5UKvxS4Ka18b1HjDR8xjSzF+tYtgURrT57FJl
rfu5ElAEqEdSxclgQqB3L43VyMFwaSufWlReqMo1dCnx8Ez1SIEv/Awe1T9PQ2c0
tUFPJaEoneNxAg2MAatZsrNaBn1hQ/bK9bWjvAjPiu7A7FixH6fHfcYnL74a+o8S
cr2QNICwm4X1EK4QhABPvyp8z1taI8DgGr4L7+N8T+agV1GD0e9L6BceiWiCJUTq
sLQeE6Ia4U9X2PZkJGNCqGTWe2uxVsgwqgZo0VyBq2IEFSSoVphJZBHqeBnPzNjQ
0SMzm+cLmq1DX5XZwEN564fyacfLu3IRLm1+OwC5EEcK3Cw1x+UxKMK9tMNxVqVg
Ea4miXMOVjoeU5WNAegM0ZpwnENmPSexic0goTlavsFXoFLkplkoV+5vjWoeJW+J
JRxklUJQ2IOLsGuoo4ZIpzhEOzYDZ55Ju/0hi4iVF87MJYSOtl00KP6cABVeiUzf
VL7xU2OBDxdUCkLVXSt5ymJ38qwKuKyR/yV5XZ1BJPtUDIJ1FIEkC3bFaQQnZka7
EZApjEfFiGuBp38WLf1c1ORozE6iepELW31Mp0zw6iC9G9gDmfrOnw7wwh3b+gxQ
HbnHf5erDmqbtiMCcqX97+wOZ18AqBSXZz5oEVAhLJ/d90W0pT7C6UtoVjxw4z4r
y4XlmY0A7zXKQQ0C6A+hfKiMI51TP2SPDDqYuUkTdqEOrX4v4J9em53wEQlz7dc5
zI130S6l61DiC8o3a+ayrTA47KOcy6O94fl8vW3j/XBS/jZI8p7zHoTtXdGmI1vD
fMXDmmukLiBkXZPY+NLFCGqVIj22jc6AthROv0FSAfAVpadebEtwtpkAmzv96z3T
Y056k5HOyZhk9mvt0M3BhOwKIfYEzt8DeQM6MOEDI74wuva8Vfa1PjCLMCuU8SeO
wN4xJQwA5Si9gSzvS6Bo6E9tLBqgnf7m0z5zycAvORUtATD4PrXc0Skc1S9kAY3r
lhGe/CqCLYEmxeum2KafjXXnmbe6omS15x15Hg6up+4Bffioi/KSbMIaiPfKTHTP
VMNqQKuJpoOOuBjZbQs1SyUB0bbdpRB8UXNZoUHCCzm5e1DA0F4IhRD6T1IVlWRx
9CTmIxvl2nY73CRQRND31mTgj+P17uAluJ24CoDNBhyTBnILlgRNm5L0stnMU9hJ
meXhh2a8BqZ33yw5U5Eci0kArjWWUMaUVlyDfYnhiYR9EJtUk7vD8MQp2KNxHBHX
/z857/Uq2+DFjU+dlze/1V1BEQywm5FJ7Dm4RoBkV0cuMUemDhqBeRxMJqb2Cm76
waglpkXTVuu/Z6NMnWZYseTZCIi2TE2fmZAsc4SvkMden4cjyVmb2LosngkeWlJs
SORtRrHJULKyiybEA2yIMxpFktKZI73Gu1iSAM5thCmJak2n+zpHBz884DSld3u3
v+w+L5qBK4cR5o/uHKODOmh6Y1J+ZRN0D7bg7/EsMpK+EUmwiH/xPmbC6x3t02EK
yCD+3NqCZJ5BtFsHS9cpkA+h81S3qOFTaafbNqO0756/LR9XAC0VLV4qehdNIRsm
0zPY+0yFmE1atxQqBiTObYCLVUb7UftM13xtwSpNw+kKgDV+SoF5LGtXGH2Wyg5U
ENrC1Zprl63mB7A/7kxqyivvipfCCE5OQq+gAu2Q68z8/p8hdNsWoOU/LY0UETu5
eV26+ZGjcIxQJzqwzx2dwbBXU23A7Kht6JIcXoTGQjfUwrSwy+rr6diD9+dMDg7U
8dVtTPlYCSK0AZDb7emsbLXNDTKvXa4ob82+EPrRrckLjwKKCE2oTd1KfuRA3IGc
ZNxPzVCq0oGPJcO2VAIEkcrEGFezjIHNYiQXbY100fFIR9C2EL4z9PCCrVoi9qQV
om6mCEyVs8N0pVozU15bLH0CaHY/QP2BSsmAiEF8wOJ7cXV10RE+lCAm/hRxeHkW
Tox/ShHnA5gbjOrxTSJ7gqDZPq8gmQm9V0l/B+yRaXZgYbId6aQQKO6EZRHlCJ7S
NR5zZ/xJEUJnXZPz8nj+cpfinDR7PCNfSYGz1pdtIw3ViLbZzKO6sCbS1zd9r+h+
+P/0+caSyKo8k4SyMoThkQoFwyGMBJal/1tLc4HpdTFOob9sosA/GBphi6smNWL5
TQEbtw4LCbI/zPknIQOOj/tioHTf0sxgldRRunZol8o1+2JUqdScFn2VA2lnlF7q
wmMSVOMauXlxKMNlpI9Q//U4KHsJScJc7i7FFYviyLzazjIwWlSfumdCtGDlqov0
RbEe+KiAJZptx+rDcrPaNFjzDUVJr0DqZu2LWpuAY0RA9Adr78KKyIokpIeuD9FC
BvwquLiSEKyTm5zM/s4qYmg6e5eUzM2QBAS6EMFHKQOkaPaO91KTNBG+pD6Qmn7Q
n+HXm2Th/X8HQY0UEkowfwRFhkg5FVJLxnWbqvWjBsc2EQtWuwvW9hv9rKcTElVE
8VpTwhuSTUsiccCLqRERI+NzpZos0XbI6QzhOJQAIYMJyQle+czLj67ecWzexvmV
FLD1BcWYAezuixPleUM9nXIs8uaJdCakvhY7uR8JSdxXzLj6Ex7+D0k0GaTOaEe3
SMcCJZ6kegQKB1s2OWSYs/d0BYdIwdZ4cLlmOLkDEoNnf14LVwBqxnJGDDZW9dr0
waRL6j8L0UYBiX13goLPVtzvJXGmd4lion2lGfAdDtAbBG8Olhsmsf0t5EVXoF/q
CuKFc8ymfHoJr2J0IO7wENNRYxcX/AxufG9fZIdBSXyBCf/fK6n1IGp2fDz+290L
C3oEF0Nqb+odzfclnRS0YnnozbD2MpQBPzKzCfkO7d7h672I/FGZWt5Pe7Gl9lqS
XM4xnHvDH4y+9Af1g2467DpbWqEz/dJZEQZHQlMWD8gbNiZd/1TkeejMgnJ2mzeN
PISFK0BNk00Kj16aPJ10Zr0vYrl3Vgm13PnCScYznXQM3y0tHwJsQEkVnn+x+4Ea
pkumVZk1ZYfGlvGvMgdhHwopIRTD0Qrj3sIWiVtf96MJNVdBrwL7atepJMzdX5FT
2qcG5YNfwMoIbG6e0Jqd2JeqnfxP4xuQSF1tZzxE4EsBKhBt2XEKVl7e5QzX5sXB
4r9rFFVit9gbz5E20HNxXwv58o3/vhRWgzIH8csXqOFAt37UwQunrDH3e8c45iCP
xXRPzLnrIwPeqVpq33/9GpVY+aQWsglXzZlOUbaZO4oEPA/7y+hlv5KU2DjOWi5s
CRz3xWUmID+cNikL7WXt01FS8LPcWERujJokNngdsIATfiuNMU3IU8rbldnEYRzY
GMWny0L8KyvJQNSaotTX4Zux2EiVtoua0YTCNZN9Bjp59zC25oyt6k6KRvVCaUIu
Ze6WM5WGx5gva9kbBu3XDer6lp2uDoFPvW1fF+HtHvScRhQuDf80Wzf9bioz0DL3
PvcCMfgCP7CQ1P9lqynaYFFyMBiADCIQAnIO4ARGTqA/zV70hZcjG8rpx0boJi5P
biPs8PlXsCeM05HFlT+3+qPVHwhQTN06gLake9+Qd+encLTSVMU4MbGOLRVfBOIK
TF8EoZ9u3SnnklYCrqVziXGwG2v8d+0eAdMHDMa68d33RVppY3zIdgTAr3SIVLCm
W3BdwovGCd1b8lZAhPZG7WZLU2SaiOUoZmvMJ8SElkW++KN8Lu+0IEcajteQDiqT
NcpXWaYdr8zp3IQFOdodk5InssfCZw+gy7xK+PgphTd7PhkkOguir4Gt03G1wQdX
PL9t60LEe28uDzmm15UNPw2nFVg2JUtF6hOsNLLpqaqVnymrfC26lJQj5UOclIwj
hRMtG4i6N576I4aVHpXfGA2uybuD52Ibscz8UzjuCk3tktwpePfP+WdorAyZpmzj
AxNKvhurJvrUF3QwjMgbfMNQZbCc+tIVowhglkYOohLsN1BYArIvB+yE0Z7pzCaf
7S7eSqM8Pa31SJbEx8KTkWIfgR22OUKF8Y31yQrwK1IjyIUVeYgJz7BsydoH9NF8
dn4GQWSfTe1H0GdM7v/jh0bGX+fHyMrW8Kixuh77dKY8Oc1mDlwrk7uyUhS87m8A
sd5MPkwpYIlpLd8FbBo+Japy7I55WtOnhQvUxr6YgTzG62LtgFpRH9bUFLWr/pgL
tT8OxG+m2rytK+Pkj8sNuu44uA/UPEtnzEz91z6XE0dUad3GHTkChuwsmqOPMvM7
4QJpcRcivcjwG7g/1O2stBU6sxmLq5VaegwKBWn1orQpfOfB2vQC1iPsyeG/Dk5n
0P8Cz/vMtP+5tcdsuGRGNCusXtV6QFHwqiqPOnz2R8D1aPqLZnrnpkhY0plu+Pru
c+xXZF7iY6D8+W3BgFGwIZPxoujgYWiKZ+O3o4MgMu9skU3Hv+oMXJepgYc0VBO+
yfUvxe+jv0Z2K8q+ymMRoWuMeFuoxfa/o0gJ/orhRr0C4581zK6+nKAj599xBFgD
VMecYKA+1/39BPsO+qoFHCdJuhhdGtYvWTAFG2XJXAxKIe2u8gyG7i67JJJ5MKlW
ZdiLf9/IIrXdFI9JKe41nYcp93zw3cqKzq178geaRybs2RDdCLdaL0Deb+miSjzy
d1azhZqCnt0s7imvF6vjobbL8j4jXpUG2VZ2WgXqfioBKIaadzTH9wmrCmfSsNS5
T5RLW0OQQDU74dum2Crzs1gE+I8QaTgkGB55NgSktc3oFSEQUmbhXh83Ekj/OSLJ
jNW5IPqSKD8fFqzG+34NuRuqYnVuXaG4iHMmGRT8Pn8UZH35k5l0xK53xs2AUKb/
wj59Cw3JD+H98lsVRljK3xkM235tyUzyjq3DGIdgL49N4GLdzDPr+tPYEpPyjr4A
SddDOCqa6EQnD6Fkbhqt/mWE2QivcHGCEcW4DBQoRU9OBiSB8fomduA6kWPkI171
/TDf0jq94fsrXEvMIZWeT0HEhWphAKCX+mOPb+m0hwhGuozAT56f+vIJf/pYgqqs
5lTXmb3fljMTdcZDtqHVUoeMFWOE/0Vy5hnxzBH7xZI+5rCNlJD9CxnhYuW5T2Rw
T0tdTQ/YQq8LgRRcfA4Pj3Pk8jnIbtu1LD8pXnxlEfpTCp9qOqo9W9YOQPxB/Tcm
p++Lr6G+hooWAgJN6772v2c6hMnMK1KqYiS44wt4aroBJhn03ADgdhU2o5DGagzR
rVqv7WvVbcPDYPvbgR4aykomu4VjPWyniwqSO86hJl0gnsfZWXuSb3jwxUI6zOFT
/w2c3dQ5RhBxPTghHllHOjwxiDdnh2Q3GJUN5IWsfGwqSQDqQSkcZTd1DIZy+5Pu
BIHnCmcLY7/C4YdjnStQY1/RONSEQSSfZfHRAFG8QlRqxJ3kNMRTkrj6fc13dGtR
bqhHkz6WrWCY09r/3cyZWN9mrHWVsuJGe6TdjZBYGD+7bw6ZLmzGjWNjoFeZrEbT
T4PR5opt/MIAkedBklaC7pF3emAkoUskHpi1k4gr0DwTr6ZsYTbzlNqYPHE12sjU
IF8Isi0Ba1x51LI9ohp0wEMXsDIgjTsiH14aYb/LzTWTqUacxdFBON+VgKWaXX8l
rdWeZIM5UhDoyW+Vr8sZKibaVUCERg9l1eU4bL0N8NDD3/RJsX4rPPUCynxEQl0E
9u3Rb/aMUhY1daXShCgg06Ky2WbeIdBKASU16proxhg5LSYVczCT6AyXQPg7KlGl
IOvQrMMV3fPREztcxPa4nB5dIaYZ4dnV1PzwtT85O0leblitSCGasDpOa38DVCFv
PVApFJz/2Hv5BBvqnjK2OvBmMZcbAuToggALFljdlE81gvqHoBdl/sA+vOcvust0
alJiRk3zGhrXbcUiKufK+RzYHqXh7pZ1oHwtGpeuwxbFf3GDqcWntE4ABaksLWyE
H1zMl8b2XrSHAci2qL3zMhKmxa8oqCRa83664XgqFTK4PJeXzYzDi1imyPQa6JEG
FcJi+flhPZmAfAB9W8U+YNXqkTWUvTH3NmWXfyVd0vVbNbc5gKvM8yz/FOJgbeDb
KtzRoz5kL2uawqSu1mo0Jw8SWGTxrMwIyBjrIa/tVVIKCrtnS8o3GQR4Z+26UK5k
XX89pWTn7lsaiQY48LvGVqSIkkRHr5nIlPyoXgNz2TE2WfFmWp3OOEMbWg3ohu3d
yA5PWGFC+9cvnR3PAuqb/66VOwWODslK6r5qJib5J04nZ+J9zfdeBSuSKMT3YQra
IMYpHDqz5ChALcPfh9azGEN7/5TnrNmJe6y8gaLHbUjuMgxuBrzpsDM3mtCVuZ6N
gLLftymbhwjFw+huayrKV9prGQLdDE6yBTfWoDcRY76b0PeLFK5ivAfz8YJLmDNq
KoyRN4YU0hSLPd3r29wDFV0KDoybpJAYbps5aHQ4FBLoH/d6CphjHEwGdUdI+0jM
49VfVMv5rApC77Vi1qERJEywCr30tAmVTWsXOHyRGAfum59DGzkqFoqg5uAgdpi4
SLx2Y5XqW+FTA9SjyE0MhEO1dNJGqzx8EgTyBjtIQR1VynZEGIwjCRhBMlpNRKxb
LEkusOlA+anE1xPIsBu9DrkCPo55RVnIf/Y56ojLKRyUs9uZPYgonPPONGbgIxv8
SIovTr0GoGzrA0utzuRffB8QNdzWXem8+RNJ/tS4KZb1sIzuylLsoOlCnBp/uR6x
FgPWE+S7RFyXKcvILUpEwCpFGef0i+uqZtCkVY7PKdpfYo/6UfnwH+IAhd4YrA/Y
afSjI/EZ7KphOBmHArwWPSEM8mktK5eMIwZZ0EkTQt2mNYK9iBZPnoTsRUdpW6WF
xvX72Ygj/nYEUipxbdm7EvdDecYZbDxbMdoyY1hLk1oh3YToSeNod8LYLbetqdON
CF+akflXaJ8qSLpajB1cwGYw0PGH3Kms43Nwy1U3vHD3y3MYtNkGZc4uyP9Z097V
xiclKyTTrOz4k65v9JH8BcUUe6p6CLxZqhZVPu0yS/M+68MgJ4nizAaYGJsbtfcr
CEyrumQRmCKkOGS00eQqTmppwWvBGyzSdcQg3x7PXDLTbenKqf4sYO6v0VElr+yo
vTncat5MWejguOlU8mvmj+yPA4j5nXzMPUHBr8+rohfOTFr5uzlU40CPK75EkGuE
Zpm6j2XwQRdC/GtydB3nAcsGtLEOfzLviADsdtGo5sY/YpfdluCOUWe3tFujzmf6
wP3/7FSV+tRa5dZ1hX5QoKX9pplH+DMWOIuy0N/B8JtyW80LzuePWVpd3CYw8/YX
Fzdy2jpyvEaz/bb8EF/Ev8cRxabnHU+o7r+vy31raYrYVJfOqLL0jOKrJ1LdmSc8
vCe3hmnmJ+lquzcgrJhAD4PHqBfTEGLXda3OEQ2Niq739KJ/HRnbmTk20szb2OAU
WxCLbkhNsMGMNCK+6D9Y2ajw1T6WwAlgM/WioT1nLZefueFKPejT0wamTpBgWNEi
qLt1xWkRABN/c+RFNv30rd1ByX+fnOEU8Cgp8vYrjzvQnKTISKTHbYA6Jg5sVc/q
RNtckWLUPJ+Q55N5rQQmXRVocBVzZfAe66rgc5/DjA3vEKEhdV/QK7OmO7LDbs/g
ks7+hhlcAj4bIWsIHRWFriIJ9r+FYolReShx2VWeOTeBjdXLKfLOym3nDFMSDKuO
OKgZ4zwTlk2kqiy7QcOVpJUQXbdyoECTNA6PtS6tC8mFhnsteoiXzgMRy5OQO4z2
frBthmcNpb5sP2Aiyx6xiLoA8lbOgyAdXE7X6FHlXMAz5/5g+LP7IbzmsH+xSJ9X
m8GbdsDr9fW7QA2dgkqvSacRb7qdENl1U2OkXIEleWchmoABBhkZdtjIvorJbm0k
fzbML7rieTQFKuFaQPFFQKs0aTZRJafL/uDn2wcPOh0ztHdQQqE2fGdQ4xwgyeYM
ZpGuSRqCKa5x32UxOcXmV7ymgKRIBxVN8HqaW2D69qa36odxmFooi9l15ADd910r
EuwybWtrcg7mu7L7K9f1DhfB0YU8vLfK99tiXGzazAeNqYQh/v+5VM/pRUjrIiPT
PhkvHCbVHxj+dyDYVyU3biXEz0h/rJNleFnCdmt9PA0Y3VLjSIOI+gfaL0AzcJ2M
4Mwe7Ks2urus5nv06txIb2irTAMcy3Yy9JPt3psJswm+wEL8lrwwvI6km7rGUP6y
8Y7ysovW1BTkDkMmF5ldtcFQABkszsZk+jTZwxRjzUHP9s1yprdBCAPni4W0Op4R
l8t6w4jdEAOCvVJfa9LFDuH3pckVRsyr5NvI/FUeyUye6GcU8Bq4jB8sk5ICCw+p
8XvsDVrtfO4sqJDyy8bATXmC36bc9kYdkoYbT4IUUngSu4wyJP/Yw4Tu1NCbamUO
b86LpOK+c0u5RmyplGmSA7rW/5b2Ll3GBwbJteA16ZIfneAmMvdtrIfBmpaTh00o
HQ+zManqfFRbUxA7Nl5xewslBk0sbIDQnoSgsjCKSpfpbxE2fZTz8iWiEmwSw1oY
fuZ2XS3R2hZpLcRs412OOAkLF4VPw1Qdm/wSoqIYWghG10VZ0NjP001DL7lO6u4O
vN+Us6ZJthHpypOd26B3ygM5DEtYaJEiuRNfAPhVFgedyonCfjbttebkncWYSTBU
R63ZG7xeDDOfchQzsg7ExSeYbuYzvLy16bPlJPRoKktxA3U9D/Gf1x1EliuCULO4
AEJhr3KqOHc2mXjSLbzBA0VeugvC0LVvXdSqTvZIQiV+gmnpoXTOzYhMpMoOUgNA
pcsLRVwHyIJGWNPGBa0iEEtNXcB66NI5a7LXEcVObnKE5uVHAI+OScdPyv2Jj+vH
1pd/V0/aNBHnDRJIvT3rnlmCOpT0dUXcZdW/R9gl+TPmVCf9CCRgrVVy4QVLBbJe
ftQrThvIXCpyWQONt9f71pvzN8Gfb9x4GGNkOhCjWoq4OPQ3B/pnzfkskdL7hlOv
w8t2QvW1NnDg9uR1EPAENkGLGNxBrlssidto+qxYbbvKXJ6V8iwue1mziVpvghZd
05JWx1vwCVcWMDrYQgeqLtK7ZiYm/BjKs0lAaJLVYoCcdJKPc6pEOKcI82SjGUjs
zc0dMLZstSV0njqs/YqcWo0QJSiOC9vip4lIWHeqet0oignbfzOj0s1EArdh+lx4
az+lFkCwORjsegezYb90kJjBkNiC39K3Y062WXH0AGMtb9HONcH1d2ckxp96iVwL
+XId6eZF/FJDrNvjIHaNpHnmaEF6rBG0zKTa2XpPXM98+7NCkJlxDX9MqpMMcG+e
k1sm6Wa2wdqy560S/c4SMdRGGWIpr9virw02Y15YbPWkirUj/1tRiOFmpgmsiFZI
UQjaYpNIBzJuN3mlKLDWDTHC8hZbqpg6HoEpZBrYqJ0PwFoTxqbRHWrebROJeLuy
mfpci2lxcpbWWGEY77dngGbZ1i5IRBIKvgSK/9wGbf7NIvoYTkmEan9Fmom4JnP1
DbNVQMBwVXQuWgeENVrrojvp+lAlmMH5REX8zonBy88y8jzeMKcCsmRCa3jwqHF3
UQrFwg9dokYEgj57OEzYD9OQOiH8VQTkht4jBsFrp9t2+KDMkbdRML4/lXm2vhg1
yC/gTqz26v82UWlK9bFk7rfzfGdT8gugyE4AVJCqRtvhw97lneB/pnUGHD/8J7HM
vYXldRVRXZsKSUCbOxMA7F5rDL857p4tMshDSoJfsFLUZp+UCTesnIyCBwvyaeY4
0Du3cuGPnml81vyDJgmQDtE+Re73Zt11m0WA/8R2KmjfdCGqISR/a5dGW0F7O09p
Z3ZZTRfjDeoGFfQ1IhD1TFWn24uzKwEDG/eaSI7BVXnYPLX6jmHF/R3JnJ/4t6n3
YU0+EML0RBgwJwbg8oarrKWbgBl5+8GzylJsbLLHVvRKnY/P0XSwJ3p7ujtX5JTs
CnkbGwX4StjQatqg2ZpT96th99MvqxSHmhPMFXHfBD8QXnNkhf5nBBG8pOR+eWEq
OfFXxjErF1Vj2Ruam+Brfkn+rbKqmN556qBeCN6NfUx5aLhUc/pNPjxQWxnd+zDe
q92ljnJOSe3r9Gs4VIZaO58hj6HqntJjNfxVxdh6E+yYgRWB6qNW4MQ6xu8XjNBL
k7kNqP8NHGsHyVbmHmRiWb6YdKKDCBaStyboIdoCfCUwGpkDYdOhkOU4TfwBkyl/
zBykNVsjlJ754KgT7OIJQiLsxdbz9KbkidM+KwibZmbdxBDOO47NvJg9aZA1yJlM
294ITqA6VldkflYUq2FXcFQoK+nEzf+Dj0M2anlXLYxweEvf+GwxaojLke7DP2BI
RczhiGAPC9acyJRh3Hpj+0Q8Ma+9eXBL1U7sw5U9O4GuX59HQCmVbJIxHc6VSXOt
DC1sKT13Ab9AVLT6oRpIq7zMzBqUFRKGtn8Y2fy8NN0Zh6FUoJ5rtWbh2bZhNEaa
2yCADraTH5TaM1TVahEXzF05EB7Gz5ruta+JTEbP2d6r5Wt7JJ35M3rfath9wd0U
skaNPFKsZgiMQ6r5xfKXimzudiRlcxbok47JdJflbULK4izSUtjb4kWdhyPVceSf
mmZGOAq8tVt0Jl4uYiYs6jx4Br1VmVA+8ordGxUcDro6vO2VggIiai6ZG3oHdkE7
aFO4ghcnflXlHH5YaBRh4EP6HqFD+BA8MRq/BDD+LeE2I/2L0lEnC8E1/tVF8fJT
p5e8GPWap1cFLATC+ZZN+g4qhppn5IEDeiBC8aXku8uphr3MIYPhZmKUyDeqBX05
8w60ckXrb6Nl0sSA6GcPSkXsS7y2EJi2vmrbX7LCTnFsLnUdziJRkCIerHF4wmKP
mbUHXz91e3I1bhs5Iva61QUMmYW+fFNCfZsojaD4Mv8jDuwkFNY+GW0hwZPybns5
MxYpXKOBIXkKTfhGGLXLEImhhLL3KtYYCTdfPS/jfnjggQcMLh0NHYvNXJ+iXiJt
62tobt3t13VE2U5p3SB1Qvxt+ffD1hUU4f+o3PcR25ZiSwDWTA9y5Toj1UrDimZG
Sz7WlDqoUfpn26UK7C10xyU4QHZODeg8QQ7ZB8jy+ujBtnBCPA96BkFe2PjQyQE0
5Bl9kKRWXLFLnisBEavmk4Vwo1RUyOInnvTl0nazwBMucuQMKRBW6rnFNWqYNS9w
SJ+51Dybd4tNt/0GBcK5RGj/0JKB4ia8OgF0284GHAYPc1KHGMtHHXW/Boq/AIz+
v3bVAmA+vu6bXclC9nKP7X5tq442FCU0JIsDF912GAaWRLojWXkY9mOjSX8KrWgy
dYmA6n/VjICE5FIlCe0xpKziArVVFaw4lEtzzYepy+LGLKUtFr1BKsS2gRQWl6cL
bpB28/OjtSuAhwdUeZcvQ2B7hGmCRFFK5tRkoRkYNXG2tgf2Sn76KPfzLqXZ4Rw9
o4yt84mTKq0rJ0RFxNEBKMf6cQo6uhE+JAxWZEwqV3u8QuvpYhAOqetVZnpT0u0J
RK3NeTMGKRL7Z9OG3lWSIpRNK5PVob3NTWqFAPNw/DfDvdU28ZOYv1/Z7lNrwRgF
56S9y6yiM0EbIrgoFL0fIOC62g4DWkX6uamOTd1Z/pMSLEVB7PYKLgcOI3D1RDvC
csBQc4P4e3QOQQxyWRra4Dk84Y1r91p4tWZvcufmF5wa2brIonJVSWD9faxNRC/U
U4gTiaQX0pxF+lrUSweQyd4RefiWPC4BGZFKRCu12mYhXQP1yyzM8pnLi25Fyhu6
6u6CmpKwXGuyY3Oo1ulxS69/uwHjGop77kd2zTqg/cezUA1L79nX5zKPKZBd7RPK
0ieOO3h/QYzqCAQm6vya9VbkeoPArQ6QWQt4hj2RuLXyzssjGJFw3UX0SSuXw+Ae
bHpN2ubTWFU+bPPlO0+3aA7qgM2Qr9ATCmDNZgNXuaTxhmBc/9sBwXu8AaUlpBa7
EWfPQBm71McnF5FWmgo6K4GPOwmzvxq+ZqHUe527XRXcw3AquJF6Xrrejima2NYS
ubt2ZYXVvlLNyVfxprAfo3U7UkU/+TOqmaY481o+DH6k4USlmr+GT/h0BQwnGmMb
kANkhqHfss6MvPKqqnOmj3UAT1GbSGbAoAlkxt0ix1VMIU+PzPhI0TmH/3yI4zkP
7xwu1wDKUQIT2CILWwqmoXXDZWkHkvc2ZfXxLvBiHqdp5jkIQeLv7BZgu1KDLm3z
R6uzPyTGlRN6uPrZ7vwgCI0o5PYkSE/MZIENuuY2a3oezSog0ce6K6F+QhegIX3W
I234OXP008IfqqFOreB3bFtDl9ocCm3qrV7QBfmYWOv9+jP6bL3tMkZ0uVadTVhC
ttdmGHDt8PfMgvmS3IRqnLwogS7EfhRhd3Do2akCICYU3xOt1vJ0h8Rq8pYxOVHs
5zEuWJ1reaAYvvCrh5mBFYk/zhu6VYqNHRLM3i8qeV2TN79k52TnTcsTQeltF6ez
hBHOM6N4iutLHg2bbeTJKLREMcuqiT6BRFINhfbSVaB76a6UdIL6CRZKuIcfPNsb
JnpnxGPSwTsFAkeTXBh0B68xumRk7dga9QEticqcIqxq7bUgsUCVaL/t3eUPKWaa
l/4IZ+xZku9K5xLxco1wkaeV+8/djT6S5RtqLNdd6qs4AHnRXMRxQot/NF+mx+AD
lTtaGMJMPWctWP4WnSvBIs4v7Qi1gJTrPaOG5qmRouB8hnqLg50XnNnDJ2jbPxCX
S3ETm1QKhZ0EnM0miCnSz+/cCviQC+FtEQWPNtw4YU13seyhyjScJ6xssX45E8Qf
abZsorGVv41ps2GDeP+iuDr8zRMfNLmeWixHn+auxtMjvnhXc1uMokj/06FbJFP2
Mr2x/ydfeLxs4iDKYYFOOkJrwAFxe/5o2fUP/NlHYJNbAVvCCJxtr+q55rdljFVX
89gWRuJ+guaddffOYYoSnEbHOtNbX5aTxoQQtX6R1B1G/w5tCAuHIuBKSkd9J2rn
cM8zOhzUzri/AJ6j83CQiHj4GqdmhBvrD4XA0FqV3fK/hhZWj/ZU/s5Zso3ihVsl
/IE4Jl7E9sv3PUmuLqoRFWsa5gn9FDQQTd0Cx8cOQtZ4IQiXiRKL3DjOk1n6FsSK
/z4qwNwW+lQctcXrih8lWi3cvqO41+GaRsOOTFSWVGiNZjeYlPkoHlBJ7thxKveb
B5mYAQEY4F//qI6vOVP9U6WVBvD+iyvbp/R7pgRP3s8d9I6SXBjWctdgHScLE6Wd
5yu6Hr97NxC6zq6SCL3tEyTPBnfCMydLByP2MJRP0TT4Qgeh6eyZiudwMdiAhRdw
vXxMjF4nvTF0BGfx7ByRd0gtyJPWSZac0Zp6t6w5QQvplzgxqEoJnPkEvV+6YN+D
t/3ayEsCW9CYtX4KL5SDs2ZrC6GohtjGVnc3RKJWwFIJtWZP5Gwjlbbtt2RqkHG4
jAYp5j6UjcRGzZ2RNIoCIsjlSnh3vP7TFcMKGAqSHjkrgU/CKChfrlEbtjH1AHbI
uX6bs5LdxikidbQ2o58+G+iinQHkfR3S6OLl8gxQzCyk+vnC7hr+APyn1dNMLTnm
aEkOBtgpT1sKMF27lPQOEDvIOrdDpKHP9ARApKvRmlombQ/4QgZ/OgCjpzK46tIJ
7uPx7buBWuhVymRkCg++rW4cLxdZunzT3vawkx6GKuYNh0laCDkKJKYAU7NTKrH4
RFpv6vWo/9flGmGhxER6dMeMDu2ybtXlMukzi7+B00xFGzKnjRCdRI4OG/u4P/tN
Phcm1Px2U4XJwoxWzzy+PIutgDrgGWcGVb0gQ0wsDDP7S7i09DzkL/vaBas9uhqM
KCdcNQIPvSBlyhbjkJGTCf9b6eXfECYjqfQvxOOHpdKq372DtyI7dZfBLx565WjM
VFmej1qgHy9f6kWJHM4CuyA2RxDjmKbZSkj4p+yqUTKR3dwtj1oGdsvPol66wKpD
Q4HGGLhg3xhDoUd40JegKZHE28M5DHZEustvk9b7649WNWQe6Yt14xvuVUmUNM/b
zWSdJgxfxIyrOkFdpvhjK4V7ZfENSpVMHleMR6yurPwVJxQ2jp+koSg5dWIXeJl5
o42K3zncucmwVpLT2w40qxGThsQr4FW8zDiDhPO0qfjFc4+QK+xTrwkEteNt0uX8
Vyq3nYIqWmoP5f18j+DuLKlooXQq2LT+P9lz1wYWECR6mcy8wfWYzBkdrKYkAMkq
wp5c0RZQN2PCujPilnyIpe7lzXGMLxoDub2fYZXD5NzU5zT18sUYN8T3+s7gABTK
WUYm/xRHER4o/z9oOZmf9Gyhqlr1O83Q5JKgk5uFQe4p3ZWpSoseMfuT5qSpBuUv
w9/W0xCZk8bX3vRa3W61Qos72kQxvlvKDlRaf13ynXHWXlSYpnuU9aHRigdtPRhF
ISm47OgD/rbIDxNiF31ttglxc5uwx9PMQVpcxa29M4AxAbvo///D8BXlE2k+SvCq
btZXTemN8MNuyZLDSpyRCH6Xf0uTiwgfwsnuv0WyREPBA7EDeOV3n6aOiDIr+33x
w3IvIQE4OgbuhUubdQjWf+q8N2q4HXjdVm5/F/wcrX4I/dqw+I4GmxsFrSyDl5qR
RIiv/O3wFR/7z/9mXa8uWBK6z+hcEnSv4HavIu2RcRmsb6umbIg/txQCkEBEooaj
Tuq+NP9WYlqQj56qf2WeRgLZTLj28twWKnrto8P7aYMFnAlHl3EUPLZ5CtaZ29+4
jviHIPBeq9gClOZJ02GeTA3w9NHTCTGVU9Vvw6FczH6/4/4fl65ORSTg/gL82fO3
alCKKkJrvjxjzbOHvWo3zuP4KCZXU6WPKocxnn/BW9M7gn9zh0XGxO7CRqHuyzTb
oiT5GhBOFyf+F4eR6CFSlmdl6Qi2BH+Ur6S0xyiCA/c2RGpzUpq9O9I/YBimkStc
I3wpqOXJnAiq2i5u7hBb/66lUmhpAh1jmnzj6T8+bxrmm7jAp65vTO8ByH2mCZtN
aoiCdtVGq++nnB+51XTYlr95TDiokH5VaEiSXTwWvdOtzC0D+JnTB6eb3zuLUsCf
QWdPcWK9v33RFjyRlQ0SQKbYMDDGjIKVHr07aknokG2Tq15E8O4/XSr9U3CIMDOI
aRT7E7nXxjUcukRwIpWbQ8O6DDW8XZWI25bokA1uN5eWSjm+KvM/pJdAjK9GZuxE
m0jqKm1wfTlLrPFOAXAeTkwKHKTHwMbDvHhsPsifCG8PDc/WaCX9BuBl13D5dmi4
RULPd0z/jW+EgtYwMNtyY13Uj8niyyvBv0SsBB8bu/YdZCoAytEywKyw6Kh/pCD+
jH7l3uufP0nxMlzsmzk3VCSdLhmBK6HnMg+unYmFSy1MQNjJESdCWou9qK2Znaox
1JaqsrORpCR+7h+3gAdSHiXNXEC7iZP+jlbo5V+Oiod6GhOFKFD1u1LKoC8tut3n
GZRVKMzPfZSrcMEJ8ejciTmD2Vx+1tjuKhf/KHWPb25iqJFimlz7GEzu/GvBSH/n
J02DwqZLsdK/FBP+BJPfUO1gPd3JPcaaGJeUBu4ysYyRx369DNGB61Zaas5monya
6HgqKJMQ4WroP4VvThyzL8+GW4gHneaTZBQHYqbFnaonA5yP3P9VuQEPHaAwWKC5
xBOAINMx/B+UfVXXy8v1AphTVht+2BtW/xp2nxSMKTOwn209j9RTYDTnN2cKaMPe
5WUGKKBJhZq789HhsjezMp0ZYOun1Mvx/KuZedX0oAXzxUICF/1pDzpD7gWX3WNq
iCs66kwA2yRAPP2SO3BRFYPhNBmBCaHltBrhQDvPuSB8kH+BMqrVPTqsfmHwCZFQ
X8EkJIw1G2RyQmiQtRwhB/COpvqaS2CxLlJvMYjfleXrKnClenzn5QqFaW3JYFH0
p3Oy5Z8gFPd7YEJPGSZOllQfj3AGYP7lgjpF7LRvYgjP+49WTz5H+IiLUjyFdN2N
WOjTbWGVripcCCSMYMHkZMN+5ktez7R0dPeAkRZnwbR0DT6FacBKa0b4poiyIGPC
GU3Pplc270YeBN4V87vAf+wySnNIm3/ZfCOS4Vz7rMctJ//oGxB2cVyIFgH0fAMo
QXPeEls6c2qqA/zld8AipKge8mOOhaPT8W7bEBersyW9UPKKJqYIutydS2p9soGB
Kq3eepW63p1zClU+sVe3ol08cHsgUhE0X2UhxHcKBvekZuO+7TPWajg2QRKPIsMB
nQaXY0IcE6Z0Mt/r0mgiKDIgp3Y79KQ8XhreNKuAdl7Mx4tJ35wkB5aO73zJPmEm
HuLAH6Xlaz3mTlORlMncleKLbYBFeafb2NP3DoRgUi4vPhXYEqfqi5RXhTmIJXeR
8ZbcY51pbnidOrrAA5BeUJzHD8K3ELNxX8EFNdbo0ani19oMjooHJPaWmg3VaULs
o2Zsk/ElGBhlyqlymErkYyM1LbMaF5WkDv5ZQS9dddPGEgjWYQFj+XkaXwQCB3Cs
OPGSIdF42iRhls0a3WAvzRmtN7o4WIST47ZrpGSEjhARGay26X8fB1S6OYsauPu2
t/VAdlslKwyut/MEIYJTSs7b3QSER5YSc3sXju4GGUhi2rjRH4Eu+HPkSTMW5HUP
of8pwjUWj42Cep4MvuRIdwrly9SAEygAgB1xedypF4gul+6nkpPT1hQ+s4mP5rsh
lCctaPTKT4aAklMH4zY8z3s05fQyw4qlsm65omFT9u2C8i89O1ulBfgcK1WOkSzu
4M5HAuyfewyiyaga2uZSPuGN896eYWoOCwQ/49fV8pEKmV0XiHXq0K0WXgACO7O8
06pFi5+mMCZisZev4z4HMbDC52lGF7qkpLAvqSnPftXSgdXupio8sxalaxfOrE7P
ulZorGrya8vNNYqlpuaoBLwx/JEAEYb+sIr1ZL0cy/F5XO4OMpwnULZmQNvvYuUM
BekrxAahxgqRcZTJLXhQXTJHG2ekeGy5IEtKXLsT2FzLMl1KEY3sgAvUCfjDtKBe
9E3NdsoexBzDX8Yn3LexhLmXfaSS7cGUoNYFXRE9S9ILhXcKP0j6Np41G3TiFRab
zMk+lq3RElUjNLxquoRzU/3yj9GNlzIWVkCJB4j4SB0WAXFskmhkNDIYp4jihS3O
Dyo61BrIiKhKkf0b7tHIfkOpOOtBnN/A/EAIYZIeFIkKl44S6sfWKfx0VEWkKVEP
NPR7X1sH51thRqReqDxavCbsLxvaJwpta3TDOydWbUyOPsmxmtVm95TdvQOHFEbH
wKAuK5imNsdZNrOv0ZnLrgz1MkL0qVBrIzHUnctxIZagfLczryPVYeJahemuD4iW
AGquhS23cT9gO28/T8vCwWUBOorkcsQ+tGpSZSjkbqan29nSmUfAXbELFGhp18Jx
i5PYmGH8WpmYF0gJ9S2p0yO5wkG0jVbOfhU/40eBv9JLit8KOc0c47KQyeG7IoRx
Z47KGg2+jEgUTNkpJbFUjjpHgOn3kKdkaesxY6eug8makbhEd13TeUea+cCaXVB4
75mlLJc8aJTkAvtM6PGADD2AexEKhUd5i64jaxG+0/WTW0ZlRDqAAVTK+4ozYneC
37+0CkFDahPEx+ekEcsgzWVYJQZNsm0k/15HxDHsePVJrxoqck+UorUbTd4IdMsv
zPZebsjsuRirycDrm+HtMCzNqlTSrmMVu7U8SiUzSvEREnewSNqGP26G09k5oPG3
FX5FwCXJa2A9RAPps7RRcKRWUX+KUuDvDZQ+8qs3gUb00mT+fFXSemNd4swi4wwp
7i42TZOZ2rBrU+NZKsGvCncnjgHlW07GejpAgYwEO1sonY2/JlCm2Npo6LIqCRnX
Aa2V64diTHmw+16KnIPMTOkz/isQvcTzir792YhGRTSbdfNXCmcQOopKDs3XtRni
5/2dvc4zsfk2PfaPPTyFmZrY69FSOwE8dNvF6NSqG4yYz2kg0JrIEiDzl4WWiYev
RIWEd1z7QdoUiQXfQTfpz+lgXg9xhzfETJzAjf2Tq1GpqiOZRAHokEI4P6AFLddk
wWBilb9+PWttDCVKmqSsE2r6OuVsmaD0Ylo7U7A4GsYDuIm4Vi7GsJpW6y2HnjUG
GKemTIl9FR/cwpM1rRgeRBn+gtZeFfsdEX9/4S0+qKXHJ/3iOGcanOfKmS7skd3f
guolcXbQNftB2tZk/jja1k9UbAo6TxBfk9ine0AMzWRod4YLTc+KOicFJBRWldRU
fgFGcWVrY8bfa/BTCma2XH47yo4dsqKskIu9+4JAfg9ug47bmO891EnJiSIXxKgQ
pB/AE1SVWUDX/nIPoTBcy5pt2OlUw7pmBkdLKMZQYEkgUU6SkfYHfewDTW24q81v
OETccRBHH4vVVjpRSA8xUg+5Ghh5V7Dtzfur9aNSHA3U1fPeVmUtWjKw770ZpuEW
c8i2lx7K9qjNsAvNXg7mj1cIUMaZ0VYJKVQOtJ3Jce26ouZyXapS6vsdvhLmhpSU
QBBqIdplyO5Ft1AEQksUKdZb/xfbT3E8LbvXZgALx2PzonXkO2X0di2S+KJpx/5g
uMXU8ILLI006uxU6gIdE5nNjVj98tSS5fSzMRkr66JOlrf5ikYL5KOeNXmMu0+5u
U5X/utVfnuSYK9FyGxXWucWqcuB8AQ6dVE12PUyidy1FivoO/qeXOca1ZT298ixS
j/hNZTbmM3tlaxdo40EVe11MwLjdsuS+RCwzCrVCsTQ5KSnoe4f5jg/TJR/OHFD8
YxJYBwj1gdBTqmw9mamd4lKY2+4Jo/y2fFKX/brMPeQjPU1Ur1Vam2LZWu/o1nlo
SNDnTlKKvEjnpJL9bnnR+rp5ezVZGtiNJD/YTBbBtYdugm78FvjryiFM27KNUj0W
58ilbwIlWCGWWdxxqM+2QswmEV3WhZ+/rjQBBbwVbnHfQV/JyNKkc/NWgCtPJDxc
A88VQac1xB1S5ToCcZWd7R1fEvlbTwbogmUDeX7i7TzBURFrUbOEB5QyGW/QpNXz
cWfZRTByVpUfZCuZ4XsOkVge5hHxm8JvjHAYuC/iaAiFIlEJEVKu+3JsK+bNg+dM
lvT0N76pUSio9LzQEcK4enR9ZcKvR5bsWzTR3sBjM++4tGuFRsURGdL2grgvElSn
YAbgxVfkFN4Eqf1n+hiLpRgq62DX0mVLV3Z139MzevFf/jbT2O3hF8a+zGR+gz3q
RN9zXlrfh8Cmc+FNE2jSRgD/zb7OghU57C8SKY84boWkkNVmcgTvWo6lsKPwwKWo
mxSNRdBwPP+9A1XFPCdsiO/UieBcfZTWmFsO55LOE+b1I24WiDUNFJRklXE6/NH5
NEMuHCo0ndfjxySUe5P6itzl+cAFG71cWUdsgnpEPMUtpp0w2bUDyMUHzKPJQfEe
OkoF6FpRzxqBOH9occpr94azGy97eN4mVXTprAdhXjHR1DUy7Ku7Pbd9n8XP7m1m
heSCbrNYCHfCeVfVco+v82wdI2Ej3tZ1FPXUuBtNu24wad+sxW5Jhyo9OHUuiMJ+
n+GEXK5MdBRVbU22iz7DYbfgL+D0xcGUbmhoRnwm7AS53ut9hkiIAZxVrWaD0NMW
BqEAgX2NxxZ9SSXzNJ15i5jzckS8wNF7qVyMLwaUOIsXcAweAogbnZkDi4t4Vkb7
ujzgcMd2knSyKGjuYnND1wVaC/X7oIhGT4x5GFHHOlBzAbiAZY197oqA/mgbfGyb
lkNOVQRvexoYZQWjdTEe2T2BWNuPD/o8YV2XCgeYWgViFelxYxAS05wCE5P4h7hi
O6oYI1bVpWKLRVk+f5arBi3OH26KAC6AhWXIKkrkq7ZuwZ2aPfkDqYLJFT0f1v4c
A85F4vitoooo1CCvHhFyguym6ylGuR7uHtlXB5B5IXMoX1F3kFTrNTgKaG370Tcz
sbpSdf1vPh+NiVWyUeBKHX8yTVrO/IYvmQjL0Yvbzlo4H9/8Jusep9sadYF5LPpT
0t0sZb/fcWgptxlIgK1jnBpbxsC3dLiRIc/c0IdKS1ipGQYyb4MgMGrunIucKfzx
Ggg0rvn4eST8wUYzG7d6k+edIQTgyWLFIVBnE/ZKPNL0MTAOmxeEH4oELyrt5zH1
5VAt28Y2I2P/T1rsjmY5bFYfOiKct0LCtEpduM1tSC73LxaNPoV+YYjdGCU0FHqo
Ow6+CLyzHAW9uf76GUyeb98kdGaL4ps09tEWswfitdKAaYmeruMSak2bvwqQ14Eu
RBJ5Ya//3h12yUtHlTRVKfqowbWrhsCi05I4VDKv/ItAGRtNtLRVshiWeyuDStAg
GjMYoA/nMMM7vfqPiqlvgDZZyOAehHC5Jz8qIWMRUtFE/INNKUK2tFsuJuXj59uo
iFYzueGIssI/Kn0hbO3rV+v7QWTE5UfVv4APZkp7AKNPy0PsI6eRgWXCYLvXapfB
Ce1kfzfiduS/uqluqVCTJ21DvUojp3Qv/yO4X8jbjhMUQKFkZ+oIpbD12ggXAajO
O7fOlLGQATiHwoW/e2kb9YtrCuG2hvcNFec5ehv9kKgYIe1OyD+igu1GNxQ0A5z9
Ng5QqEiTPkuttdJG2lO/sZT5w19Vux7xCJgKFhgFjS9r0gdBfcBsBhRfiXgzj0/0
cZpZuTNnALvfUX0SHGGmfcq9fDnnF+9SSvP4MJKCdLEf1fXM5M2vvg8Ju7eLLjy+
dTTvyTqu5P9D/0Ttwgm60c5QfORMQbnwtofDkB59I40/g83HDDy/TMe1q9yrHzuQ
EOuGZFrbkkDXmoY2H2w0I+O/a8a/CZQF3Q0kT869LIXKZLIcrVD5THIwOFi+p+IZ
Snt6cXhlLt8gGBY+Y9TarYDisSRkzgbL8Oabb2loCepA6Cuyhg0IT2nwXuVm+KzX
pjvrtdJHP8R5a4v6ZPUcMDDZD0zw0N3OADgw8eJ6yvqrXS65QmqEv5iv78Pr0ynf
8PYsNT1x2vvvxVlKphVSVBHBNdOaviBXi2PMQj56A/FPca1MVi3Ju2ttKU8x1puM
hNnRO1DfD4+4LuQCAg3uBvNcq83o4ZAmaNHxwgOWeWP70a/82v3gtSGZ/BOY0CoU
bx/XAgpmnHQO8NhE922lrlX+tvpmTcCCRBdacOBzb7TTMBUKB6V1gR/lUzJODC/s
e/o3S/GQzV4Kmrls8iYIEUyrZdq8Jvq3FkU+BGIYS49d5SPTZSVf5fzJbJzccF/a
0Fryp17qQP+Njd50ot5qFInwnHO2n61ZT27UiIGgHob2l0Bu5ZbBUNZ+lSSiUdeJ
9tNj1m9W49QfJROSvl+jaQVbOY6M45IPryucc6zIvqzHSLWJwh5GRlUojaP79fSE
lFc4g9tNlbEH5/qZT5trn0iRR2FW59lZsNugFcO1VoLLRNHuQKIPqqP4vyf0Ha5w
xwvJOYWd1rSLe+3+3+laUy5lZ0N2oB9aFoBDeuXU6QUEbQYafiGUQjU+SoFZYJdL
lq84kwZjL3QS5ApWkXXoTtemIAvKtNJwhzpOKeFa03XqiCQJml4u6RuoGhEwdw+O
2N3l7CeVX9dZWW+oqRGVQ57faoexAb45NJ34Wv/1l0UdfMH09Znh6T+WZsSgOAHo
iU3kjAjKz6oBZjR48g0SMkP9EfpuvoEPTJ82YAzs4mzeVZUG5Uw6E0S8giKaFsd4
EBVSlzcAHgWyzmlaWPYNThd3fG3gU26gVczN0nsiplg80uGu8Q9kiaKnfgUn+fzV
8Qdx5igWugymgschi3ehW5c/a8DWimEWN6xpPgYbZyEgOZ8m/a6lKmTl+3BW75Te
UF8bWKwfk7+WJ4JrBa0Y1/Mkthitot1Rb+dqiyOwwxyUsmH/NfUKzoJ8mzB2bIBm
Fx8vjLplUJ4HJ3QD69EGylxa3ihfLPWK/Rw7XvoBuQRYZvDurQVvWSEqZZo8TgV3
4az804XJmcHiR0WC+TVEgWKa39KYeXLFuG30lc0me7fkM5t0KF6IosofoT8qweAT
J7Iu0w/qrvOAMs1fC4yn3hBsRde4EeTSdKMTdDHW8v0t0vNVFkWtlbSEanz03HOc
5oUr+UuOB+YFH+ZdzkYDlirECQ5F97I+rG2viTJkaQ28qltnvLnXiIJk2NWZ2cVY
zKkaX2CZcisM/KFelIzmTAeN2YeEj3qZqGnE0PFqOfUYMvG2OJuXqgdUWiyyxQnh
HdWF2y8fC9wRnM3fHmRknZSWRlsjyUHgnLr3MhTUA65uRK647gZQpyEVL2rEDmmQ
Vx7+v6bBSY4+zIjZ6SUjAD1NStfH9v8/fW8KsUqdmBTPnOAcHG+c2JUVr5OFl9fl
mL5h1WRV2nsrRI/9jhewmMvn4lCCvIuRpucgn+Pc7Mq7U+2J5n1CAvB44YdS9wvJ
mLnpQGOsdLVnaBLMUOMg6edm1Z7cx4pxUnsqn5+VxlXKOkae5IizK0TSkaJD4icF
1gH8cFz0KKpE3/wRdXWJ9fYxFm5feRij4qTmm2uzXkV3lsYBiHMhxqverWDZL329
2k3J0ObLPavfUVUL/+aXLmC/4z0jBMbSTgoxRidFusBTxYiNn12LfdR/99WG6VG0
TKVM7uNQd3M6rrgDLe+JFlaQyICHW3HHuYL4XSvupP31TARjjy9vuf+dL3fKaKG9
cU5SaAzfg6NATt/T77Yo1+gaGR3vxwBsAALQFfRxE7O9a+Fj49S6lOUA21NjRyv5
mBnWwGYyWgiu5ZHfxGKJHTdp4ydTg07TO3eGNL6G7TRA848kLY15tpNcPLbYLkF6
m434Ty9EhQgHIJVGCGvCdQ2O/XWY6T7NcHHXBhG9AwFHU3YtAmjeR4WXIl/0DzaF
unkHoJgrPrg3Qcu7UcDRF6SE45MaJwIr1uEPWv2kNEmG4zK4UZ3qHynt8XqYZAmV
NAe/woMaqz+I1jIgXiirLquktqPVw0IillhrkUgdX4ZLH+rz37KwAsyootxBIfb0
jjSsVZDQ9lXtwSLurxjBtzqk0P2maP6ysIhkQQoWWVhhrO0f/jFHvHQ1K9zLW4rP
qPXyz/NQLFhSoQ8dEMdlDmo/Bg7Q/3xysiw3mRk5ijL1KMIPf5wfDYhPjbzX31p1
lHIYmlnpjT2oOUIsfbZ1SGWa8hG+0oTHUkhvlBF2cNAiSpW6ELhV9DwCuZe/4ckF
aRenBPQdOSEP1hz2+xRM1QV/398t4l+3NHQgI+l4C5yKa2CMKCzFPHungyMt70Y0
KgMUswRT8PWKSxfQxhc08oDbas9Y7EC3QEz1ARhD3NZncBgnjQmqQQFdSiBi/J9D
XUPuecfclrKgln4f858UD+j2r+N+r/knPb1S63rF6/2dtRvIqMIcwEUsBepBfaAv
3uJCCREymgtsHRvFVryzUnhwhok1+aWBy/6oW4OlrERq/yGQkhz3mHW969fDHXd0
bzoiJ76sC3STbVXHm3ipfBJus2J0idoT0DZxtL2NqNBecP2FWXeviAmaQHiQ8iRQ
rS6GONFf7OU9rwNpXXcdkM/DEJOr8199s8wvTqNTQIx3TAoHLL8b8u51S6hCXm/X
uqlkSkLehkK33k4MgcOW4ejIXmKuleYkanlFne5tvF9GLp8h68O8cS35fYxi/xa1
MheLXU5nGkb3UZ4XKF3XnoFSiMIPfdxX06SxgtZXGr7XgaX7kQBgT7xdZYRXCj2X
2JtBbbcOc0lEpG7d/q9nlzSVU8z1O2oUNHHu7UEwAgfR44vFUNZ6OBDT9D6fav/o
yjX8EDechruldng7zd+luJb2Z6qa/mHCgwn8AafrKNi+1Chw6DaIQJ41Q8cScJcN
iDq/Xywlxm/bjO8KtaZ8L8s81/PDAx9GUS78u/o5X95Y66i9srzVQFmCwfPOZeSH
ttnuokxbynB8ipe5j4nbuV4Og73jfBBfvLtvyfb/W6UTSDL4lZmy2jRuNIl8L1mA
Kof2MSEEv4fSO/6BrB59ZUXbeQy7C/KVRxtP4hyCo7mJprf6DCBYGBi+VefFoML2
iK8kjeFey9GEBRPmdp1NMxcyKjljmEHdKiSYTMAQBuTRO7EeLP6UTvaoLehUHJ5S
bXCAYpkrhnGtoQR8MIwzKTGPp0Xkn27/hR+RekDZvai460u66tMowx08jURwTlLC
Zj10jdKVXUXwWBT3S5HOcYogt5/pwBJb/DO6Lw3tZNBFXpA7V8HF71BaWPVgcboc
1KWz54/Ft33tBPZpdScXManixVVWy4B496ZvGBUlmqunmXVKLSRh8qQQ7ftX8AiJ
/0DwxYQHhzb96aF2EtS9Cy409htooYfWr84W361bcwSz5W7d/IDVPdVsp8S4lAkH
/Sb4vCvy+5NxyrtQWaHAGim4wK66UyA+oNf5P0tDWPWIOjoeBwOYGPkRDrNawd95
F8P9yAmRZQNmJIXXT3PFl/RRu8W517jn6PsUzKUXFHomqts9Edb7Ad+L8iWkplRV
y1Ne83Hg8/jDMCn1zTb3q8saOq7kujrcBvM6xK8DWx8hAVsmelunvZw1LQwvOINi
EogdP3rxpsFl6Zybnububm5Tz79D5nAg3w97FAPRAFhb/FiivIF/skVXY/TuXzJi
iqY5aAgj6Xnc0DOoxmtXvk5aV1un4D4lO16DUAOTQ7ek6wnlyiiI5EIw6mQsmBs+
A9oUz2+AluN2kDsnPrBJO7fVfg+Y3W/pmlwwqlUHmkE3AB5RAzrwgbJj3aNeRgSo
X8fJENn0ZGq5+Br7URo7vtQBuHqGvwLo7iBdPwS7GXMgEY+9zOn8k0D0imRRUz7B
prOlZafvAA6n6ufmKKv0PxTRIvRjxeH29gTcu52EhYgqv4BJtI0Zu5t1VmZ+1OTh
OoWTIzMg9hauETCxy1rbYuOf01MgMH42RqnROiG5WThpBDRUU7wVHS1fdiGiHEQ2
JgVacqypUt3+ekyzIdmJdus7DjTu09do7TOP2C1H4BG8DxCfjgdIA1U+cN7iVtk/
fKX9kxfu54g+4M7gkLSscnz85zwi2ut+xDcKGk4SoVunD15THvNugc6nCoqnoaZK
vwV9VZ7yjyNPCEB2bmSKOEzFiuhlKUm+nLk/wuOLf8Y6wQazilq6zrpJv/yetW01
L/pcsKLd+Kr01lx7M414D5GJi0s/MmeK0lAgkKx/DjqzVhQ4qrAsGzbfccDa+B8y
LiCll3ARdf+uqCbxD3xPMv+DXdROpmu30k5UdpetAxAXg/X/F5klgw+Sf/s+MRd3
IaV7NXZ9d/l+S50P2rGzZVcA5sYtp0Qtp68PW//SU7XTt6hAZDqofbHNuMB5KcZU
0R1xFN1hHa/gzzg6NRiaqjee5STrl/1V95EcsBpGWnwts5nZmemWqsDqQ2RSc0MO
+i+ybEFWDR8XV5GMZL6ox/2MbZxweCTPXO3XqDy1pBR9aU9EMOVcdzZrwhUzb6yN
r5qC5kv17G5CHdXJc9IIqCR47CUd15g9Fg53/GS/k5dW2HtDRs7HVOCqswXKwwlS
JpwZ0zFZEvdH5j+H2PuWqTGFI1pQfSbXU/lZ8ADuB3n6Kua66OkFdVFeJ0NDmQva
b09+j1eaCudQOVUINXhN+JPyB9LqPXKteg453qeraojxMGbAWCMjpfV2rZk/ckNH
bvIKBsCQRPg2gRJeAedbYkNyXvgKZlgqYnfqftzLH4+SlXxTLc0QrDE2f9f8j/VX
fTVcdCZ9dCGt2ysWvy1OUSxIggBmefKwoMsCiB+o0jgrSAJ1JMCz8kC5c1lpppNT
Mw2A2crt5H/jTnFdm1Cq3C09MV5AWYxGwK+HdMHHxq+TtfYlelISHc2I5ELegcWi
/qzznaKeSJOCQQgI+ldI7NqFOBrUW3z+F4eI+sBTvHnu7AJYDaVGa/EELCt/bG+t
LOVyNFOYZSgMFPM4xyF5wsjJdjDVEgSw1dHmjCXzB4qMSm5/aMCdKQeh5/D7LCRd
WeZsnTHFJYJwhTQKj1GVivPr3fm9PIJoQbB9ep48ZUTLxkqzxAhjBCH+6sIPFsIw
rRssZV7KRY54sHwGcyZrrNOBUqj0FB+gB//GrLxU3ePU6X1M9WBws3p2Ytl4ZJwE
AkrYVpOuxs1vUGSLH8aD0+t168ceBXrcdUqcHUDWxIt5vRIoCBLxejcpRikJDtK4
Py87+IuOlqWD2mnmh956yRPGApclGo5a0l3cKE/Vuixs5x0yQGjUv80jQpib5Xjc
PcfXIY4yt220ahb/qlDzLPcuBf0WXE2XfCQhp4n0hnX0jJm+fL0tou+6zAs7mGFs
TaLAJN3ucYN/Uii+Jc7FD9bbncZfxxlkZjAvp5xk5C9LzDmEe2U9ZIh0G8Bp+F4/
QXHEekxsOVGInuYaElbZlkmV10eJMQjZx+DQz9VSyCylXgvEQyTYBqzypIdrSZUJ
SHWkEr59Ull30jQ1teFOYUP/vCD4DyFnjhbJIEojM5o0zU9/uFpFhCuF8m1FSqzA
rDUjffK5SULeS5KQx3mLhBXhJQXVLGai5pzdRAc3k7QXA9uIaV/MSdGPyeAWPOlH
3EG1ehX36Z18vVyAOeLW2+m2t8c9x+RF16YB2eF9Tj6LX9ebYHY6FABN1eArNA76
BKlS78ImgohxskO9mT6/9suHyCLR/FyDiwJG7vbAQWB3rBrSu1gJgimBgg9sN+V6
+ieCJP04pPSxN3ACX+1ZAhArzzfocai2QPmexlZ3l5D7BnCHRadE8wpgjWyn/bL4
oVv/Qu6mweDfto5iRF578yY60WA0i82Kt+LnOA3NL+V/z4DSlFXDwQGpPfQ87EqB
AjGhY/64aAZJRK8mfag/oPnW9Q431lnP9zeKz7LVXkRgnfmZzkOiYjZLbHknnMvD
XCJzFIU1ieV4UfFZcKU4OTKbvHjCAQiGlJNK7uM1rntMuCbsVpuowTrx3nWEE2YE
FF+K7Z9h761KQnBN4P4BLpkvEDt5jHHVc/xAXfwAsp6uUZpkiAD6JpN0Y1/o8L0/
cVI5aMGOpphHrzPQcvizm7S21eT54rw1b6fs0Rnl/rUl45Ra+IP/hE9GE1HqqXtT
xHi0vIzDzuFlBFvuppE4nRRLPYlrAcKlY4+aO0jvgCTMcmbf5LgeGDE4D1VdyCPr
jNQZWgREXT2YNXvQ7iD2HcaLT0CiUrPdjqQhtD9sM49+j+pGS0gjxudq8yB7DLFb
pUZ2xDfN8u1bS2YlyrbbxFKAM6k2Yw+pbyUK9n7C19qGR9bRA/C2A6TSDFJFO5Zk
Mzup/C6H0BSkogl1rI2pRdkeDj7DQsfby2opSzDdaKJbovOIbhVEndSQHD5MBFAm
ED9bXAle/DeZzEVY/KdXG40DZyrbEBKV9rp8ytxgHnN+yuMU16Jy7ZGAAUFTbxMt
9pfyvOiAwoV04l3dmyTSklEZojPnZBN7541i5pmOFPmc11QN4feZ60AIDAGNMjF4
IaYhZFUD1HjG5z0qISFnwKd347bXMtJ967RyqLMb7cc7hkNrLxuyChB1mg9BLgBC
4iOM2McTTlCFdTPvmdaGh10FHDtru6BkvrFWltnYjN4vfa8Nq/XFp9pCVUzWtnXc
VoQIeLXycBBnFRzklnOqRO9kozzHGUZksZmqLn6SRyYEAU9KtsZ3gRwrdeqeWbL3
ZIRx3CoRWm8lQsVKRQxBPgUecFHO/H+aTprKkjy0m3+UTqlEdF7oEKy7JhloEjUg
EnAJe9LUgrfJ3x2pBP0b6kCO8F2c26Afc0B4hubuCf/eze4SsiyTnOavqHIoTb1E
hp7YC/j0mPVqw5SjBwAShno43LGHYWtl3QS2dJnH0wY/caRwLHCRx1MkiMYmeA18
M8MNPHRoJCjgWSBWMHdWCh2EHECJYn+Svzwrlvm6qXpa0Kl3dUa7wvPg94Wiz407
Q16pugtjr/bqI6blLoaHF4LCzfJffoS4u2bAzf99F7BOCX6GPpO4havwN/81qSNj
MVY9P7wK9nYV8En7CeKR/GSOeyV9AVf7USpHCl3IHKxginx7MRV0JRyWLNRJcymR
t1ln7JbZq5Nm2awkv/+O0nh+6a7O+69m22iWK15RSQGnkUH65ZkK0L1/qgdPcmPz
Ne2EK3WAFb2+lEmz01q6ISzbs3VXUwccF4xh1lKUesfHPQ5cjqh0Tj4fQiI8J4FR
kErc7kJJAfSHcdJBRcvfn/p+HHzQnR1M7RTLTv9dmNB90o0VFTOv7WmCM0qiAIql
Og05LMKm2we/N+0eKlweMua6rMIWHkBwazBA49ClADISgXaJXYmW+cl52NkoE28r
/fCBgH2q0obLfU5GcKEFnj47/viYGyzdt/Yzg84kL/4V9u1aND/ZyBRIH2I/ikZ7
+BNyx6k+L5eteeo0yjUhvpbEnuB/xufzerx6g9OjSiwGYJu1t5c/+SQ3ILDG5m7W
+PyyDTkOW8VxQo3JNqPAAXwWMZ9HwjZZiU0TO5ltEabMBi3LE3NR/6GJFE1+Bb//
cxOIaNBjgOTmK40W+ZfszFXqoVZJTE27lVtHnJcIeIHgs46XkEid5yMPUXCnJX5y
VQO+H6+jKtWjtcFVZcxb85W7VRIGOeCL4IREcprqyJzveRI0SCwiQCqiKhYQNd3I
JylskWsaL1r7MO0d26uu/nPTesf3jeQ7tnd6qVSWsZr9D5h34cKg21HGMJZaTggm
I20lF2tskKlA9JqMkxgpuaxCtIur36palObyibdJFCRlfVddd4nXBsOJGmMb+9nI
lSnBs1XQgbZpnfwVeKovyhHMkwUdzsioT+S3T2qHD3SHRkRWmnjAikma1IW/GFSe
97aIsjpcgPTqL9TfSn4+y2x66qSiO1mSN7l1oJS9AiblmL6v7EHAsAm8SLQTSlQE
Io5dCWy5ugNFJvOE2MkV0UnsW6RrRakXddnfhFDFKYacUCmCwIxCRylcrV5ubnqG
p/nYXOyzI2/BJyj4WJKgLWeAWYJ4wnrv+Ri4eKWBa3IitJf3KBGRQrBcplPzGUkU
5dn6ThHlqXBvsLqZ1kPgyhFXCoGEjNw0/DIqGMiw8IuzELPp7+qtB9iZ2RGGGHiO
A0RJfq6IllLKV/XhcWjSbOqsSQRjLqeEyIiX2Rg/adx6jz+8fYhiD1VNFEHC4Ey7
lgU/JZAQo1umrfV2sZOxCAt8cCLDkpFQOKv9efIGo/Cu3oniJDagR9inUY/2LL6j
1Yl6Ox4AbqcELzwfZfI3mMa1+30qMIbcRKAlmRLiLGRAwvH/MH8A3k1LZkNYiwu2
qCmlDS65JPEvL9bX/5lkw8DCU9+bAd7hF5TxU7D11T4UpxAj4Rik9O9N9MgdhUPS
ldYh8MSCPzhcjsnxnYnvMdZHz9ERoqMPY3mG783XfD/kos6f1x/Xhfit9yCQKGnX
6cM6/dWqtG79dnZf1XDjidfb71FyqWSweyJ0fqUSRT5PPUGb47k0YsbaQJnHgLp2
sw04rXpp2dsHkXZ8OEe6Vaxomzrqi9+/HkCXO8WUQBmNO7i07HAJZWw72KCX4g7+
gvPF4pdhhyfpiFH6JRTUkrMWOkzuxJxcudcQaJ0HREevFsMIDOxuNS3c5t3og0jw
SXj65GCsUaSI8nBzsTXaBAYrHBe83DY+O/n0GfaJWRjgDC6EW7a/6eArIRIBTR2c
owBQx2/yty+wyevKdjKcQos9WBq6PdkiXuEaxPXQon3ZNHwjr6H8GsRipiteoV2a
98MplArzYFWTrpTxlu/Jgc4rAAYX3C0oDTZ5+xWnZ2NK0a+94b2dKKgA53MWvqp1
OVY3Q41qGdQwDZdVnErWscDbK5Dk0KAUIwlour36n1TyhbRcV2wCICSB83tia2cG
rZ7rlDnjjvv9oqCv+iCtPFaQS6H3aHT20BVRMAQxitqM7ryRrrXm6JqcrRkulPCX
lhAs2GTCuSKyW9EXmxpsVufQAkP5pysbdBfzbO4RVAm+p78U4WoImFHhdSLShgmW
giIX/qLGBCY5qMc46Locl93mIbgUisB7X0os0SND2GAcHzTkNcdk1k93adEi6yEc
Pxs+8TK7ohXbJ3ZPOB5GThyDCGv7XufVR104yaTALug7X48hgRXHNRXoMdtP6jLK
9xL2qw+lE4EJDHhyjotqZV0Kaug/oIcqcAdcIkXhq5utqmkQLIZFqEC/xsmvUKpd
kdK4TdiLu0angcGszIKQNh0a8dZt9p4ixmnRH6zNJJm0ZyiM05zw/EdKkpkHYW/T
2IAsZwOHLE9A0Sh+FkVZ2BBTVS1eN65wLF8iDfjR7c9x6vJBakgTvounMCNGOa+4
etFCwGSAv3JerubhcLOUbebnaR0k6BqxF07Xh4oM0kWZlb6Bv5kUjfJT9dNrYZX3
yeAoQbOzjHvfDYEZw61+6J3bP3A+cUynyxYY8ILYRVRWCMe+bk15TtXRzriQRlHe
8Q9Sfs3doMlViHCAZ7JCe2ibdRyrFJd1hpfXnGxm/7M4jOU1/fHAeC1adQljzUTy
Up9W/QNfttcJl4KDA+Jo4fxe+u3ShTon5wUbGpgi3++HNrrVmFYTS9uSKih2CgPq
7UrFQEHvhaoWw6uWBV2TenWssYnPxpFYQH5DZDCvMI3GsyIa6ESVj1jYClBhgtwu
ewZwmjhsSb83G6/TQTm2l7ea8Nnc9dODT8wORb0sVm1uknSKbnbnLiD6WFCH5pH6
Jg3L8ezgT+b2Na8kR2SckGeRREsTzMFTCN3i9XvST9p1mRQBodqZqZdhK5mauRzT
s7YP3011x57+UFETqNyomAi/41YcINTDBF2p55yMpPlGXFGADpTRz7eEgFxpJnL7
f/JwlxCzE3AUe0SswcocsKFtxPZlUgvM/YPhEPLDDqzPVG0ZKw/IVQ8DqXJFNlj+
Fbg45AkeUfxo2ay80lx2vL/zUg7J5r13ppcfjwPSXtucch9nj46xCVBo81TvitpE
HsquSpqraIg1GGhr6zAl7EL27eeIbSTEHneJlRH+FZyjx0gl75+8jiTe4mO6kBDj
RB4hvCxU1/8Cg6aSoWld/sRjZm5b3KUAW24gcAFBoCp49/QgVyKw4FmiWlyAiwpB
DL+enlWF1eRs/DAokVdwlGjAG/EictKkFROC7Hsg2mx9OW4j2ZydAKfXn2wucMM4
EiQJA2sSO4OLmY6tKtfvzNr/w35XKbmeSf4eQJXhbU84+tFWpTV1K2OJ21r2BGz1
KTb7qAQ9Kq70+azOFmnnlRwWjTYGHALwOPu0C8tSDK6tY8L9MZ7QRZCJNk7VHsKj
sjix2QTCz6pJ0Lvx1ZkiuigDz/sWjE0+K+TCqEVgF/Gbe/dkJMD22p9oL3BbD3b/
LwiiHdQvmExDf9V2oRIWq53MM79j9NSWgTuPP6O5d6Dn3higuwgjHpiLXbDALe0b
s79Rs1iIb5fGzPKyRg6qQFZl6tiw4oJVznc5NqnAsoWP4oCoGjivUxBDEuPUpdlT
3uBASkhXPXksvF/UfCScyVfgVkvHbgn9JP9KOLOhM31mT0b29y3XWHurfPO2AISf
2Dsf0pKhitPr8y/B8JZRA9wE5YTOPblSTn1JfldIxc0FPENc46Je+jGKHgcvLJCR
XrFu8++OyNRJ39kkfZQLRzk3pyb7qeGMwKijgNFROR/qYIyy6/FP6K447v8h+/bK
Xoxq3YoVnEKrx93QWKNS3UMCqmKUldWlJ551BC95g9FIuWVteaAcr8cPQkkzpeF+
Gtqhpx9IuenI9zgvXnFX6nNeayo7ToPodTUoLfIYjacR5WTFcEzZSRQr+d3ztBqF
bZg02Ax2h7SxYSGUUHy3FiZAw7/F/xAxROAcfokHJgUqlrL/hOmiRTMHiVVgO8O4
58gVCd/B28Uz/dzjos0X3uiyJAxxSdZUQeribp5watYvYFEC+gOC8DkbE6n5xpCg
gNgj5dxZy0oOEWBnJRoXlTg85LpxWBqmNGvCeJceyRLH1BaNx4t/QFj/7C1+q02s
qnfD9hF2dqKa7QSyGbA4J4uirludeceHfsaC5XNx9pqIYzURPMm/icQWfqL9cwuO
I6EspXJbbyuUw26uH9UpB8nBVVEfUU1n73BCRmmsir9gnxpxfCAGOu1ObR4zAXa2
8ooSh8OYDndCiQ/oGMCLbJmYim7t2rEEBn6/CIr9Mzk+tglQ06ViGbDaObMd3vI2
LRiKSghMydLyIumGRllvnKAMwissQZfezgMBpYen3mWfea2ExLBnB1O3yyPA8/az
q42SG8aw8cCmABCqBPxdi3/9FLvmX+DcAzKYkSkpBAbvr+J3FnexmkyS4uw7mzEI
1tXJ+yjkKtezlksxO5GvAKqzYglcp5nmmpG9TkwXS4paG0HdviXjGZd9X1PKFpwr
9JkfVjEjoU+IXe53OkaCLmXyUL4o1z65Qp4YfJgsgyGB7TjVbZ1Mo2hpFMCCc+vk
/KrnUfbFSgmI/8x3QBhCf4Gm+DaNnuIv33Ml/Ax+vNV1HyVla6unmV2lLtIO6LFP
9Fa20SZ0J1I1qulZKCMI+Qk8v21H042FPljP5so/P2ajCKZ6p9gmc3omp1IblXRU
wUfFPtq3lp1o2Kj6kTcfeuN+EeGLHjXZsk/GxK+2GBGor3T9OWWDUkmjGuP193EV
bG4YHipMqyF3FqcN4WHz8mVJ5D0z1pKAWU3gwM09RzE7it6fThQzPtQ4VoLDpos0
arZeZD7GNrz7N3UDjN2Kw+gnmPEkCfEbU5G3yK287q7NH8a4UnFrcSufEpIm6yTT
ahz2bLN1Fja1oZILF/M+dTw/4gZc/mwOxZKzFLJJgDbX8V8B2bOup9uoH1vp1IOH
YL4F4pdU6f4xwkBjMCzzNpqwXIEycQ38EUspKbLPQmm05Q+uCsmRlc3cvAj3wiL2
kQXmZ8ydYqczkdC5NIGec86y+hyWnKYKJ+ysa+y04fTnkby6EA3tapvOiPPMe1lZ
9zsV7zwoXImZlG9pVa18XF9MRE36BkREVX9UzJpr134EtjcvtbFBfvkS4nWv8m9I
8XeLDmygj+pfcJXE333mEpU3n9LemewF8GyF83RoFl3zoeHcFvumEIx1EQz+8w5h
XrfuUu2V2eteeZ4DGSk0MjUuikTs0jGj0eczz/Rw7csA0+JAV9hil2YtEyZnr3j3
AwfoJdaVpxmjecKrnjRgITT6LXzpL5aVY5A42NRsDt1AV0D98Ix/NSNnAFMSsSyB
Yjcuo3MPL3zorCAl7v9TiBc6OLm0BLRpnZuxFlZQGN6kLUvRq/AIs/2rZvF/fGkl
bpfCd/28KiQZ8yKOZmYoU5O6CE7hmGjnEGKOlWe3FIEvtWMJEETfzgw7bntZ788Y
zFbE60o3Z5Nqq+VaI8ZnggmZ5TXRm3ybEcUyf3RexV66uDR8cm5fJkQQ/s60mkO5
wwT5u18GiAoMuoCKckvbJ1N+j+W8K/urXPuhpxiAO84wCiBXeO0kbD3UiO5KZdFm
GsEWS+bpDN/Og9SBVzR+cUNz88WuUIE8XY0EscRYDiWLeFFir3zTuogI9T6pJB2u
rusB3rQPh1j5B3iQZZF6VtPj8mU4ICRKzzcVZpM3w3p/NEuH9PlPPQOokepXtLz5
tC+ryICf2xFpzolz/QisxUPZE38Xe0DDDVnnR+F03eGBgpoIL/dboOsp9VA0U5wR
lwB3kGgQ02SvolPAp+UEg5bZU//o6pHyWa3DwfzjKy+WgqqWUN6C6DsQ3NMW5XFM
Mgnwf3K8QnjoisBWbHFSYdDIQkcbxLZd13ZxIA0vJ7mY8eOlYUMBnMG5pnIWpOGY
ug/6X73WH7fIQTYSlp1eC+W40pNQnblLdAHtcpTtdn4CaEftHi22lVpBbV5DTFgy
X6NJ8CsSQDI3JXLJzo2S4N51G6MpQUZBNpNOCCl1eMsydZ/IulAJLm3eXRuxrFE8
HcJmuJO2jo51dLZwFSKwqoWspz60IUj+zMFJhY9xfN/UQXMxiRSx8ZvuwO+CwRp2
vJEOfWJDHIdPZ6K0mJouUmdnDVUmArVWRtGFW5MdCudEpA6TH/2Mj6S3vArFoH4G
NylvwNA1h9xFTTKSzp/aILrqy+qWXNEIuVcrRG2HOHWIXq+Eba+UkQaSYKvdzr+b
Yv7TcbIMZ52TuUKNIiHEtOU/kKeDVzDMJ7B66jZ8GRJ9nDxOxSTho26GmwTCgn3Z
2tvBcYPyUJmtbYxnOQmACWQ4bluqu8qKA646SaLgizdzHH3LrV4TTVQs4njyIf8z
vX8Mg0vt8YdRbxqtTqFldyT21vy8tGLHb5F1gCBzFv2dBkq0fkYcWliK44lDTJ1/
kj2dBOFZR5yMvGS7x51Uv2hcZTZUxNDK4UuYOTkjaerpEhsKRFvvl4OAdKvMgV/y
fAMiNGrq/sG7dAdIs3iV8NZ6yA0rk2B8ncpfgiJieDZGNydD+vF1ofgFxC30oALc
aMkOajGBJEu3VUMy4qrZWNAU1k2voc/YxbOjXenmUKf3K/YZhMOL55FdXgAG3rAy
b+24+DLjQHePcoRWfd+cVPmevg3fCXkvXiC+Rr4N/v0+GJD5B0IBibZKrxbU+4+G
jU5S+pIV/5JuxQOV6Gwjtywv6FcDnx538UQZlM4IwJPQfjAc5y3CT5z2zZd76PN9
ZDSLAx2VFxbcJ4CRSTV7u2prqC/4WfVsQXHw1lcm5WdjNapgAgfcpysIqtxsi3LI
tewX8v6fsejjHBexD+9e9N57IYbcw49n17tXx1IlwphRjdNfXX0H7D78ZsdtuFuH
IXteP1lOqh1xDwPyqLCU7oofs61ztt5QWAomglhfhcXFtDh/b4ov/WYjuY5aDRtp
kbHFWkjyRFqw0/WiUmjqWS3que1OTVwN5+Lp2QyPSyIuqrqnPKAvpaP1ENTpqvzn
v5JhZgWb60yOxe2c1eYakLYIPw/PdVCqi69SmrWhQXUUVqlfrv7fi6Hr0bfLD1mf
CPiqoxd9oWac++FkjNFITJZXQkJ2OJSAN8yAUKf2OxVNR2zkubJQ40DdN7aJWYu1
vPAYTKLN5ez4Sp0b/WGOycWsD7Ks8U8ORB8zYXUInS2sFe++7EieYtmdmsHbgWGa
IVg0LrheBo45gl3N8gUprX7Dq+njU1oLWMBNV+myyUTM3X977tViythJr59w/WDk
oXT37MdfSoaRwmoIdhecq7lI9SCwX17Jm8PnSpB5vKtNdpARS7cCM7k3qV6QalpI
iKG0ZyXPY7bBIfqWKSdzeczB22l1F0b0FRgGpwkAIzulp43RPe2k0Z72bA+iICIQ
YMSjwMTe3ZHXr/IbKMBAM+kFxN11jAZBn5gdQ+ntOuSHJI4InqIBFXUzYGGqUmYc
XXnA/+qZpdJuhfWvRWQl9E1qfAvrEvnG/4ib4XCnPfH65wA3fvQ5VqLUJbD/AE+m
LGJA7Mm/whJS3VJWXL6LycK6fo66Mx21tagMzoIYQ/tLe83uUv+bk0nwa2dJUCo/
82fi9ZDc0ZA6zPPmcrWAXduZJZT14sBusyhZyEyxaIj3WJsgjSAeBvT5aPH7B2Zi
worMlDQwicUCdop84jDTv8cHJpHs85Aue65Ist9aY6oVRJlK6GetwHqRjuvIOo/s
ig9ktKasVDZ/QRjDpH5HLkhxtW0aE5/Zvui+MdIoTvc8kIF/1oA5jGRQwxUU+aqS
hoZpPN9TJuEXbofIOiSH5yd8i0UOGwTUOFUOG82fUT17CDD+SAn8e5BWVmOFwPpx
DyWYbqoIBkEVjjbDBIxKJM7SVLPEaq/DkUvXax4vO+EKql1cu4AL1iHyZH97iQEI
0zR6MAfbzOMo+5m14kc7ECBFT1ujKjFN4wLbmsvBgIKt2W6CkMfMuuwhjMyw7OxI
vrCowCn2ZdPRNHwhGIK5nsVZkXFoGDlJrn2Inh0xYufHw0H+x4ron1KM6Up9ecLm
JOUIprIT5AThvahHy/idcdH1KCb/+ip42xk0U4G708uU6/sAXQQG2vfxEl3BvTZG
YCu7E3OoMn9TASNvBZp9EfUhIzJYtUnnvzLQ46/JhZ0Ekd1psi/5164rUP0rVCOn
O2vml83GkZmfXhnvMMfjgtTtSo070Vxivf9E9IsB9AP+zzw/a+smpe0HsnM+ivjW
9KcBw2AY7dgvb8UX34pz5EcYga/Z6EgPr+FuqYDOOXi1acd2Z84a4ZWM7BkNc5sl
Zv/qFgFtFAJc1cL53UavOCwDoZwz2dDAEt0QInAXziEb8OPaR/kwQK6odLPo5Yt6
wk1ELpWn5NC2E8MZSof4j4b6bUusz1oCC+Ll1gGHN1g+pee3liCgeIFeBXMmAq2s
tRURs17q7oSxP4n1IMGVsYAsPayt/oaDKiWEfnphB0mj6W5Bc1Fpd0D7ei9AQTg4
m0bx/7B4dMGhJB/XmqeHAFywDS7jipZKAfnxUJgja6kPaIZy9teQANkRUrcbxoCo
wIp6JGzdLDlfVJBeu4qf2rWufQzE3F6I+7fFJ77fwO9sVr6a7wvhzTHV7Em1npRC
rSOpR2U5zdzswsdE45/wOIU3FmL+3AsGrsCmSH8eZnCBdEDDx0AgufaSJqv1Knnw
HUL5SvSceoTTSXa+FBAo2I6skYhrAmnqAyk7r8iS9x78fVEUJe+JRmsu7avNkUg8
sqWfE+INOycIe4JR1yyA2UnrMbJJjYNCiXDvQBa++1e471+nuHdMqQShUIlLDRjo
A9D8E2h4Wo7+BSSki/R3Qkj0Tt4f4yvK5mWdlQ9T1oqzPL0FkQ/ZfnVQY6QvIpFu
2ZJrbLkahqJwChKtQHMd0hRwCntdhRXkMc1P/0OZE7HpNGSSei89vYYDMG2G6f/C
KM/a9XlzQW4aPF6/2ifgeag1Z3IYQ+7ngqYh/j8hAwENyCsTqmxmFsKkih6O0B7z
lN6XyAiB80Ypz2uvOEUFozaNKU2AtlsN5fgoQZqKlUGUrUeXNCNi3bqXc+fEBvJq
PqHSfQqAyop19F3hS6cbkqay9G4d2TPc5QzrqUnYWxgBTjWl70LbntqLtPV/CCt4
GmjcOSLKsrPr4vX9ILR+Ne+HRAgNtr9dkGPnU3CAk4JRRgQIi95qFFkr3+dFmc4a
Y0+/TwGc1IgC6c4z2p1uTVI9FjPoO28UXQc9tcxoiykRzQzB5ZV/BbvG0KyXPNxI
gSjEOO0goCVaY+6aIwavh3hVED4lF+bj0gn2TLHQhd9jkSYGir9QHilcUvxMdDbS
g/DO0SudpGhTm9gw5JIFKr9Sqm/KkPfiOLkNkZKOQfUUQCIu4OgDc7lB7IC+tB+N
eysJpTIPnV2GekHN3TqALmP8xifssXe6B6mY4ZY/gRhY73pIMxcmvU5Fb3aVZEsS
vbWYvh7ZUGSMRP5swweNwlp2uEqsfeKnlxrMl4i6sFar25x6p16OAb3f1kQgFLJn
DBUqZsNrd9N2mkagl1ykcGzsPOMxP1zqmgZCpJAByRVNyuJbVn2pVuJssxBjwO1K
pdPFrajL5Z631YFEg7URIpQqD0cSgRzhNl9J5xilhmUqqR+rDEgAzttfHlzCu4OW
5bPlhDy1Sy4pNMLmfRDZB3AeOYTgTOGprIqtAGl2tv8pE0Gae2GKgKhx40xU5CZm
/DbeKAReI9GQ6Ys3b9cWeEe8bdCId8AGnZpjTq44xwMuRuZQP/ycdoT0G7Gw2sie
B7e/O93ULlyP4X5awE/7P5QP9YKtYi+2OJbMHN9kg3vuWF2U0oth8sEmoYzcTZW4
C/w5KQVQqBO+W6lxzVweYOSXggipL3GAWbdMm3Q14ts4mhROesqDZOunVO4TWorw
lStbBAWO1rZFPS1YpxBi5SkjnawMSJTqmRzkqnuCHuNOK1JRr+bs1BaPNCWD5JLh
D5ZTMZZvncxuyKpD8rW2XiUoVaU/rdXr1lqBHk/o3q3KX34mFDY4D66tqse3s97u
xn5Lp1QFc4y0hfwEaO9xgV8HDviAHegxFfVTs52jvnu9rL2oHyvBsC40jYJob+MB
HP2VT4ChI/jMNAAC/d9ZMbHIj+qVcaGpbbW3s6idI0XXgn9a3BMJu5HSDg19BHij
bSM8G4GSwyutH3kp4SaeoWPkFUxVDMU20gKJv2DpUDlmOba1b/d5w6tuYwK501RH
bLfMl3EiMi7aX/s1ko+p2z/bJhkVGDtfVVG2PFrlSSdk8+ONSOClmEeZvhlS4MzZ
Q3qMC8F6cscfOKUWKeIARVRcxjvZ4uzDN0Z3wQZ2aSE1AuwBNL86rzZ/XODVo2GZ
4l1Boj8vU5ncZ2oXij5oeSFynLe7XzHL6yip+FMqy//Si7zRV3VfzBr6vESH4lmN
fVhAxJoTLse2hA4q990KcPntteTmx7VTzLoEUkY164rOjy9U+kHznWwKh1oGrmHv
X/xqh9GNB2UFZYeqfC2rhu11RPr8S9+wrghtkQMn7WbC4PaVXuVYHO5rBOh5u9zt
OU1b0CMPpfHNc/yNh2AEGCm8vlV07uiq8d5h6iwoMukLs6srZeorOcjzgMYI2rOc
82aoxG20GFFuWIT8jd8wkFtS4F/zqkF/HUq+7Y1UcMC4wwaqSMB0sh7zo8vBW//f
FpdBA+s/B+S/WV1617H+Fi5a/WmlFkDWv9lbl8quE7+1wV/FihCkortmqgDsqw4v
nGjY88lpFrdbx4DsfSOYYNYypmux2uFi9UI1krZezlVKeivnGOfH6ERz+dqCGI3e
zI2ynmDiHNOVyqd/jDGCsNHiQrXGmi7EfRxLxPZw8pybf23EANY/3AvS+D/qEz9k
7pbpYVZkq4dDvaXSeXB2lDmMhMN44vEqCknFBK+dfWQ+ZbsUcYTAyiUulAq78uEs
6YL1Iwplqj3FXqwPrdwmpJQXMQfSulnMzm/rxkznX+yEQLBG1alef2vYjYZi5W/g
3nnE5jI54z1/G/QKVlS/fjPX19wqwIOegY70bgqHblGAzhC04a5XlK/C7egPegH7
PRKT70BptkgpvMCa1oQFGQeH7AFs2Ho6Mk/PQZm1/amRCMCb5sVzhjbKggSnrQ7G
Xl8YOeIcCkympQ5AV9cxtu2oM9BRBa8rUH5jKO5YhyUvZ6Hv7vELX8xCNb8DS0wr
BnYuk0b1pIKOlp1wUy+gYaMr6cKC3uywnIMeDa6N8UFbw2IIjRsdwgCFohdKWAYU
G9izkTsJ6ChxZNT6ouyS4wCELP//5PZpF14MgvUF87i2LHATW2/mKlp+CCHYLO3+
hPN5oErHkYkBq28fUpaAoexhibR3oK3rHUaHeu64UlAvKbvm10UYlz5d9nX23zIV
OxjRH1ehcmUpTcD0RtHv+T/ZuiOiEHs+wEGo+F7kN3WsVoTezexs49K5VXSolvg9
/5Tt+xRDjiSIZ99oP0v9P82DhHkwHbcZ7X1+uNHjWzS8Z88eMm0dVnSbHLxM8QJu
gS2fRlZFNW3TlUSLzbkMc8XsdzXmSRB6tC4zjalZXclP5FWSDIxAhPD32MhoVih0
g7Xlu3ohTxPBZpDOdFBdt3GL+ciHKghCcEw1ylcTagzH/9Vt7FCLAk7sTC9VNxPr
G7NOALfIv+6+aZjWLHFeGFpD86scT2Jr2LtIvs0QRvma4tCqo80dCSpBaQgXoW2W
veK9X5EZGTNLgTN/P2POcEnV5PuVsi/YI/k0KeccNOix29I7AuzCIAjT5wQDA9IW
0ut88wjMVbRl7IRq4Hq1z8az5qSc1RCkPUwgR4v69J3iO9YaKVEs4at5VikuN9py
5nSXGhjH/ncjnAJbiDUxH1LffKmwHsSel+BF1qdUrHuzmmpsxO5l+gQG+n4LhGrY
crIxZZI45/8Ab0x05B+GXbryjkhS1MPzfEe49JCBMrAOj0lO4fHxvl2GhDFWEJbC
kmrdrkp2crFxLPA1OF+rnt2nWCOQCWywU6gUbvQ9TDHN9/ygVZfJvLKqQorMSI2S
+OoDFbrZURrJid9leUc3PlyIoJhvDzXKW+RQs4+WqHEM3dFou5yFRl+PkgDCRXrP
h+ulwnytzhZ88om+WoUkf415EV09Jzvg4jEf1Qfet5+Ll5j277htFW+T6t/Bd9K/
nksIpyOK8lpkTTEeYbxlEWYiktVIMzSo3JHexbYztN6u/hsNaCu7OKsyU44fqPaB
PAga7MPQS4KaY8nC/fukAVOpLZM9evcDNGAR8nZU9bOWHnfbzPiHarVvOQRISo15
4CCRld0gzPT4cIFSKI7Sx5Dgp4W0UYGp9fCXLvCMdX6uO8vHcK/lNe6E7jbMzrmq
B6CkMPIEbKSxCdNDjQg5BcDbxOWFPG5wFu1PbMofv0H1dYI2/lPsQy3MbpvoRTxE
VlfjgN7HMQ92+we9Z9bOMtJAGpuDEwNO8yBCCa9xIIQMGtizfmsWsL03L16Pu6Pb
pQ5q0xZFCXEw8ct1dBoKOIJi29GMzBeNL/bKTZ+oVGudaKGYE1+Xawqck8H3t+lc
Q+/Zv4CtnB913+r2foNkClH7tSobsbBSpt2inhk9bt9VdUiDddKBnvosJryISNKr
pTo/xJ6z1ZHwR2nB+WvQHr3m6P2RB4it80I5O2X3GKHW8Vv7bK50aioz8020nwIb
oA2TK0ATWwrLHeujgH0knGsTj2kZ2hVpQTGaYW3171E3WQgLIXYBL4e6akJjCty6
RemPTEKvcxjuPEDWdmNahEJqPql3rdMo9un+XtIb4WK/rNqJlPlPJmErYaSaNU8Y
ew20x8at9OvOUIBQ5MbdbSvVgPLIWRUle2NAF+w5CTS/xxt1cZdZonJ71wE6Z9Rg
CRKNsX26lv91UVfTax8xEXrUnM895lzEqfjLMk8CekWKuhD+q0SgLXNVeO471rSV
EQeJHyO+VJAyao0H2QeMxKWQey9EuNQ4qhG3vQPDE52uNaLL0m/K//uVHq6tmuTF
ttzBXYAhU+PQEllX+0GHtfHBjzcRGPSar0wO8H3oMM/dfdTy6FwXh3/1FgqDxogw
/SDakbV3NS2Ke/BUulPvh7l3xh1LA3WhqRx46lCXKwiMTUNiQ78F5i9u1Zvo3s6m
M6k5UjxSeUfaw2t/WYSn0rJ6R8Gb8LAQzst1ckvqBJabA7W+pw7euF6utqK8hOfE
s7zBkRqT+Cse78ZTeIJa+pZbluVQiliQpnxG8l7qg3FqmxcbqpJKmwolCjsUlSsL
ARa7QjFOXuDWcvkjA9BBxZVHRJje6VWKoJs2xK9O/gLINIvtV5OFOov82PlrhLpD
fomQN8qKIROclCXIl8+kS71vdqf/ep3iJ/DWw0AngXGdDGczFiE98aUQ1F2jEwn2
0XR5uzgMz3FusFXv6AAzmevbahkBXXkhS8GVI9ugjzpGQZdd3WIedkXqY1zwLxcl
LRDoPgxaubH6gThHK/HNV5I5MHxO1x0eot6TDR61TpNVhqnoIPaYLX0TYut+poRI
1uJ99JRzZQuxJ0JwEy7O1BZmSlQQUFdTwxv+pRVtjBNkRyo/tcPM57Ik0p1NYhcq
mRw2cFLRu/3Z3PpvaBPdESSEHV95nZhifim+LirxEhrvAbHxw0CozEHQowdNULtt
XRkPDeRb4tT+6/SC77TO44iGGAOUARfQpShOpkpKJnX4QU9h1jpmZL1tDQh0yiY1
nEPlrPL3fE7xtOQqo8fK56ZXRKNFyFwQKl+D0rHQfIJawTdTsZ/MQu3tPD9uiNJB
rid5d2zzJk9DNZQyiq2WOcOb/WhdMlWq9lzBPjAiunwAAEjAuEw3oFwkqzROWYLQ
9X0L86JK0P6BS1H26W8S9TYB6o5RHq/k53ge9pNkIkaPB3cAqCPKdcMpAFkO1EEa
vXKNmx6bZGI3lzQF4Tin7T5u3f3YjmTfTPH28lLIZGUXQhPBU9cRb395Mgs7lKu9
8FNR2ZQ7OfNX90SQT4ZOapA/NQEP2Lc7/RcBW9bglMcJa5lfx4XyNJ5VM6ZdfjNd
xbhlqhWJtzT+Ed1+/2k6W7lazNCUFWCIL1FY3FKy6WSmYuOLYl7Z4dgx8L8yycuk
OYFwX5I9TAPfNh51UL7wgmUfOKigyk3VGXmSgL93CqFbmHRns2BXSkaAIIVMTYhI
mMbFQh64QHCswYt9MB9WkDhGPVirHyBmfN+dn7tNyh8dXB7MpXW5LiRd871tNkEN
OLM3biDQC55P8Q1Od4WaOIobT34Y41fStxiu65zUv+lxDY/grNP0xtsWUOFeO286
r3BJWWMADNHXWaJGTEIhPpUF3pr2yhN79zEMuJur7y1WtFjJjWmbQRyq6yaZlyhC
988OMoLWhxZuLnb41Pq5R7t0xa+fSEUIeaviaPQxMv04+QJBeaodVIrQY36xwfdy
Q/FkCc/vMGVWuyqfq1/ZAyFIIngsnpr2du/kl8oadSIB2Bq4FJHnPIkx9VvHhiPC
N7QLyzGEUeXvtfRj7G6eTwcZmfqmxF1p0GCstNH/YAdyH9CGd/O6ly1AR5X2adng
SEe/moslPZJHZ8tzMhs/XlkL42CyGOGu+JclTDxsAdEGxiEbIm8FCMNsrvXuanAL
tJGpvJDzTfIozAR4F8yzJgnOJpCy/v/b51wwqislUuFTPwFpglHIVOdg5bZgr3bI
lxYKO3ZrmYtz75JYe/bgAeFVM3hPvXpkCrU982BNrAOo4/zoYfrILWHKrs/IOBjJ
IBep8J+mcP1WVWMm9mHwGwuVQa3Xv5i/HrXDlO9tAOtmlwdjSh0H5oi+K/PqfdO+
D9KUtn+qSVWmflEG94CEzICtVllTk/aIPNUnqPmxJG3wmxZOh96hWUqhYVtiYLKv
se6ycCg7PP+sXhP6er/sPNBS3vJHXg6LENHcGesocr0kk+dyq7PRsShLaXWc7q8H
fMBo0hfXHpFBFYB7+Ps4i2d0AMS0ZHUCQ+2aBTe2R2XdR7xo6pwaD6hmDShHctja
ofc4TOyNh5/L6P5V2o6TM1eIjBWEd6qMxZr5O90BXwjRcp7CqfnXZZdLM8YRp2Om
v2rGMjsoNdQKistpn5I/yAsStFViD4YatSbIj6SU0ny83hQDemBbOk1+Np0+RFR6
py09dLjyTRnKqT3nWqeHKUu4kRG2aLSHH14WXAXs9KXErv2p+1wreQOS9y+lT2c/
NvO+mRkND215ukzlY9wqReOFbLTlfnWqL3FhYUMoji10V7mUlVV4I1Nln7jodPTK
aTHlLrZ9MYzdRrRYvCpi0Q+5X3jRJVEAX1TcVVMVJdVdLQvP6yHz7WEDzH32vYWI
kRsH0U3JIEvAmYmwSwFgGl/LoPWX/UZk9h4VMYoFgPhmwTe6iVwWdgEOSiezGSk3
VDwNQgdByv2OEC1H2dMTowzsGFOKvXis+9159YV8QqH+hg92ozxru275nhI0L+fK
pew9P5St2oABQ+HREBcpSXBmsQGyC0ELAoXB//yDtg8foH9F/pB6IWITBcFSQPhq
lknuwsOmOd1ldzM9Ji9Aug81smcfoRwyo+vwcaNCvopdkQ7gjKVsM6vrS2kjhIBe
YVSHfNSTm1CAMsgtGrG547Bf8TE/Ac4xQSWE3TwUPxx7hg/EX+EVL/XL7SMJ7loA
nzQuJ4xWnE/A6MCdTo22Ob5O+Q0hEswx/01EHC/R98nkiq6MR5lNMz+I5iPbUnFz
Fe/Uht44IL3pjCHBLD3Bg0lh9zt0EndpvKkl1UIb+Ljr1iYQxCJZsSW2rrzHOQhD
Pt8jKz6h5G+ALgEy748T4ezfXwjgha0WGGdrQ4ezm9B7AUe734zvVJOFqXClhbKR
z1hnVzvLa3bSBFhD/eXlOAelgZcnhTv0Hwztt3hpZSphp5LzxogXZFLUJ0rHn03h
x26YmWarxpDUifbwU4/jBSjhv+1R+7zvCQRPoNw2p82igJ8ebY0AXbHOBxQACXWF
XUwe9+B5DmOgpTyl+2CS4YGKql6tOwZnxTMghj06fXzBV6EHKmFUknmVBkoCaSM/
V5xkQCLMk41lh7r4HE37Ew/2S90rFoIUatL+UDboIHVF3gQ6uOyc6wi2LE6AspUD
0Lv46n8V60Euv+5uHJY6jis3yD13Go9MwAAybDwHxoczYDHKWW0sQteaE96G1Ilg
zt+/x5S92LqlDZzhEIvnUMnFiIAi/4MWMRE0Up7D3DLdWVsQkB/LX09Lm2ciPnyx
iPdBhdPviC/9pFENG/MVmshW+lsX4HOuAB83zaMXLXTozQw3C/ILmHGLMPa0PntF
kqZunIH32FKe3OkaCdoBpHTyav+agcMTsjDYMSuNyEtAlwpmp13xxZEwEity2zq0
kODk9rcnSeRKP249OEmprtOjTAVnQruzS9eQ8sNDq7GYF0PrYnathhWf5fbK1wf7
1MNb6J0waKvV6QKocCRJMGHMbI0OZKqRUHoWDalCb8kKHzt5OTcll79T6RhPGPA0
GC3gMVLIDIeGs3ilxWISzxoxqE5ArICoi5Q156Z5Y+HguUOqKcbn0Q/uB/DKoYu0
wTugNRh+AvBnnO5Ws/FoYaNvP+VOH02LmRzgPJcAf15reFpY3XpDLl81bpWl3W2h
hlYFQSs3Karxxu4zhPChHfVz8dYUKQJ9Jgxar2K6EsPQ8ygObn6TKfzfpzsiM2jE
SszYvfAPt1hWWj1+o6HE/FVn6vgy+MZl0r0Tvi3FgUtGj+PaRsPYpkrXEKodt7qV
1hmrCgLh47ISiO6TSa5qUmVgpZdE1MoljQVv+lICt8eb5pJXZOYz402a2j6x7bI0
YzjbTcf5A+EQlOkBxKZ28rWi7+yiDPtHulUrhv9b0Gp1OjL0cI6GPLZ9zRlC3d5b
Im5o71D1cmzf+V5j5tddU5fxIAX/JcYvgi8dDFfjkNFnojQjrewHQxUHwyiziaSQ
8gQpJaeehwBsQnx1uVI12dIy+O1MtZqvPgnrgiHHvr28CBqSOFhUUG1XaoYXKQGB
j7+UHaDCvel2jVPjJ0gTwR0sSK4LGobROrSknoHRHiNQgUYBsSVr2gw0wDzb+e2m
6aX02bSlDhbqw4jdIPO1CKUxoaE6lPa6Mb+uDeG5JUdiUmtpvLt3i9vV7QbVgsC9
EC8eqaoMkoTnZob0R0MqmucW4SKK6mZ88Pl2038JFhcMFe80OOfJf6aileh+ZA7Z
bjb5DW+nLQ/+Q6xA58zJ7jIyQeJ/3eNOaFC6f/w7W41yDw2gBwyOVfzmp/t/0cE7
W3qkcNaBEGz7epn1tcFvk/+WDz8a3RagYqEcR/GztgDqCZIVZSNwei4VxAiYy/2b
O7Knvj9iYXp8zQwiDwGnDgWaNlXOYkcpTgLePaiqeQp0i6zlQgTaeR+ztzNWPXtn
UnJjqS1AF+FFiBkB7Hni6GlaPbc7l1jqPMHI81sLUuhj9gAHWHUWqs8HFMJ23WVn
cT4IYgNbFfXQroJ+KvZ2GRo2Vp2qJeKBInhIgcDf9Ul8AIv3SmptqH731LcRDT+f
WUBN+IKcXVjVK8c480VaSMwC0wTwNrZTQGLHNFTBcT3fYpKDePmYJpEsjn4pqu+/
dhGccQKMK8NgeAVXyN87ogktjQnlxfrsNDRdGaZ3bJA0aHkDJLbVC4GTSnafP/of
LEFEr5AvA1JoNmf9sBrUEKuweUiK8JmQVSr72/2XowUr8eI2KVT4VVpJ+hy36uPe
H3T4AfmPLcCGx3WKYro4tMHIJ5insQ8uQKmEC/BrpODSYpmJCiLRv+gSk5+N2u/e
YtbHG0m3VNmXXUa/d2n5iM4Lh+EtbYj4IKzl5fS2wt/LLIEOZ2B0odKxGNyBj7MR
mW0PmU11gC81j/xJoirDOJo3cjv1rF9VrMhwCqouIhcJ04rPO/YY0ayzXclTf3K/
lzcoP+VViBAPrxWKaiOXkUJKydTTn7dYsssN4jhpQh/GCMP8I53H/Re7d5Pd7N3Q
+VoQdxH9+dJiX/tjQn2/m+Q4uo/vyEPqyk0z6/SLZsd1tq1hRyL4EGNSL/pGSqE9
ftTHGXoRGaFHz9eNtsL92swMBUb7wOLCRYrF8hyktyWKP7loch6exUjP9E6KweKW
aPkupsVN9TnMi71KhvloxOOIsYIqXV/e/m/FLkpX3vODo+LKX7uxfqt0sy3XZ389
zqmOX8hcCuEVnGBhvzXyDz3FGyVkujxL64ZUxbhiwwoh9bq5PYfihHo3WXqLyy+q
P5JLimWv1Kl/NfrkbqYUk0/h7lzw2YfdybQciachEpVl0MJRwuFvU+6IaDgvDcJJ
lPY2WSfW7gMfiXyokqwlx+mlWQ2blyv3XV7yfi5468fZAEmJw6+GxqQM/JLAEuWi
bFqm9kej0Wi7AtKziOo/zNXw5WT2RknCWzr/MpN0XnwSTFFIUliXuDD0ApWtmkcI
/5jnpybi/jGIrfX/qsccdksJWMI1kBW3Jd+lCYCZ5Ohy3fUc2pyuPsdL0ZU2gzKA
yMXc1Mz3Y9UTcpouqgvZkuSGWJrUhMbe2/hoFDpkLNn+tR21KPQL+uGJAqB/kCPZ
r+g2iEPJ6XgV0g21u9pJlYlWfjITZI9J6BS9wfekZk4TWc/IFhSILkH0U2gOaBrB
neyTso6Umkvf9tMyQL6oeT3O0Tn4QLpgAqnrV+seyHgk8dWQ7heFkzJ5Yl6egFjd
U3uwYP/5NboaRga/d+mG1v88yKK7xNANOECIzH4rdK6FRbIo/2kOngVBbv7Dakd1
B5L/4qgQI/NFU4KVwqgPybUToGQhqG8K0Ch3/0jw6pMrLNA0u5FOMq+7QDaUIN5c
JNLQ0WKAWS3uUWw0ufAb7IKNngjLtQ00WdvWggCVaSlQA8c8YJbGRJjbDXZssd9m
NG35x8knqMqVXsw+RZCOyLvUmoLox48ezoyIGmK2waAKLmv7gPpJNLbcACxALBWL
JH4y2YKIDhQH3KHftlyFHIUt62BJr7pO0rNmous4+iPVj8+XWtO5Ux+qbjV+oFfJ
Px+9489zKQSsHhzelv2PboUjI2l767v/D2tF5Eti4GI6ldFyVSkW1HYV6Tky/49+
XHnZBE2zMa7/zB+I6Xpce332EDlyfMmJbl6HLD5A+JXU7/EIy+s9EKvxutNFb/WJ
xOUstvvyJgfv8zUGWzav0afi2W2lF5XIK8JhrckaanPVnaZG+XImejN1Iew/fDQU
CHlaZ2RvFAqsXLrN+1mPPLELIi81Aqgpwj8X1MFbGGOvfNU34lSkfb3BHtRF+7Ja
74ZXxL4iVl0oC/pxnwwtankFT79gsjsiSrmVKNK9T8WZgZrTI+j3vGfkGXtQOnXL
HgRPF7djxbznTotUwBgO3GcW7WNuFu0mNCGmgVMa1T/ddquQQOKT/nxqI9P50E6l
TOjFyIU/Gl123IOShB1pW0EEliZjc3RdT7Uk1IzqOyx7iJpBmvTduLMbQ9eF1NhT
aJrL1JfaQGSxvfsQfvx5id6kIlY4JvHihaAQ5A/7zzg7Bvadu8wZYZzIbD9qGbGt
nLtI9cfxFlxvmU/yt8m7Z4ZtzjDqihwRvEb9Zy91fKmY5sfH0qCZPgVyHiuBuyVH
PbN4m4Uq3q4NxJytkzF7CRWee+fnIwJIS4eSQNJWx7dRWLwAPQvKbi8t2HZjNslT
mxB7vXPK7Ib6NzzzBQlfuLNF1zWxUAQV78MZz3wM7+W0NKozFTgXbmdHUVWkpPMT
gMjqO6GouiojidWQTzWQrdo3Fst6yGUZxMG08E2l7nyIdwaN3cIE8+HIhqEXbx4/
571CDe7br9t43g72i9Q2KFi1dR9IWvJGNE2klDiYctIbN9n4b3iba1OeU7BfEh72
+Ryrc1tvlIDnHvuTs7uHZEbfMP8kGA33/rGNSuMNdRsuQI8mEAgjaAYXJQKgfSZh
3HNUdA775L8eIJnvW6dIYYD72LNRVjw2fXUdo++M1+6zCSUqUOqpqcSW07D0qevL
SGOQbNZINL8pigamYs3Qf7HalA9BR0Kxtz1SMlQ1oRRg1DIVa/dWXsW1H+x4nY+w
TnisuOh+UOHWJ31JEw5+M5tscNYxLCDr0msHlMwjX3GOpO+3wDMWUWMJeGLYk5WP
3HJpQJM6b6YlQRjFX4G0u73eVkr6Ho0L4xMhtL46M0TfUQdcwRxFhdTQR/tsRGfL
9zgR3mcygnfGbk4Fy3xyOZaT2EzU9KRYaLlrZ3camM8Z+MjHEOBKlXpXLSnuzpja
SSzqMehvzEGG0cMMOogW1Qk2NjZPv+qOaxiGs9oYtuNmWIWnO6+HmEghJJXZR3V3
uZbsQVdPwtSuFwAprZxX490q47kV9rGS6qE3+zcdlbHY3KHD8Le+wFUGRStOseme
mVKQj2GVtXdVT6gf7ipkYf+uR1bvpEzm8fu1ct+qJLaOdB5u3z1qAqQUlKRunw5q
2yeWPHUPU9+upGwqtOn2TozbTfQ57GlAaHCUf0hmvPq3MN7NEGH8KjYkVfPxJQSL
ivU+IaTq3VhCYjqP0m54kPkLsXv+oO9t6xS4wAoXxZLOlUD1c7cqAVvN2ezNOtia
9lcBValEi1qc/eyLYN4d7XnOxyy06Hj6IUeYtRY4AuX0BLGW5SuRMiPqsmkm1pj4
sjNP/R8vTXKM+D9e3LhKcRY3hiq5tsczNea8yyDit6iulBIMm76A/lf9gl1UpQJk
7Au8JC5uHG4I6wvTpRh9ih6OMGXI8ZRuRM+GeUtkzA7GZDkAwdRLQ5Dr81Bgwhdz
W915jP+ZBTvr8rB7KtA170cqseBn5j89zXghchhJxhcN5tZszqKOzMQ3eWv6X2Dm
UBVGAj0GqxqWfZymV6vfaOWVLggIftCSAqoT1WD/cJe/usyzu+B7Rw//k3GlKj1G
bmuLe8gtbOJnMXkCHd18voreCpQVNqVQreJaRWLNNn/Iy5Ajxm3dCS0oHFWFLSfK
5CUPe3WZuK9iIAS1CcUBUE+1USJzr72qWpAv4XNghs0+XqfZZuqgDGZocpEHz/o0
s2BS5T4Z57jZkrquRPJPIJY9d5aF6KyFkJUgxMuaBBnzt9ctfthyzGEt1fHCQQFk
rXYGrcj2VPLTE2UXA4pEM/RYmO4+VYiyzWuXcr9ZQNmn9iRIF5p3r3UcLp2cTOks
q79/skYnwkOPdTl8nPKlDkIT7Lc+wMvDLp7TKNNOMbeCgeqQjfMzS31lSZbeKKXm
i2wUjOcFOChjvToyiTo5s+PWSl06wsUvdeqmjvqF+OCcPYgXqXWCLz6aD7wejdz3
rUHIy8agxXBYPj7oL+TljWkbt6OJ0s55Buwnbe4dGSXke9b2kp4J/z2LDGoGfVWN
bSlx45QXzowIt3QKatsXIIk3/R/Y1h2dIi+jL3klma0b1x8B+LUaEZBznoS+LGxv
35sB5O9+RsFFva+ZPyfLinuMcmEO3gzWCO8povPDo4Lq5j/0nP2VzIDn1uSQ2yQm
ZLOpNKAIAxAAUhXWCVXrwkSgZ04mvmwx6XkR8p5kMsuKFb/WNTdNKZTE5P/j9Obr
U4q5B4XDF21kM9oxyI7t8umZrYQC6rTwNvRbGZAiJx2Rz7aNPelfzH8pxMXRPq9D
o6PMCLAZAGRLbmKmAeKuoZ4ow1P5c1sWbGioSnxwfWfKhnUzofBmDH4/ctTo9skH
fuOEhANm04lBh7WPNS7Ia0krpQQNy/J3V716QzijYSwEgJ28E7edn84ThN3MB8En
anX6YcXs/yMe03H24Uvz8RY7ap6GlUEozT23N7T5cZ6DQNguEXZbWX8+Zmc0WW34
Z7WPZ7IWvkugxdRT0bSp/xqieLaCXcdWhs36gw/v/JpOUkr92hhHkNVywSL36jOy
XZw08TucZZRnNx1p44VO35nSXN2TCJZnqsQ2W5paEjlFIvYwI4XD/anRdqqD5a+U
vGAYZvESeFs/83B2kxR8K5nrtZbUvFW3MDJ+ROO0jSYsgR7qHUkMrwV8lsmVwwhR
BPRntEvni2RNpcibMkeBywyJNNg6stp2bh1wj/68D2QeYm0eGHgt0Dh0jjKEEjPu
XoR1Zjh3Wc+CPw+SIWANGYYWTTD14vd/ZKcQ+00TL3wbRg/6AYxLO+8O7Urlnr8h
JjdI+U7n9//VPgh5YUxtxnUSU+DajFWi+WmdNMmLgI5+VlYa30U++flCIrCmRv3C
MC1yMez8EIz7aR9zz1Q9rErzNo2t/0CfJQgIcIoL6MFm0wwwIvjBBe7bZ3v/bhgE
29ikt4bOTDD5SGd2UjNVAF6kNSXls7fIIeddi5SboFaiV0iPo4POM7dDo5LxZ8gN
JYyaEiTohw6fATJQ2Vw9B+eWJE2j2X12j7vFUTvKfhsEu4vyUOmMCIrODwDWSd0H
YhB/siFXzOnY3yeVejE4ifgbkQTnSJUv3Wi7E/Ne3fBA5GoZIkweJAPQGIvRVdUz
OkzHsdo8LrPpc3mcrhX51RGnokNcWkjMJyQdIRatxYCXHKsWgPyJ0Q+L+boGs19y
Yox7CShVzkTxQw8IhGAI4vYj9u73ZKEE4FRsOa1DycBV7E8nhXpUQ2Bi4U6FZ6Z1
j4MaPc8x5MFyj3FAPJUfcqFe9vWxEGFbSPkuqKrwp9MFcUCgdqXjuBwjpnTfNH3w
+iWVdq0XYqFA48RxMci/bYZRr9fpyGuENM00gBDnH0KVSnKqRaLlfehnPQYOfRma
7xpYq0ibf9yBUcSejjiUxsEWao9abs1qETDb6JxixL02JuQ2Rptu9Sd2CQ+aZNNJ
h46DQN52CEoKXLYXpJGWz6d5jkme8uEU0btsufc44CL2FvydAaaHKa51giVmOKsr
1kgI6SSYs4g6xGCvDmbcOCcWfmB8AuDAonZjzLk89bkt3kwFuTCLL4UciQLpau9W
8F3Q/FMTRti0UyThPYCaQzaypGQmo1QoVnDs7pv3aOqfmrDLb3LbrykEJxzJ8Ldj
pARPLgMloKuddFpOxPTxIP599R/t/TH8tyfxakLC7sI/WyoS2+F+MWYp7JdZc2iq
zcEAzzjsupuzrTUfTogDeippvllrCzOH90TC5CYigfbOAaJtZRv2kz08Z6YwsrJh
j61NCxDTo0D7PqId0gaLtv3DMCMykrzMrJI1KTcFNbm15KbNVV+QxN9lphYmXoHI
to0UNvj3V3OS3v+gPs1S5r2b0WmeOhqp+82Fk38zJVtkQtws5thLbJ6rpi0nl+Tv
vkzR+ti4GpamtM0p7mpOsRLHIi4m+OA5+Lcu83mXmc66ivo4K4ja4YKx9gE1GqwQ
h4mbF+rgFfv1zJnqGN3yCkADITDoqi80wR1cQ2bAsPWKN2AvJsM04K6Ja8jkcCVW
S4vIOTVQwXeu5jv84uSHkhHSl4wme0XZiqvdk3sdUEeeakcR474tnCnTtas6DlXc
G3FTewQofBu7GauMOld65nfLdCWUWfyjNZKjBR14etcbRSxue1tcKCdQNVkQteAT
psqr35JwnhrBXPEwGYIwsSXFgw6XWwBTqo543bG4YWYcDqh5y+iZWubSbi2BRA4/
ZL230ZiM5IwlX3KM12e0AbgRfjfHyMkVCIJEtk+STU34Txlo29LKKnSg/LfWyMtm
XkYTn1sFdzpbCHBS4qyNqd5Zaw7vZa2KM+uW1cM8YoBxEzPWToqvarMzfaReF4AO
/1CMWR/qbfPSQf81fr+x2BuHn5d7de5WwCbBQd8R+5MhellBLtpMnECjGRCtI3ll
fQRBy9eRapzHgXcQhMyQFSPhRgaJK5o6YIMLZ23X7LFjJrBSLCXXQmn2ccLpJwos
iur4eETnPe3xpNV6BuQ05C/XWMpj4LapMk6CsCt7Xx/Z71wCijzf3FhhyiVuuBdo
Htldpt9/aAV0Pj1juOsUXbbbAxousHsutjsIRnuFBBFOLW+33C2pt0JrMZsuGOCy
lUUWAJBRRV4jVkyCni68iCxOFeDKR6j+7B94wPxNSfyZM6DuiHHtR5RkFoOG+JKU
qEEkXzyA5doK0ONCuYaTLPohXh3imTE7aIt1YY064Vm4u5nMsyPB26TKNeC1FsMc
hYatamQmkRjmmC48bAiz6WoamRY/J691EZ+rw361BFVAlMhLtyY1Szhw00OXsm+V
2ddJaFW0bycgLss0Ze8AJnRENzqhXo8pG0f+tXlZMmMBlpYam2+20jvUVN43SPth
3CXLgZtcRqhOh7FV2/xJ0vdUGXWAl4oe5gyOXPAOniUBWXyBFcjJfxCS+g6/0gEB
e3JVD415/J8qnjdoCk/MO8UW37uDkIV0ZZ2sY7I4eHGvh+6IpBhahAhTbtQdYtbt
SxMRwj2jWTYfe7w7nN7YEa2xyjDuhNgwcj0aHnXNQ6moZudmacAFvWZm9sezxJcO
vK+FI32Yej0xMERzAuUOlUzExTL95wI2YqE5pbem2wvvwTY+Gh2X4BXqZTcxzUcd
3QHB+L4P755t7APIIzpg4TEZeju2HKwjFz7WZACRKtjZV4H0iT1VsAawfEesa7ZY
umr3KnqjCEk5vuWG7jnZxyGI1KybtRojJf3Q0wwkrfKst5cvKV0MDxj5ACQZ4hwm
ZzPgB0PXP7O797nZtkI8F7sb02/5dgsExV2ULunNj6E46GcxXp3jnS2ZJ7AaEHKE
APZ4WoEM9F6hWBsOLw9o0gw3Ei2MrC43QWD9HLH257k4m7R5KZy1rfPnNAqLClhZ
W9ZwidOmDvP+K8dRepLSIwpWWNw2KBuoxvVXhAZh9IKmBYIxj+B8aXPI7cA42QjN
0CYZk460KTTpMLl9CPVWXP7itSjlWj6wLTOisFgTYNUhKikAI63gUqyg3ixId+s0
0gBfn0RekRgJYvqsCkN/5toqWkGKHRWAwPhUlBao4EIRom3CiW48OeZ0XOboIah/
QmtUQcVQ9cmRICmWxhj8iQkk2yb+36Q6tulTwv2BsBtWJ8pwXpTr4auAk94ZRDd+
eaQLwItaAphNzARLTkGsojskbRFQcaje3QokXG3IYY91RcfVwP0tjP1QaUIeKwgU
8L+Ufbs8SLmS2j0vhbmV1xEmchihP2x/+TgYERaN8989UiWdUakHlF73yYNfVuO9
nIHpiB3y7mKd0UQg40sdLeu2QEn/avL7ERXRgflQXXm3tFQwbP8nsrR0fk5iITbw
abRRXUJfiWaO9pb0Nd9e+5pZRjy5EtG7fqshFRMhLB9TmYYNGzyNLREgTs3sEB9g
PM1d2O0tWvTmwl1kcDjvUAUb2PLcCpUq15Cmz6HOyU3LCTw4+hha+flVGVDneLct
joRWsRxSSNEQxSlfBTf04ztCCX6o4D9pah0ilbbHTd9u5nBgIzMP9GcEx74PVlIP
ttTnmHZaudwJR9HIIAx6zofGrg5z3TZSA/TMLzVVsrdnj5r50F6PHvCcMOvGD7jA
74wkLe3GprcQtn0b95PDib+wvoZJxH8nsV46GCyWMmAPn9Ir9qgArZnJVeeGDvhQ
seons4Gn6xcxRIEAVoKKeCUpzWitLGKK0UcDQ/tJLxTMyeVHUp3RompefUYv/9Gd
C4waQk8CdczG0Elvl0qNpnn0krM8xjuU8/sMDZ4HWrlCU5aPX9xeFStoQ2LxPdXo
S3m5WymqHq266gyMSjTQFaN3vOeJLXh1NtbQRFeEIYF8xwwNgDGwwKBBFtr87SsV
DhiLE02rKSLmHsDci4GF+WWvQNKpV93QT+nut7SdluVGWGssrKOrA2BeoXeG2usM
n3BBwK2dq4yIABRMy0QzgR0PsVYrTV7XwpvO1BMSbwe09e5dgAszAM4kVy7Q8jWh
5vGNfhjXay7c3Ol9iPGIeAdXQwyiC0SSmDpAx7jc5nMEjwO25tOKrqNxy3EMuuwu
PTu7QOvSIM0uKb3jCU4MnfNjsZ4bOTDPH9YEFzHO6JHLr8yG7L8sKMUFyv1p4RN+
oIYbnLPWSJBMwZDa6K4zRuZA+q+GIC9NP5aaZOocsU6FkgC8bRkf3bYFQV/+hzxY
hpz1Tt0MmfqzMDBiNNJ3zui7gTqQ3TM2IVRQzQvlPfpEfnFs0sQtac7Q4dQ5DpIM
RpZveWOsfONw1o3UJgjQwiEqWs41IsWKTR295HJAmQsIoqQ0SjHw+auwO11u//Ir
zCuMR2gv5uEsJok37mKMqQqTwMic0rCk0g3YpYX44gIT43heZLZpLytrcMyXzyIF
TEwEc2Ogo840JjpGCoLjrZwmqJs1/QSofj/km35ZD8g+fAa9PETnqmsjcO28L3i4
oh/V7nTzu+mDD87hXBA8sw2JYlVHjXl4AJiY8Ovjhfmxw6r0AOkLUEopOaupFdJg
fJLLSWqpHCHCepefbT8pP2grnrc9q1ZmN8vYV3JMqOYfv/lK3xkxCIM20tEoKqs/
y64EMRyHgcIhddl8YzzwJKnwHB6WIRGe4jeXgUbMPJERbPcgsD07IVVIWno3ecEP
GkisTHAq3vt1JQbjMRP6/ZzpY/jwHfmfewMZRfxpbXCJ40zqcM/IkbwnLMN8BRQe
EAyebBw+AetTfNFab7yezX7VKRiT6Pnb2Fm2R+5ucXiKThIE7fC6aL5KcEkJvtZQ
7xH4ckneKe3A7snmuEK+Y07kh1rhQAfNxtHytFZD2PyEleXiLXSvlqqxGOl/eu41
OHx1lE0BEHg9W5BXelk28oiRFr4B2sfSVznAfeQydjW5BnjgpWt8/h4LRBSlVvFI
U5hW1yZ+NEvO/pb9eOavvWaeeGCU6UmaZHpCZvm+nzvwXRlX19HbRVtkHOIOwH38
JMguQ0+BQ8KOh8WjWlKoD83SEbcJVLQZ+agdc69XTHPdjVYYlVj2A0ORkVpy9HVc
k9ydes3MgHrzwlf2NQgjpXSBvCCpA9TVg3s5R1516PgPgqiFkwl+2pa2pR8rHW1x
k297sNijUVfow7sgTtHr+4vM+I9tNwSocKyqpewt0B61ySa4svCD4EkzRbSF4HH0
FtqsTJlhKg8H+RV1mrODwUUdEWy7ByoSjCWuzXkTWMcJR4cGQz4G8lQjCWnJARWi
IcH6imZ7GjmWFrS9Edi4Ad4b7/kPCh87rTrgaVuebK8IOLLRoWsddDgrOCF0iPmg
hvzt76T6XXTzoa7q+tb1XLLxwTMjJcCFo2oVFPjCbOTfMUbGXLWlMmVfCURbWbwE
zvLm3lRzM7mQaxfQNYR3lcOAQlKtizBRQcOX1nm6BXPiPzUtaeXWmbC2V6DiR40f
t9rI/zThyWhhngyV4Duz5zRf4V9DMyPxDjzpHKFV7JRcJQLpUqLESNZO0VmCRyjQ
ySQbDZO2uqMcDiT7oArj5iV8CoyW9/WsgUIYG0hKqxZTcFVufWosB0N8QkR3r+o5
EHE2JVnsrn1ad+KXLZ1A0MKoOYYDr5yEX/ALAZV2Jp4S2UzFavJ8/q4HJYT54kGp
Oi9Ty4m8zzP5IP8TQ8rwWO6wyniTavx40tb6i/xJRoQAW2cdOdRAndPm2gWenP0Q
BJMNaf5EhUQDi8bd2bjdysHm+sK3cjukSXYpSnMbNX6+0GySHvOAI6lBD6GjPOj0
sCuHO1WrnstAD6Tz6yG0430DfgK5itbsVXqFWY2I+8xLkIKrUpfCvwH11iL5xbLz
OGYwSM8ShumdSo8NW4Mtm9FQ+JThrx6z7TIZI+c2TbdKUaw73VIUuBhUd9cIu/83
haorh1p4C5uRgbfvtu0hrSucsv+OAejMAHbf22MWKHJcvNwrYmJTaKcbtJiC54Qi
jSh/KgdslKTyUZxDziFxm/jtzrRmi15GqGLEoiw/mE1VDGhTXZcJqygCds94kSZy
MZYvggBZn07pHir509BPQqZsZ+6ttt+/DJDoMT67F/vo/hVPn5Q+Q41ajOpZIvNP
98AuTikXtfEO+nVPBhK+x58/ItX0wGodp5M0AxggpJAiKEPSNZyRK1CN60wLiLyT
t9+aMx7f/IUjswbRBRp9LWv0L9aTynOD62wWXia8UVm7n4XUofdN122GM20x0Yco
wq/CYuK4B/aI9BUIvTGLz/R+mCNz/DZUGB9znNU9b0pudC/tzpoQ1iJGjzKLIYBH
IEpk/m8UGEHP0b3h+Ww04XrgNJuedzaQ3/Ptwm3QAU6wyPvaX0BvbBf2kE6N3lMW
1hOutt6Hmpr0tisJcXSsdhh/mSPiy9bpY9xZrqpOImhZgmyhDxwZyNVrk/V4sqZ5
QE8a4Hue77hh6PAhhWeYl7RA4iYf827uuWcqeOqXS6Jc9HGCXQo7k/gb7BoIBS2L
Hv/FOdhREDm7hTFA3SfRt806yviRlyJKEtieDyY6HdIB8jLfZ+rauJkQqXhqEPTD
68wA2G36w4yTJEkqmqXX6Yu6eVtEjVrSum51amnW7psiOB+GO7O93VS6UOjHZDai
/S3VjnNWmvkyuMS0F3D6OCsh4ZLAXywEtNMENJ+LjRCU8HX/jtCIaBrUKeCxZQue
Wht7SepWtYPga3OdSN2PkeWuQa7AYAaeRFBqzQePfRhsbZzu2Ll65ExhRvEMhgaH
CTBbF2Ymlv2NdeK0Nofqg0VT8zDKdj9NbcVe5ZypWDhGkdO7YuqEw3A2ShJ7SaFq
MjF36c36zmr5l5E3uHz4+IyhagaXcb82qNR5GMpGM4XVxx99uBz0NA5WWXUrvm1w
5+Rh/KOmoFxwe/pyPu7ntBL7tcYZSRdrOZWZQSdbmWh3yzjRnmorJFhenctIPMeH
OzHr0MjMg9//QsNSaoO7fU2vJ3Mhr9bfCGj2WhFOq67vQKBHUnoAzwgi6dUhYeWJ
2T2UcymDONfzAYBKPYzfoXMC+f9qiQVtXmDkNXLkorlfVZsHH0NkyfMjk1+ZymPA
66cx6ZR/27yWMVvg48IpjNYbvswQ021pyO+ByD0n/VvYInnnNtKgTdJPpvJrMUXB
kt4Ps6/P6DcfIPTrcerTURK8JrwxNUsaPUvw1mxlNtZnQ2D7EoOwyyYitjXzyMkz
7iqvqd+H81ivTzRVGb5LsSyCZ3WyOxV0orJO3+qkHv8WzDY5GLxyzxoBP6Aef7aL
BFzjCsChEJ/fy3uOcT6OmJcRMIvKN9NOoGoT6lrknVHPb87bO1/J6UGdYh3yA6iU
4g7ReUxZ9DdDqlfSLQDxsiPs/vLuF4vZQtnyYnb2Msegtp/uvc2u2KtFG8Vt2v5X
01UQx65GEVV0K0111QmuGjEoUQRf+dHJE9d7kKC9blQ5qR+z9TWRrBluusAIoW3m
joO8YmoGbqDvLHbGGM3WgHKmT7kpDKfhk6XnK8y4+gXyEPxfeGswgI214Ht4wsZw
C5rUHdvN51oKwj9e+Wn9JlCD+bavNmWX61hR1+S4YU5xP3QRkGpac8KWioXln9fu
sRnslKpcHmG0aio9YgMHc5O1Amp7YAORbrhlLQmZioYTAnN/fztvGnJbnUz4CUSr
v+fJ6znbDyuE+B9YXIPckghlQnyjDASjG1epbr/I+N49gUs6fn1QrgyAcHFd3bmj
RdTVijv36+1bDo2tET26uNqGjwjew0xS/hyjPV8mPo92ms+xsD6BXrNBr9crRMo6
AWtVKsKAEfzDSi8kUvksn0YXxYe8P6iYcTEseTZUp8N+IBsZsMjaUseqgA70fF/A
8R27WB3tlK5GSrnG8+cKDzjgaLUGYw16RraGyOdzomOm2zCMPpTSEKNt0HgQRAGu
sAC+dDNID0DRP4ET1yaW7YjaXe2ingMs4tsUE8uiYkCq20jJaVS64I9U/DRDhga2
l/heq7HMUTNjqvN3olkyvMSBp/voB8NyBzFLsdjzViU8ZxwoTQkAsyFa1PNabolz
wIykDSOILk7UFq8DocT+Kg+43uLtLQKRh90tq4rWvCjWSBWfN1sf2R2+IyYQJ1UW
0ocPZrH6PVcpzPk0md5OmAdj+IkAM1t2ju2zcQt+GiR07RHRCsy1QGYUoiGI4hzB
qgZ1X/1G0KpjV9EI9WoM20O05T8etBVfGRuSkSC3ZW0Vhg6Cp00DSBgYrwBuSlI/
yDHbDx4geJMSVz5Ep0Alga+yec9xfVAWPq6C5nKjq+NTnjwFpABj6LR7rz4wZcAP
CkX6DYvy6BcYK0a4/AgUwyp3soImNDNnpwQgIx7JJGVkf+ORD//PrQux5QV3tbD7
F4hezR6hTJ+61wCmJogUs0IdCtfqsbgTNjmorgNMZBEjOqELB9wNIDP2reHP8Wua
ix/YabGur1zzPeLeLKanRvysZNKVzTLEOeqplIIQQ3UMgw0Jb42mv91T0VevJDBY
En4yo7LiQFsmtrANrjMke5KLouSlCu8wHehy84ePzHz9r3z8wcQ7ZCruJkWhN6Sz
fZfXtzSFc7hpemgXJgNT7ZVcEhmgFv7eRB5K5ZVMQHfqca+SbdKQTpbfPST9h6Ed
FKnx/Mr4nkaC6DBl32uk4ATMEW5dMIufTTohx7a8hjuyJ3zFbBdHwHjf2KmNTEs2
meYqdPM2fzC9gpw9YEGPAtXqy80pMHPNHgdpxANjO31E6NwJJuQd2XSJpFX3Qyhz
7otc3nALas6Ew+bhvrzdd+uFxRFLn102rr7h6SDvcbQeV8owFvji/jzfO/z7+9Q6
N9spzB1Jf1FqvV0Z/T749UIB3arjd3HN+WZHg2Ag0WO9Ora9m7d2TFDnG0ybgsfL
MUNp6kxWAbuUycAjurbIyZephz/VWnoHouDyFvjvzWKjF2guZS/5SgbPH5MbjX3M
iY8lHHMNHdjKgAfXJmMPmAXhSuO5JnzDSgUtP3dlGj8wvFtlT6mEPgdKiDsEo2Ww
PrlOhBMytA0X/ZV/s9SZ3Iu8vw4P0oX4aRHPl1ww9oHz8OJSnkB1OqJ0Au7tGvGB
Z+E5MNkNASTDGk9hRd5U5MtXOu/mgYnZ1f0qsV+/xgU4gcRrsNPVuetcPNg9Jmqe
5gLwsIKwrt57tM5OPXTbR23ciVcFq19IkVAcYhRfUCdM9mZWTEqDYJfHiFtU2I+5
Xzgacf/MGVFu966PaRU6MzgI5UCKoJOt4omQwZsRUWh1KyY5kOoy7QOFvSLtt4kY
QhmO/ib6Zo2qBf9PyRM6IrS+UABpPcMpEyDpQutFcJcVxuEPUEzW/rAMTlOqXPZO
YajR04dZQ68Y0Ny/sPjZ+PcJYcMssvqFk2d0DsnC6Eo3S+H9uUNEm7F6J6NwIvKy
RPqJpHxBUTd52+jk7wLLd/BIKxZUasM3qi6T1u5oqVK2fb8kVbNOs2uDmOhdQweQ
ZKAUkAcnxpKYSfBaZ7eCA4rEzrTjOknU2DIUD1z6FPVHZSU8XZkWFUuxkDDhc3mf
FKJ4M8GCzTlfhUMm9hjlvcrGs6wrOTJg557PsZqOnXwKOEF3MYwfSnJo6vqkAo68
HUU9hPXjaOZuARhayaYp/uAIso3zMo4nWzdL/ubh4RUzE8cYTrsqBq331ycb9lFq
Y1BdNKLjmE02HWn3sxhyTzQYJ0Qic4uol2CiuObC/IcZUVrGeZ77Gqn2WcjnBjjQ
W84FjD1CTk/NXIzeoScKCo7/cZrNzqxCtJoS8GTmTCK4eKcuCXc5LnoIndcyMptx
WsjhN6eBUTN4gHzMw99AaWkt5OUGp3VknaH50JTrqAM63z3mIb7Fe8YysyzHeaXW
2K1OlRp1BKbQqbTBDQyotee6yVrNx0hTFUXq8TktjeE/kbKGInSjHF0Li8t8ZdRv
cp5doMgqCktZoEBkbu0uWaIaXbSA25AG84+9i9SAK4QB8SntQpgiiRFAKHi++kd+
7yYc9CiSHZfiI9QiRPQxy2kXzrzsfcxjfSbcQhoJnLcZ8IeDwmSLMiipmYXasGBR
yB/yYP1QDPFP6m9CDcwef7uHy+q3OT8T6q1+HDpYXs8Y7EpIeYe0Pj2eTHsYRCBJ
x3k0i4aWxFbnVHnAkamtc3ouw7hR3r1a2GBBsSmob2MrljuwroDpmj8w9qZ9/Ypo
cVvrc6ALM9mVOKgGmP78c6VtJGQi4zD0evT7R2SkDk+XtbuJ6arAaab+mGziLgVx
lRmFdJSb1+9+nF2YJ/R7XVTsVw+zLClXFzpUFmzUkhY2BFe289t1Q5FHYfx25dWL
ZwZrN+IfeMonEpO7ha3MrfscWaJAAJvsFpnhvTT4i1TVxnSXtlhze7eImeMHXnSo
p9VRu6ZnGi8gA7nxduVUIh2hGeHNT5J5E7EOC+Q++YYAbqWVsop5B8mHPFcwEWhv
b9ec1hDxhyUF5nXVAXtWJa09XxJR73bMiuKU0TiF3ac06QrRlNSqEDlyZwNGQoj7
R3Krw6fCg1uoaQi7ufTfQ1IEV7BeVrXHtBb4lOABzI6//QOmKpnvTjhOXx+l4/IH
P5tYibRGEaPQIdso9eLMJEldRtuimEO+N5LoSD5en2lSYuYXqYMyUAZy/qDK+CME
FinYkfEp0zWopG9mK/EWkKqBujHH4lWXi4FIM3A7J+ox3WgZFwaSmpd7I/N1ru6j
97iwhFuInufzgaaWg4COUjsJ3Kp0YFalCz541VUnqyDAtqJDrFAvx/XfWy0ine5F
GClCD3mZxDD2W9qh4sIJHnN+XR3im37IMhTADCLhraSnN28Xg0j8wH9M1suW0LXW
p12jwMzL9FKSazNDh1FLyfmky1CaIq3UfMqtJXdyHNDZMyust1aSwV8wmupO+ajw
V5dDHIRqrbXNVNhhbYyHp5C4KnOFk7s4J1sMoBllXvnLQzI54wdwRnDmdGlt9LO2
wLCM1bghd/3NbodprqD6E0YhIVh7cODIaF6QRSI8rlIe4SG1A9bdeM2yh/OZYk+N
NoHjZbd2xc0c9uSAygs1akQEcwP42bDXjR2hduFvzIxzXLVfIzdjyrAPq05wbtbA
EqTuLjS/jb6O3ghU86ifShG0HPWHw8WPLENlT/Lf1mI8R/bVEYGiGo18br5wTgEl
a83kK3GaTA3erKTRjZadQtPh6/U88sS2h98fgf/ZC3pOm9HdyFkumitqGsHaltRc
kwYjLLmhugv8kMpf7N3lbhfDYmQzjpd9ToNwHRlqIRpa5R5Qu9cOzC7JhOFb4LrD
GZ8qbh8YonY1Yf4khpoqMa6umOHeE7ScuvC9Iu2RmnGrYPdbgcB2uGyU/ya6bEpY
sogBP5CwfLw0hkObSWhT2hOMBWPTyteeH1llZqWZK8fK7eXWvHUl/g0Jk7JR43K0
CUPHiug4AD6fpyqS/6Qgrg4W3Ia05Em3hlAeLFceU5ut2WDeOPGvmiTo7t8Y9zl+
YwTYmLzMhbXtNrskmVpVZipewz4p9h6EW4qQGV9JKp36u+V0QSsQfYEnn/XsXHba
1a5ede78xIctcZeA+xu1IWwlaj/3rjBEUibrcxrZJOFLoTziS65rOJ394oz85Q4u
lU0AA4q76c6h16fFFln38pU1rX0PURcoiHGF4+PohrOCyExHsEsLtBssv/kfgQzn
45tDLmLuRuuJylpqhY5rID/oHShGpIpNbW1qFibQBvjsfNBs7M/PYjUN12+JPoJP
C2i54X0+JaZr/HFhpCWk04EaIb4E1F0TLdq/O2XQIzYuv7MoM3HCyUPcSottMR5d
2RYG5YCXlYeTt9kG139ocpadAv/KZrJXLIqYs/b/jOdJobau63X9ndGqaMC07UN/
N8uXnnWpK1+jXxcB1+k7KnRKkFQwm+9Yn3NbB9D9JvquLas+oNyo1cIycFD0m3QX
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:34 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Duyo8tbgPjzYo1wuK580AqgdIsMEW7AvBWgy7xYIPKnrL7WCFbvCmY8iqazqhzFr
9iA+kuYLxF1f1JJItcI8EIz2Rzm0fCEqm3tTT5krRDcpzN3J8mdsbggtF873INUd
vwsWorq74jNb4JXuOmKguAAWkvishJGjzyni+QgcymI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1888)
jHSck3q+177Z4S6jLH7Gnub9RIQLRT/8ulzmvs0+BKClWgwcLRyau/JmItVI/wVO
gkht5K2aazxMlcm+1rPhYfmDfqGbRNjImx3xPuf2mfnG/1Oql87iFIcwckeh0e53
PtwDp8/MfjutpN9pXFB7+arTo8FQlMUctuobuIcX5W6/2kX+r2ntlApd6dRqi7Mc
+rC2F9zLz/B7mtifFlWGrvVQku4RjNL1kqsnVXIKVNaEPaFIfsFtOsxkh2nCvbK0
0ffNDbZxxWQjXyW8WyoD2y20BOBtnyeUkguyPXH3vHdhPSC9Ean7Z1dJ3pXPMbdn
k+29tEYmdQZD2x8zcJpqmC9L5vHYgTvlWdyc8VjXQjQ5a1ERQE3QSLpSN76PZhw/
jwhWw1nSMdEjQxwcocF9LvUAdvom5OgZ9L6P9PINLJk3sfZQHykh9fzTt312Zy6N
nCw/z/VP/AHesfiqxsbUYBYxFMpDzep9+PGuZoSSOv4jdgHCmIhOXdqCHUFsOCPu
6PpMnsDcKrtLJ2v32BYioiPoZSAH+UkD9ltt1aY0TErF676yPo8zrBBQ7BfiJ4IP
uEowOJlLbjmsdX1H2pFWBv64Bm5y5iLAH+tlKK+yky+pDm+CRlnDlNBpMxpTNqdT
nKhl6TX4E7VY/NpxKYl+wZheRTvRKs4D0K9dt99f16JpAHyIF1KeAhXgG+8A1kvI
Oe6X2XPn4ls1oMJqFVB7AhQhmfGiWfeWSCQhMsKmrTWv2uzcvwVn0Tf5e4cnFUYw
Fl5nHMJ415K4nlU2ivvb0vKrnteRG/b+hNhnKhJC20nxAhhLVmgvK2GHkv8u8R/m
2sIIXkTcAuFqPAyBC/iv5ofMBT+rHtJzB907L36zyd1bM+mtR0eDXxcl3+37si3v
flLnOyqYCWapFMaJV2tLv750RCIALF6G1duk4ATqDUbFJe+BwQsmv/PWvZOvwCdR
9Uh0fa4XvXtyxzU+1lfaCepPSBzREHg2c4/se03lVYLRzvWPl5w2WbiPTYVAqmoj
o+hB52a1DMA+94Sw44ffP6vMAUgVm1Vux8nB8ki4hgZh73af5W217ywD9woB3oEi
d+K4R4h5hpwghMYAw16eaj5z2vwRrs8pz6qJtvV1UenALsica5KkruYOGoXhG0+L
JCabyBus+uAquggcoUrh/NjQ//34UWpT2op3WhSdmChawrZDDzhfZsPp8YPIadwq
IV0DK3JKxw6VmqTY4AGroPRSGyO8a+FyW2UpYOwVZ3ktAOIhzWOODK/1svfyoNjN
iNU4xGIqc7gMG8AduaILy8dVD0NPSO2y/fWu8GPsHNBXCS5K8ubKvWR+YBtHJttq
g5q5m4dDa/m4+VeLHVKwbA6wZPlZSgg0z6SvZd95jKGI4SUcDoDjRiwrkcX27f4y
RwdVTG9wcADqfsaeDNFlp0ZyyU9RUF7SWzp8zOshklWKerEcrrLLVbZ4uzlA7y7v
ChaW3R+nAsxA4B26aE+EbB3TYIwWKWC3gzDufbyfeFrekSWtvjoXb4dPwJcMDLif
+IQH6dPtc/8HHbR/6rAHNncTSIjt8dcWbgCPeeXSeDIIhPhGfw0WPnaO+Ba0OruH
gqfYZdgVqMXxqC8A+/zvPKKcN7dPL1yYCOXIPTwHBASGiFvglwBr9h28/ijO5koo
7XeUqZFRFtgyX8g1GAgA+oWk4ztYL2pXmeTAEXyWozvlvU1D0BXDLran4N0MKrZ3
H+bnoY4mHszUvQOWYxafBU7hShO8HUqauk/FD4Q9X8GyLqSY8yeMJkdxRMyNP2A0
5ca9WqpNgq8I/jW/xuNPVdQdwis97xZsZglPZIHoulnDNi5q/SQycISHDd95UfGg
dfceIalSsEz2xurZshXgZdefyIkppEpKV4DH2ERBYSI3uz4gEO8ASZUZ3g3Pz3pv
fgnmz62+5j1VYrVyFja1tOaYpilMM4NNPJzGqXiJyNZsucbI/3OKlmkcRds96jso
1juM7BcQauyS8BGhSDM45PoHJjy81rk4k2YObU6fsuzqon8NlwcphPaDtOnEGsDk
yzyRhdSXCCcBWV5frL/n3obUGtWH9hnEfDF1jVqbX1OEOTLDLBPw0X0Cmm12vqo+
6UJz8r+2Eo0P36qVsiSxfGRfVoasQne+38mbhYwfpYFVHkiTYJ7pKy8tbNlsMM3u
HA+c3SA0XGqKqOhelcZzxZAazF97/rhgNn3yN+A4qRdIO/d6TgWw8/SFsG2c3JAK
M3bj3og2KV2EmfDcGFScNAFP7awEb7nIILp+aXxXtndz8PE8sEu06R72R82J9eAt
BPkdAGDdK79p3F98fprNic018NuIdixy5inQWUnJ33uTkPVfJJKWJxmvD2zwKoDu
3R+MvJ1v3nPoVoJGITZ+FMhRqspLj+6EnqPKk64ajxu3UA6sR4Lc7Ky5mEgecxeX
VUgIZOAn2P1VxqF9iymSMiqTy0RJGKCWjB5AUvxEUMyyPLfwP9w7zwEtuwvezEkB
VUreLjxsr2zNIomJRnEUSw==
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:22:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LsEBB1H2LTpHd/7lrs66Gr0t4fDV7G20FLonNLGNo0U5aZIm3u2hKN87d+W/gdyj
TQZsKcm5rviy5M3lqI8wYMgWV46DV9i5an1ZOhDv5JzLCYJfLLVPp7pD09ife0vp
6Mdni3gn1qzu4PTBZwJYP8qsIJbRMl18GxcDitw7gBo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 49456)
2bwVQa3jmvlO/aYyGoy83OlEb4EIRW8p9Rogv5PXgvKvYov2WpY+kKtgIhUybpE+
Y5Jycy4XT55Duo5QD4pxrgoZo3xSJILATyiExsLOGgIl6GWokdOm5SgjaWB+iF2Q
WbRFlqqOvPDtxRMi5G7bTg5gd2c/0efqD/cMoA/jZbjVK+iZe5Bmwd5C4XyDfm5L
QOuVjedP0RK4xWU5xsggx2aVbDerfAaKxHg4qMC0hr6qb7csCGlokQlGzLCiCaIw
NoRor0BURE62e63/kDwsn4OKkTbxQ5Lznv8G9ASmkjYvPnwpRD+ChdLRU7kwmjyr
ChdAcKDnJKhvpKoXVQN5eSsVE2BREgrIILoD/okzoQa5vhw3P85zQWsdxUamCt4I
CGvDw1/p0FF1wgh5n9AFHdY8G8yy7H6Cr+vhK/xg4b0EHySqD20CEThpNn6lfnP3
RWMv2a1yQvk6PY3xl8BNK2Izf9wiHO52q8VLRwEb4ivFoUDwRrkFkt7T4g28ys1/
5LX8pPsbDbzcXaqh3JAoIC3m0IDN8xD5TO8eL9iU2SmIReqjMboAeo4i5YfiZrdF
4Jae7R/W9vf237ldGobm7ZFPuw6U1T1IVdAq6IrHX8/3jCvD0UUZVeFhU6/zVBrl
uiZ5jjsrNDUpgB5YH6blPTB94cuBIzUeHRrSOzQAeMpzNXEAJNl+CH6YKsHnky6L
+B3c7ETwGywvwY++OZGf1iTR95FS7aSvl4sJErlK86UQ+hIPKMZg4MllhkT8XOJ7
9bRIeFz2LiuN8X++cfzIY/WZ8G85XwRW8pHhweuKgN8zYACJITpI8xg6Z1LAS/ay
vUItXLn/+W/+IMDhRLKBMTQyWYDKzDnVUywsSq1C259ZDAk5f+H5VZX/IJDVOLZQ
xomXBNtYEdga6kkY9qnvTP7707ww0yIOgvgSLoiHPo4DrqldsGIEOyPqLuS77XWE
I9TKrqhq2IOo/BYcTItjEqzSoqiyiex1/h0bdoTfyDqiD3ppHG91PJAq92+osYUK
O3+mWSUxoYgwfrKp+j9M58ivG2busc2lr1Nz/N5rDxOBef4tl3p063l42Td9ee3H
GX9LoPV1heRg1sWsSFgEunFYRFPfhpMlNOhgfUhcj+jtJ2eZwu7QOHzR9ovr9pM/
ENzMHX6+nMmSoCsCbQMgDVgdsTfNvSsaG59z9sW/07JyNyJBW+V7pQ7fpzmd4EaW
5Lwx4o6B7kfZwcnAcFys5JC5xpzegM5LRJlYV6Hub1UVNo2C/qXUeKTddysj5nGE
4I4EuvbbDPB6iVkpgEA27T+s+Gb+o2QN5K21ftq7o9hkJ1x65E52Fi2LLtO7L5Rf
LnGcGkp6+f376EExipi3huTnL8bLOmcss79uLoqZyM9uIXXWR8AtUtMROXrZi/UA
z9TRa72kGxiYj16IKigqiurvg3yBIMEI4Uixz9XNruSba1VEozHApgsC86jEaUfF
fQ4gH4Nu4OA2Zm4vaWeR/vSLa+nl0LnSsLRU8l1OLj5CXka0sanQGAhaNXtNworv
AZYENNCpebrXGeibcPt7FI93DqBULkGap21h9vddLYFY687U65kbmOz/XOqvZT0E
/LKbzssAd6W31MPfF5MCaoh/vLkBqMaSuyIUvgxD2+sEIAM+AQKMJCuqjVnA+Mtc
jiXfEJclBRO21uI57LDSv+2CAwNuJQFqIFdpjdRdMgryF9TTt4FheEBRn7YuQjPL
C0SOG0VePgKWfN/m/gVwHqQHKVB5CEh81utLAyuqHkqywMuVEhOzLcdFV3nKcE8R
rzwnqQSMHDWQAYAYh6XOXL5hFb98r76bZAfyQ3ctaLUBmHkXdS6y/7hX52YnnYGq
TG0huh87Q7863BsNCfX9qAFkc6vTsyGwvqEGULTLJ/7exTH0+hKr5anHnetkuRxe
fWwTVRjRaIcgQAdtAghXJD7A+wrFep8qiQr2sV/TtvxOTvdOuIejjrIQnRcPBv2/
YhjvIiSOPxWEffYlY+I2GDWIAfZmeg05WFvyh6oKHgT9DbjT0zF+PjorwL7L84FN
2hjMzOs80VtIB8YfzY8PjmUCd/X68rKL3AbKtrUk9h2NR9G3hct5jzX+kQETajpc
CovyhuCT+A3OxXzYVjnC77DQHA52d+8SWBRjRA8GRDKnD0jNkLZSONWQ9RE8UhRQ
ZMah3uDtxRHqleAfPXaTMZ0VIq7lDmsUuow2jY9XZ92V6PjdlkY5g/s5LA4lKgLV
WbVeZi9e+i9RNMpOfRow+P1dTKo1K2ZhVguu2Gfo+tE1kTsWtmflNqZ64ixNg+cT
f48bfGXKZ/v9t4tk23ASWpEfhRKOuRo1wRtEcFqZweWRe7M4x+U3lcMYH/ocMtOg
hs3ULptuKC9HL7Mpa/BQpeK5snlF3Bi5oZOvV10br1VoIIAHVuRy2I2LNS3YCt6U
Pi0A8uO75G+29qOT+E0Hwm26Lu/DDs7LGqBCwA8eESP94V9BXgakKWl5q7OStsEy
OmIbq12l6Uu/M1fq1nLobr9S1IXF1sogTV3jK6mgxey3xRB2zGf/RWVf3WeV0dJd
vTMH6u3PWJw/4LsCMywpAAoy5gIncvr+5FWGVJoOBN7GfLo6Fbtj8lCCKQSVHwjZ
/CqezuNrEoIO970/kNDOgCFvLTXJaXc7ihqLYtaS8Wfr5wwZr6qNbbBCM/VXvxbu
jgzxbHw8jUbOou8CPqWsvQqsdoARc98D/XOJSsrktWTnCktvduySZA7BuPhSgWE4
5DKniVYXjIYY4CC8z0phu5cX9BeDdeqVcDD3Wfy1eihNK0Iy9Gut+i9pomEU0022
1nwTaL+m7TsTGeneWST78S3fYmX50RsbJcVAKjYYys2Qq/0ynm3z517BKHHMp+sf
UP6Bka6DRkzm6pZ52hV3B8vkQ3DFR2wxyPxkhn+SaMtzjRC5eKW5JSdFZYW2uOAp
PkuPjf/q0Vpr8pCncBcMk+V494yQaAEO08ByDY8LednHU8lg0idiTNC4M5ydG1x0
zyRx3tRODIfsN/6hci2dZmhMOrsP0ds4/01azGPF9K7ZDsiv7y+5QTfB1bkiGvBU
xPopEzGQ5CiRpRQe3tQ+Hmho54F5P40l4jbo8LvCH8UM3gXuZlGEdvO2mf1WQ69i
oissXZNockdpRMeFUSSBgz6LlUaPrmyrQbVHN+3293X/SzRUnAgKaeJ/QxPMU0dR
+BpEZXV9D0XabYUgxPiazsIhjhAMovOHRAiadDQCiNkk3Zz+wWQ6piGmWkgQdV/a
VxBU8Ok356qfsCrvn6oRCIAOlI9IrkmL4AP7jJlQK8Tz3j9WxXknURjAnL8tG6Lc
w5COq6aM6s/jMVTRovQABGEWNKob53isG9hRS/gG+++kMJ0Ygz1YH0pAyeFO+z9e
vDLANKR877eqyFBRLEOxvoGLcdtgATOrLfbChvy1JTW6ci4XI61q6B14Gy//rlRW
8y4Rb5PyCZ+fzN9burYn0ARdO6B6DMBhG0xRunySbbga23r0w4guxrBpwk2RRBK8
9m72nApeppeYB16isZpgHuFvTTMcly3GlgXzlYI+OAET1e+n/CjmpkNXVchs4U0M
byzMaT0YOt2YOao1023RoUhgwL/PnrWTti1TRGETLL0a4A0iu06Tof4MuoLTGoOm
uBtLK+VPHQuz302c5r9mN7vc9tpzHzK4Y9SM0LAIqa9rClUYpfBsU2hhUMogdLiA
LuE28WlKfK29r65D4pujjy8vNtwUUUlU5ibsaSLE/bfJ849saDgCtMzV+8CXLIz5
OVKbiPTywYR9nHu+j+lHPC6XzehT0tvSS66ghQ0ApVEvvCfNWqf3fzKnI1fvZPBk
atFHlE/PU+/pJm0ZCXw7zbX+X1PhqG9nzotRMMUVWD84Wbx5nNCzm3gv/Jxe4Rod
mcdI8qH2zUm7hm1qKtVXjB1UeedlxMAhCBAW9fpJ69XjA1YxI1jjEEmqJqd4LlQr
i23K4r82g2xjulQhpAy+usXPkwwnwdGoa9THja5aSOI5JKEGzNoKSxJZUTk4B9eG
GdNxqSgN/tWERk21Fg9ER6ad4GG0+pDx5mo0s9P+BrXFpbIpZI96oro+u1NdCHa1
zYMPayX+Eu7F8W2QJ4oOGyKJZHisPQFauTvytEWPyjQuil9f2s2YgKjqW7qsiSq3
xUxUHlQbD8YTUFSVdpXGt1SfD+xDp/aytdxr/6m6u6FyhoskcrqKuqrKncLf2Mb7
aPvwq09ibEPqezarI0Lp9LWrBZ2e/CwkDujkxGzq4glFwqqWVKfS5uRrwRgbaWTo
SYB9YxU9k41iAnWgcM+yEomlFI3Q6r9sGfVHfSjt/EDO7fTir9HIh/91n8pjp0ju
+ia56Hvcd51pjV/UyvSHsYHanc2SPMK0H2UOoJ/YuNjKes2DZOnbYFRnr19QJglv
wdE5s/BDYW4iwSCmkf64fMLSb2LTjBGxoCZpUXVVRYb9SEIZi/5/Eub1ZJyzA58a
uhdx9GbOoNwUHu9PF3oIOmSvFp+bo+zyu5e6q4PDHlChHIsFggqrPrFcKx92Oydv
ri3k40G5RpxVyuMNifbY7YEUCSVGUMsK0mQNG27SZAsf+CUN2Y4HPrPd0Y4WhO2F
rfbg8IIfEb5b6VTdnyH32dIzXh4w1ch8WST5u3RaAUDw8tutB6rTwt5QSvA5+o7a
MkR5aZgMbpqNVLvUPB4e/AVTohzo02C2pXQqyvSPND4Qm4S4uRe5EOI0BT/9nMPM
G2HRoOZTBXi/eMI+7yUcj5FXsLoatfTYwzBQbzNh5G9C1fXz7d+yY7h3PeacXrA+
G4aJlP0eWweohqTYgGiL+YLC+VEqVkQkyERTDIKrMcq5jKuaKVARLWhach3bi1Fk
Sabo4cC0aysVcPONq00STqkA46sUnFmmxb9R9UsAvkGp8Cj48BheU5Oembc0RMjU
uWz4SrxzoZItEmcwCHNQsxXHDdJkAZp0us8XoxnPXDI+bUI9NrGa1cnihZaJe1RL
8opQUMCBEVbw84mDnfLzM/8zspugHbb69U14H8v8C+MRx5hxVQkv/Imv8U11pK8H
4upd+CmNvd/1MhDDqFhj9gQ4emu3hjikmQLgcqY0BZC15maHFvSNhDBkGJsfr371
x6RrjYXqe8sGZ2V2HROa/6SliXDeQoIFmXBihFRQJLO3qcNVt+innuPHxAxYgUmm
eUt+0U070fGZV4PAc4GDctF5oAFGHS0Q6K8k7suqQDSK54EZ6scssK+cdd0c58OP
ep/6MP5i8d+ozN9vXV4xbgZOhdShSuKH9OcmKpgNfTLLS7SVjRbBNFApahN2z9Hj
/fCv6ccZZg0uvhsrFAWVf3Hks89VcSFdsekBA4v4/AHS8KhH+NUHvKNW1olMOqJe
XOFqTb/lxnHR8WbljWvhCaAQxGB5rLrEH6u15l8tsS09pO+fFyV5Nhd4LUWwY4v+
qDSXmYaRy8TNyyms+jXZFHUkTvG/TPSMjQx3uR/BLT8h27bLnZOGzkh5bOd/xr6w
4z0f/JK4j5000iKzXhlyJcIIpqSvS7oLHj/wBQPgTKz7Kv39RTTYnsvngMORtdOp
dR6DgCPqkDNxczBLmKMObTjGvpp+6mYyHcETze8jnMXPcJp4W98xtzmqk+fKKFWx
cURdH1XCzzx/mPmhthwMbRkb2WRzx10yBl94ET4CgoADxY0AfwdNzNMGmNX9wdgG
X6RuA4e/X7hJZA6hGpLNArjdyBiTbOBSfSxoU8qZAW6KOsdGyz4pJIHoPrE8cz1u
ueE+24pn+8TZONLMk0Qrk2CvX0bvL3JVrlTYx/aZighmUziCWqvztvZuJNNE7C+l
VrHVDruIOEDdQRkntdwhjOX3BPxLsRZIh34EinwBQ5CeQa/cIJYKqCGWUmz/UtWA
GjG2Q7Jg7t/dISp8f3H9D1juWksvY1Wfdyqg4ErvJINa3X3TV0My00DKiSBe9z/h
Kf8wTkjjrVawAoH578OvPGVnOXXpzcdIAdzK9NMQ7ZvkmY5/mqxqEZwlBzLN695G
t+ALpxWnSIPKlkpnafW1GfPcxgzdNp8WL4qJmFHD6V2oVcop28aHZ03MOoRsPI+X
UHkaMwZObUeaUeUYevhe6hGUjnl4DhC2PTwQtG2PjMfcr6JxY9tT8WfCb/4C0uLT
DuKKNuMcu3bdEKsmyGPUjVdVHp2slnxq5Qksp1hEs+IUgVFE6LZ4npE+xcSe3lbi
tLLOd2ixS/lv5Fio9c+rmLPVgYOVTmSylzH8nv2+gl9nS+s48iXC0sSBRTSk+cQf
lD+ltDFtdSk0gNCnJqOgoM5Zyo5yKFNN0aCqAX9L9CoSPyCxcH5r9nVkZ+afIsg7
LCr7Q9nrExOhsYq560VPrZ/fOEavF/okkdU7NuYsMidv1tBlqe/nHGUosAfwFb/8
jaaLkqIPRKO7OzXxb0MIUsMXhHYD9mQ03Y4jevD+oaHuyy6AJmUHGv3++fCapjSh
gkuI4u/66yM7Zi6LEC1NPBmuL8b4n8GIpHdoLspheYMPuWXe28/Ynu+eiuQbmue+
JqAs0cfMTwbCSU65cd17orxGYM9OEBPrePdjsZoIHxF8QlEsxgH9a98qk2ZLITRS
9Cre2RURRMExwdUF0yOPMYYq038XMnOxLWcoyinnN9Eb+ftjnOG9LtnRqrHe25FE
wq9rDhysnQhraGmQKF1v3FRXvtVPKwRiNN8wKwibCIzB5U8YeowrzksqsEtO5m7F
DUuGgW7egE5a5e3JrvTfRFT0FL7hzVODw/LLBvnbwULpmI9ibMULKmEIgKoVU62Z
/mFO8uRb5JSzU+AUqKk3cMU8sKdVNBCFTAC7KwjyH4YLp2dmHKNIPCwVBfeNgDkl
TOd5+r6YV7e+gHkCGsB4iO/5+wEqGU1h5JbKb+DbL0iwC75FMO791CLPvtRicOfB
XfTpQ+lvt7jaNoOoV0WzIGpp76JVoUvicBI13aZw6Lvk+xADXk70cEXjOTOEFo0z
c+y+mHdUY9zjgZspDKu60jXKuN8nI3HHropiDr3BJuOJxoViQM7MBk7VhUfAlXhW
ov0QEzHAr5cyi20L92ev3wkhRWL3RdN3eTVmD5L0WKB0geik8VrAfkqt/QokCzHF
CFgT7sgc0ykBvnQtHSjKKxSYF91mxI7FzEs59Aah2MJUgSaAgzWJZlMQpAKNbRvc
GFXdiPokq/E6KDksqZHQ3Rlr0T9/428FdgDU8RIv3HoW0x2UEhXKEdaIVfhIKmqB
6ppc07gDJjOfXAQBIFdW4Xmd69kAztPLDVY+Vn6gTY+Es7eTg+4O7+2KN1ggWw35
u6179uPv9vOSyflhIotTWBwxlkxGTVAcYAMTM1gGr8uF9nHnMWB2iq68+NmuiXAS
+lvnmD83WTSSo1bX3capVZYzBh6c7wc3H39fMPNr1jxqdtrLVqmHmP8b93ccPeSt
ilzspZJ/jT40nVqVo+3N9xDKs1LK+0irKJWdr/5pz+qd4g1486GsAy1dnuQKJe/I
lK7jXnDV5bIk9kkaYQwX43/JJL427xVazfpkTmoibilT9tMbczMNvMAwk8kkeEEq
HDQBeqFy8cvWxZdTan9prbeRxTBvhL4Ol38pL9tvqKYPl0h0PB5L7albu08kBVT8
DbKagbVuTXEaDmYlsj/YZRNYc1RDKuv7dw4m3WAgFrSkRdVUc7FN8/LezzqxaK/s
yfu6MUB6UMNrUSoNdtlZktqdr8R5AuaOsg/EIDneRpDWituLgM2MXlT9UDr1HyDP
MJayNExmJ+3nL9hLMD+foLAreP/+cCfwPFe7hDjv5Cu+Tk3pyufc/P+/sfQYpz/g
93JAaMjpxgkVnrIFydxFYHiSddryEW70ETNNu6wbmkImj9DraFet2FpCmlfBQkdL
8pxJrQ+H21U6JPkMaTPzyO29XAk5RGKVXQJLklJXPPjJLjFGoewh5N1j7a71eT56
x322zJkuZwq39FPd7MCNNV3O0o+WqpYVOa+pJfW3TW4T4as9X4ldQ9nEL8AlxAdO
Bk5fejj3lT90UBzBLPFQItvB43LmU+8vQYyv70MNDxRW+g0Y4ctz9hH2w0qv/6VA
Dbg8Se5qDPhxxOkQrB+X5DlLRtHT+Z/MEdnfMSDIReQcUrwDrIwh33p4IZ5WMptv
XOru+gQoTbDPZxUZtCnCYLwFLTQByiwDEyYSeXsfYXi1Vb0mq2iNS1mfPGzWPvDT
bRZv9fZ/hp6j6EHPDwqkLZeTvzRIHiQT3zx6keF0kBbSE83lKIksv+1A7LnzHqYC
DGQxf/iSX7SyWAmf0ur62R23ufs1/GQthTf2CHNwQosqZQdj1cViRwDgMLVCv2+5
1XHlHXqdVbKJtfkvk48JCF/ootnKfm2LIPseMI8x/6kFKpYaZdb51ypoVTEN4emh
SisslzzjCoRk9LIQh/EwShjAy5hBIQDsyxs6foLBifvELfgYTa3DfPcHk6WWPR6d
ik6owP1klD5/K8ut+Xh2HvuGxOD7PUqmAN6R91Vm5SaNCP9TttujymBFfnaIuowj
d992GCc50O1GRofzKBf6i76Mlpx++hnub3Hgsu+HS8KiGJG4OVAioahrXwIJ6BYO
q+79lsDsPOk50viC4JacfOTkqCfcKZ95obt34lq+lVjAis7NTFGrkciX5LoSvitR
j7K7Nl6RYW4LRdM3W2RWwe36dC0WJlDlecgW3sTpcVVLwG+oxQlgFQZNAVMOGUqt
gmzIebMN7U0qXatsulW5kKjMG+4N4zEnVzyGWWrb77IyxQYa00MZWadQ3R52JT3n
vhxGiyG0+AnAmkw5A40QtN3zsad3AgTkwJTjL4EmF+7LDaXJmlump3EsHKS8PA70
BdIMiYzqEPe+75zciznHcJ/L76cYeoWkkJZiXodCrdCNhAGavPZ1SaVpNEpj8zRR
vQBG+V9U5ojGnN2PkbbPtiWQZ50ivxJSShpAJhxXYJcsnmeXd7Bb+jA1j6ZL4/yY
Yy5tqXBIDL/FHqXwqhuZtGuxQIxs5pdtGBb2SfaZs/ZSobow3ZINHijfIk0EMxGV
MhmbRVkcSlHgZhSPXT3KoaozOvZ/rWDIxySgTr6bmZX1qScI55SKLFIuZZktIzFT
FErzyHjK1gV336BGSuCUMtGbzWGZth6l+mQvcpr+RAnloCe6xQzLnblo0Xb44bVw
s/z5cji0yFogZn7NYp+uS4GUuiU+s0rsaNWZjWu8RxWfiD/ppLZvMOozX7tFTJsr
DyTeGmReAu+CwSuKWD0wFkPpE3iARCkgqEDZmaGZehY/g3cFgglDDnE7pKEdFA19
SnJCJTrIjN8JSJiPzBbSlxIwi3ZNancZ9Sx/jcxJYvCLzXlhErd0tPH2LxPDtK18
yi4njDvp8cvkKIEkW8T2oHPszW/4ktRGdZYV7VUKb2SdU8V5SSEHBFQ3/iad8mF+
lP/WsI5INkVu7eE5c1ZtxtsPbA2pbikl/GsmCIF4TolIHzYNGcYWw6iIsKFUF4uF
jA/cDDcYs6J9eAP+vZnLaWLrzCqEEu2avXwhtvqiYJ1yVZ+wKPgw+O75EoTs9T5w
SAXPWrhmHOweYDZr5f8UopsbvfsL/fHQoDH5l6PjC/WLO0JX+XSOQhnHWSSBR0vs
bOKief284ZHKX8ksqZtUWKQkmj6HvHr3OB7mTKFooh1pPQyjKUMxWQR9a9FW92XH
CONQ/dJxyxNU82YNEo1I008c+VFrQx9C7gfCOvk8uaG71AUCAbA4/IXwwO4t6JCI
CnaSOwA2zxlwrtfLYX2Ykwtq3WutVOOqUeYqEzxmUcEwO14bC5RJjLw/dGeqwe5x
7pXkxofluHyj3PMczRYu+LvEL8YWOaP4y5N+qqsaIGshWcAxHnhl5Kg0p0lhVObE
3H8SNgiWCXOgmWU/EvhixYBIHcKNNW729yCzPhRDIXJmvQiJGDwi8d/O13jQO5qF
0GkXoHmOKZ3z78apq04XqPCJ8YzWNcwqXvhpp1fIgaNp95hRY6627TJhArjcv39n
QUDQTNmImsSt7RMYWNd86+B9SC4IDaHEtXKJFvVxKLvQOmWjFR6O2nV+IPWyA3Gi
9xa/DWRqPsz698of89t/ABIjFw7Q16dSp9l/q2J02G79+dDRPiwV6TmiogCLUeTE
Sgy1hUDbMSx/usBpxJnAkEWS3eOgAtwTloVCZSlKAr+Iv6MReWs6FTswkNJbDSWA
1UgL+DpJTltH4XwvTRNR5HZimkOdZ3viZe8dUKYDnqPAPI+7Hxw1m/LurVsyfGC9
DflL7RiuT/WawlfmZ9gEmdN7O1R7Yh/KUYDC4l2GG8pvtbS2Z6DX7u++lJVlsvi5
ZUbHjX7ocEewNOBWvtr+rO5BksMGONr2EZuGNvzOOeY9ZTTi4k16P0iR+bWNHiqf
1Ap77S/vv9EGo/CXQTdSMowDkeILvg91o4uGNIumGqK9sW6qr9d6mRbeaaf21+bv
fFwK165Aur8vnH3SCwLmKsMNec22bcHetqWlItMveibRkg/MsLCYI8r7xzxfQ2Fi
AgXC2kt7lzkrL/nw++UYH4Gbfu9u81UQDUVhVIg7I2yY+46HiSM3h+j2xKB2MZov
7Ou8Srrlv8wmNnRPRt0pzDgPOXUQw9qw8w6DUbydQARsLSqR4mAxuimRSwzs1u4b
OGgadI482LfNzfgQWuNReRv+6M57NBSPSEC4WfJYsLBSNz2WCAb9/612rioQow1P
HfZedZSl8ULjwf3udA7bAwE1ZWEU+ONtRnCzJtDXtGAunr1wJsa6G9gtUkflSsDA
eoZbDrO2A83Hgwf8wn6RJnzIJ3EKFDXAMSkazxXN8J1l7wmxkjrlAcYwrQQlmXn4
wy9QAo9L8slOAqm1xVwlDbujq1e7xFPTPw/fzf2T65Rtp8PsIt8iLoM0Nu0r9S7H
4GapeG2vaQQhFTaRAg8iYgOg75F3zBnFLc1+y1PBzl1j2Tx7adMCMMCe1k8/Lipd
Y0nPuAdfVlWpHv6dinaJjdD++2TiJoSpeJbt45G6Slftru6DncBFaS2vznlwZjiB
z70YaRQa28nACFy/ONqy+EM/tmkDHhNYeKr+yJbgkvRVq2IboemUf02iTc/1UP17
VIqSPHRhNwvCX2ajD15133AUkZUfZIrZd1pyXIBPolPv/odPfVWlX6Ul7DxK/k67
VEGVuHAGPSjbpzYLsYI5PiMk+dmLlzkLl829VRNLWGPy+knJmOrJLbSWaxkRhJnx
4jG4J1WZF1vDDyKIZJzqHBWLGAGdPL3B22vjSm/UTpF4CRmA9gHG7BAwinSuTt5J
BmFzdTCbgY+zZw8rcWuU3J1G8vtQgRKxficSZ3NxfhhYtZwU1OwixGV0LzDEUiVn
dM0kUvc1A+VhGhS5xLvdowNFqvmZsm0c6mJ3fVxifliopz8OxW+K0PKqGmAF/5xm
tXIibm74uTEv5FTAEzWX4n/vvgAyNjOMF6y+9KmJ3DQHQRz+KOhu9yl1MFYUiIS/
lHqstBgnvWfIxbz7py2Vfjgg1uUVJ4L5gEclfHNrEz40WKqjgB7KLBflOmHLniGj
2+K4imvUD9qujb7tzyCbwXXHiTs8BTyGDzMOhfDa2ZdMENW03eQm8E4D8IZBi9JH
bJV9J6rxBXqQ5X1gKn34Jfl/IBMeYzkwHFndfZqexluKiCxrK+gnIRcJwGNNbzTE
JclK6DYji6bvDq+yvKtDvnnfKvOycK5XyrzpWdOwkKOglT/qa2aCBdgY3M3yV15Z
6rMs0/oXtDNE4MTHng2C92fOzzq85Vt5RcjpQi9IIZz9A2R2LLqKcc426CiWfioG
MpEE9YQhOSnsB7eZARQmQdFCv0h/1HvOCw3Q02SrZyuMJaMusHkM6d2KQfW7zFKA
/WZ0AOMOvo/x6GqcByco3qnv+GKAIuODr1LxnYE/HPhY/4H/J9a+JEBpM5jmJvS8
u1dtcR7jmBt5ErpgloMeXx5CedeqmlnGOPavAQcr/goQEz02I2DW30ScJZf1xUHZ
S2G7NYMmoyv+Di/zuM8EIHv2IJ8JoOqR5IONNCdSkK219WpQM5KNB9lxbSZDsfRo
5Tkrz55fU1RkHNaojLPWjYXvUsXJdV4NpsujpWSeq0ZeXP/HbSU1sWVTUYsf9IrI
Z+9v14HSWrAdpLEcWLAgWHeAeyYVqr45xIe+6QxE2+SazFwNrJhnHq0RH27VyfTa
dpILGow3aaa5795bfLqxSjzyZMr7dgLCTh3m5LY+vUtKYBZKmFnCHRzlX+HZdLKD
JPYQZPqnj2U0urEu2i0cUFfys8LysVX4AZHyGYsrkJOEsjHVo+0SSnIox8cSCo6H
LmGEUapJSYJHCV+Hv/HPqQV+4pZvBpxiwyaKIalycD3TUnsHB1/l+7Bl4Oog9XRI
nsf0mkk2jQPF3xqRrvZr6hqJM072tjB9RIm0ztpzgQCAFVcXEhs1S2Xemk/gmGcB
M2Qk6Js0QUdiswTECu/VRrYnbXSv5mfEssvCWO1I/9LRbyNz79Pz2jvkGm7RODkG
WaCkG7Ikt10gam61r0mkPXsGPXJxGdSwQLAlJUtF9ii5UQL9zpjF+Zf8Cm6EwTaO
JQmOnhdn0Lpxy0Od+vgOZoHv8tK+cxA9ggqtQj1M5Pzqh+5/xDYDXXB3EpuOoB+n
R9R8Cg/V1LTEFPJiyVAqaYEhdIwz6IYPG0i184xp4beyWoC0kyBwo6Zz9997etaH
UyzPgI1qB43qqsqfDw9+K79TYBVFFW8V3alWMWG2ZTaTMDIVd02Ftb3NkIIIA9T8
QKWyBFywpddqHxvq1SEz56IMSQCGHMtzee+ibcnbZw9R5HVtgI7wOZ/RPYnq4qkB
Meomq4D8RvbboI6lyb0fVvPd3Kyl490uiFZaWWIMyEB/U5Y9j1cWhgt3zKQRlkwe
ew/ySf6VMoWq+NsJC2aMoiJKGDP4V4gcSL0E529ka99/9TsBxsvS88E8qOpt+YCm
AzBL7kISy81vaCyn+wMpa1y4ryJiL7PxMCEuaj2MJgp+1J60+P5WURUsobEwsVEm
fKkMRg7RCdOJcsRrUO3YvEG7ltkjzqqKTXefY7IbdCerjjZoHzCWW7PTMlm2bUwO
LsMt+T1ceqGCPq/oP3ZuraZ7amLu6X0sqjUZZw9TlubWRFyEbsA0nS05pdw/Xxb1
xpkNX+1EmMkOjo3yweXT6e55txgGnDsEsI/IJ+7GmUGM/0NgQhOoLBVx34Winlb0
1OLY3dbFHR22qdlwClWGugttlQIOU9XZ7QNiHsam3zuOoaByNlCoEb+wZv2p2Pev
Z/GIfSPwg8lozWB9q3/65GFEnuMmIqaZWhsoYCpPLg7ERC4OGV1Z/Y7G97HfRDU0
X7+gDHXziLYB5yhwmFv6TER4PLW747AEwcYbPlXrpCZpP/JZDdeJg32ubQ/L4aNv
QS4cOYeKaiBD6m5mcAmkjK65lgKx1ocJjGFHGQGMYKERRDqfO/EPHtMWviCg3cyF
bbRwXGWVMA1B5eMqY+vPz+UlxXU5+wODjD0Ytv5q6v4nvmJXYlZW3CsfVOFLYjGA
wKPyRkRHPU0v6Mx+sKVkQQShuJo7PUvnTlx7jTG7v/MJoEk6W4AfBbaSxGdl2p1u
igtUo35hfwBhlgaEYI5FVKFiQu2BdXRpJ8U5grbT2KlsnKaEc739GAQz5GxPg/L7
GPUSspA1+gKGHRrypxcCGMBGMUIrjSOOTC4dA5NZiUf1yKDCwx51+vYNPuSI9Eoz
n5Vz2Bv/AuuNStkUSn2tMBzlk+8LJmqy+yU5JHqBa4GrkkVOq0hFVsrtcpkGynbM
SFBUD88AFL325Xyj/nre0GG5VdEKa69eg446SlVgWHDNpAJE5ziGwQVLOCzdxb2B
34L92dPigzMjd1bLftGTHDHbsmG5FLfun3NakRpCyLzpXdYNi7QygSicdkuOpWQz
vVCKCG3SPHQuNCJa8nbnXzfuzkdesJRIhpmK+ziWTwNPj6K36mJ/bvGwgJg5VHL6
GwGHC626OjmHe+PN/0gAamf6vJm2ta9KScoLBoyGB0U7YMOIPn/N+KF1bq0XcvG2
2LbMr9xY6w5FOwCu84+cdNIZYNjPx+3L/a5FuTyhMXrYFdfiaJqIts4Vhl9OgsRn
L5fEycjXSiIH5YUJKpvrUPwbm/laiiASP6CbvYmvqN0DZ2ZtJgwzi2C2kEaL8cH0
k0lfbXKVvH/vqIIZIbBLeNOj6XL48NvKSYq3RFo2E7Is73JiZpTZ3BjTdrDof8bM
b5IRiSBWfdeE6t+aUECwXDLjlv0wxlNtOxvC5IteO5vHIFCuxBh8i6Q/jUJKklr1
rGNauMN0IHfmy1kLAtaYAM44+yjq/tWi9GYkwktkaEL7xTRQp9YbQ7jKIpXG5Yij
kr/MFGfgRWR92si8oDdbpb+c3pbWGPfYwBID2vZi59JoBHZCXlgIsSuDdPuRVfjG
m90OsRjzrmEkmC55g9vnUHFjbN3oAGY0+jVHNUcKioAZZ+EedlvNbH+PheMTbqNZ
qBbWgxjqqNxUvjwlZr6Hlc0/dxT9F9nmOystBCY0N6x/X4a84RYxn+XuN0cE6hV3
zq7GgpHuN9V5o8Rd/bcP1D2EGbXdAPli9mzmsAm+qwNCvxSO3dVVBddyP1E7D0rt
wtuuwAkUMoNfKyl+KPaiCT+Qkmg0HMu78ggndrVUUsi1FdCyptEop4cyC5CiVMVN
xYtaFflhi6cX67zzHqPjP2R5TLY841IPl7ZKjyCBTSCu8TMywK3RANxSfa4HZqGj
NbXRroWT655LszAN1FSAE21YTDqKtcCJzLf8Gfdth+k6HRV2I+JD5xqVl0OQGw7f
A8f37Gh2U47Do88nvyP9V5u5xCHipolXQnEbxPJfVwBbSR5reGvzZ09ntNpLPR+K
NIPqajsoL+kHj/uWoqmDX12bqpzcCix68LdZe4LEXEAccYR0Q1nQSt9KOJmH5xqg
p8695AZZFroHN3EcXDzKw93rWsBH/U3osdregOUFY26Sqw3sc/ovvsPye39FOmxJ
5IreXV694CQnV6PT5YyQ7rfYobcNpMhPycJRrt2I7aHdmmJtiuiVliegjv4hecPf
0I2U4H90X6cFnnaK9aOTtihKGgcv0ZJEIlUsOy6SI4dQ6V2TSwWbFAD49MC4XCho
jytlcHdB5ckgl298rgHqDUTrwPj3KhC80olV57orxnqemr/pnnI14tZRKh6KDSNT
hGkxk+Y7EX5ezPqJp+yVaETxuH6O3Dhib6WF0wrG9wqP7/DoBxi460spv7Q6jzk3
SM/y77he/aIP5Lhk1OBLLhxPiN7G2qi8Rdb7QIw3kD0fwwagb9WSDOnThzYsSRPF
KvB9qRH913Ca2fMNf7AOHj8eX4O8yGXnLZpQjlkENwtTLu+z4JoaBuXt1+z1xxhc
NTvmDKR/ctQSKtjjH2RvUSdygNhk0CG9gXA009X6NT560cm3hWvE/MmcSCkvEN2f
UaXf9udJT4AzhCMR68Tq1CwKVgnTs35xzWWBLPHb68R4kwrAHh4bTEDNu7J0Zjm/
l/AZ54EA6L01Ts/YRJ4vMfs54Rs5MGUzMci/xtryCMaOjFD8zjnOpqBss7SX0dgp
2R0ehQXoBpnMXnnCSAwV+kfN7vW8ZTVL0XTdAA9HnTDuBNaS9ksT5UAONVgqjT7m
9JXCn1ZBgNqzXP8lRKcW+Xf5bvuCifKNWkdLHJbHhxAvmabRV6Du6Iya2Z7OHri8
IwH0C7Ol8lgc6T76EaNOran89EjXcQD90ieGoU2BeoJ3TpU4h9mHUIawNR5/+Fwp
+CCdM10YPqeYm2rReklU44851r2bwLJ24ASDLqWjDr4pPx6AkntzSLwo1GsgBBX+
5TSr7BDzFM2bSx2esx/AbhvT2+hqntxBr1BF0U2kO450n5YwwTXG8KgW0YL6msVf
fO3ueLMYE8nX1kbmUGld20LzykS9qCG72H2M93txTRxSsm5oz87mNSFDQx6+4hyr
RN3EP48bw0Yv/Nydx4vWPk+7tcLVsGZAC8/dZlhIgCCygXcDMJWSlEr6X1Jkz9c1
ij8AL6xnVhHkLVOf2NAqZbwIZZqTb3Yinatg6wBdUQeyBMdglcxUOrPG6kFml7tC
ZR2QzFuxd7c8ljU3e83sdGTXBoAZSbEStGIBPV/N+dn38XmMAVRc279m2EpBpGx2
3lFx6ooVOrf5OocOOFCDX5KMotGbiDiYmd85Wu/aeTZB7PR9VPEymHrV+65vTgO6
aYYZZolC3h6Dw4Ku4g6dNKO0EpVcmDm7fCbUhHkhrrL+slum7QrkebtqrwDcJPLr
8SCmyM7EKS3M0K+GIu401RHPUGqb2+WU4VGdIvgXT6StluScWvBlq7ZEUDacm7OB
W1J5GLt1CwMKcCC3sRYenu7RQd/MZuWlqQkfwXu8OX+BsN7Yszm3mGs3bjCBhQRS
M+KenZRpBJBcJFKP5f8Sn2XWuvgT+Jc6LFLXTtNK1R88lxGT7lYfebOaDQWZCMpT
okEYZJev0DaQavHRLTUxzjBSFNjW7TNzdznOpwALyiLm2v3eOmhLwiW/kKFJwZVk
y8DDLrGqDQ/w+VzTXPTXANOci7G55sNn4iSF/O7PQUYLQucQf8aV4UZlaPgliUjR
E7aSEq5V7EqA6c5w4Al7cVyEZjNwdt5RwxyA/61qShksV6aur0PovL1WAE9/sXqQ
Wmfepnuq0MQspaEON6BD5IuNV/WjLon5OjeFXAXnSskHITv/epQwGrkL3VngSbvg
LFg6EIX0Qb5CrrGsVptFPV/pVdl1jKjrEIU2p6gqU7I6ODy8GnnQbNCwtZ8KRy0a
qQpv2woyY0NHLEs5hailInAza+RvBCdpWHXJ8dFpq3SlHWoLTu1SVAtSfVaEs50f
+uqqRtof0fI17k/m2Xbxu3BowWGe3w9gtET5FJVrPUsV0ru7N8iZ9EDDMXITLHFO
MQhxYlHWWVZW3t2DxWnRUC7gdhcoPmKuhx6V9S1B+nZE45KRu6Qg66WO3wn2PDHW
L7urY6UFwmtbmW3veF1m0DsaOcBDDTEqkSDmNNlaMQ1bvkqvXD2fPeY25RkhlbI8
OncnLxScvYtIdRxw2B2FbIQJPwBTSBZ5Nr05AFVwVJqp1MVhwPgVlSQHJi+5No2w
sfvIG/Ljvgj9Cgt6xg9pIPgh2oDawvsRdhUN8get+tLs3fj5SE7JbyCr3Ogeu4KX
blLggDmWIFOlUptbmiCzPLj0fSw4OhosRL+tLp6o1ZBxbrGKAYSau4s5m7cBhYqb
Af4hs5yjVp1Fv4hMyq69WZes5CUtE0hV13cllDjyPku6hubgXN+bA9syeQwRwk4C
2Hes0mX5eHyaO3Nd5ptV0Fc0SfDtVP5Emq9gLGr8ju1JxFSNdRoUzDnBATCv9Ion
WRECgQ/+pHH+wkVr/pbKkU3+ggFpDHQwZ8Fzup5YyAFg1mgEycPndtfOiZ6J3Hmc
wOz7AsTn32sXRlIIVpkwGj1sy7qzF7cKKvOb8zttmDycceDDjKxprO4ojKxVKxDX
rYYJxj9SWRBXfLHzpJgf0sY142SYBILqkAGI3fyxcIGeSbKidPdrfGoRka4sxZYv
meLkzEi+1HsqX57h0c885ySKqmZPt/fRR2ZphKwVZR4777l3ww/bXcNtOBSr4FiQ
gGkZS/93OsnlU8Qx9KTxd/4uoGD2qSdcY1jGmPnJkBPsKOkEeV9CxcivZkrFqkrv
dQyOIDvJhZWVp/ZPInmWMarJ0wuUiw84/Gn0yz230cYzYr1e8Utxgz0NVWyXSOEU
DIbb4s7rwgD07rss568RipWIaXgNoonLymxrI1mRS0V8d6H8ZfBWAi0LGo3GRwzI
+Ao3sfVSNW190FHBtxOPlNzBNbkpe2Wy4tvYT5feSFHG/GWzOFB8qY8QUKHfXw0m
/v9x7A9HHnCyoaxh+N1nAF4m2jZdZqFfskDp0TRYWC3Z3vY4lsNX5bdLq0VoturE
e+BpI/86p69glqWQoUKsGyXRjXIkeBFRJq8wGpocLIZdPWmOMuRXbNf1MdRaNrTf
qsKoDZ93KClF1Fy7gvCApRIyM3X6I9xYfhc17tRBYXVgsHNDM7ibVg+u+ReuRFt4
8eqd9TF4M+th0L84jabLcBNUjgBKIpuBdA7d+epkKG76dlIyigWTQwiiREBOHJyT
zU3kihK13gBXnzLQEKD/dWZtOFMZYMvuo83KEMZNwzhSvXup2RJpYRGPkfkD3sCQ
HF+5h2SDUO5W4FLnYaSb82mN6fWK+l/nYtWsuc8AipIxIgcX+WdSaiB4eE1zRWjU
m8waRT94zgiNqtTtA0LPCJ3dhxfkMys/9EYsJvIcElN0ViSlL+TkiCmFUTOhPxWx
FymBWExgsZURX6lkwhBeYpeXZT5Me+6m5JlVFsvd//xu7y13X4Q+W5GpcjulhQlF
O0/cSYogsisCzLog+bK2ItoqWunUxs+UMQy76iCN56IiffYKtAMkvjb0P4JU8hWP
xmmKM9EVrh8JbHyG0KToI9qsu04xPRLG8vI+ket74/ovkP+tvRtuGaUrEOaf5YNR
+5igIF3RXmZrwNsFXQDN4iH6MZNiBzW15eVm1Kc7JeNR0v15L4g8xMR9pKYkV6zl
UaNRFTkYI1wBCW4/xsWtGxFJtAe/ndZsp87KBB3Ei4fzo4tjMOAr9stVHuvwDogj
B7mGSAsmZIUA+GIfftv323P4Eecv4O8HU8iYrLlasxsqHgxJeestigUgYjDQD3cm
vbkBxkpSH6wtrhxPTe422j+383yTSbFMGFhYso4gld19WJQZ0og7/jVK0ZfIW1zW
PckhHtJEtg7o6IzXQjFpskgyq/k4ZhaI30dB3r+MDp4nJsWMInkFtfAbT07UKw1+
4UAoRz+9O+/23FigOefTkmOLOJVUs5JjViYVKUv5LlxGY/kICjwxsIY7tT8WmSVf
7C60BVhVKytIIon6APxp1sdCtAO9GKMqNOEYMAVfP+65B1RotT4QAJ5FFam7zdqy
kBLveIdTvOTfCg9umre4ax7AhNvVkLmntad7qUPAKP7Bg33D2IS1FMgYaya3ycsC
PmZoVSFz3+pT5yJwHZCB7tGn+PbDfwcatx1Hh+EJ8yv6B2exCnKX0QQ39HZ3i/Zq
42W3c/BQo5RC7aEDadwffsns3M6O2JwefUEB8aKQruMGKjtZJOsFE2tiFD6vfevv
zod1j5SAgOFtHvzR4pNnZeUpAh0AnfsP6TBJJaFcAfd9AJPxCrsIKdnTkDGLAf0P
JeuRDZKLPgIVVoClaXjWYlE2l3mejmMm9pBdcih4dImWF/NwVvwrTWYuu4FRP/vx
eH+sRmY7iYiJL3bzGVETLsiNENEbLfC5EZzXJQ4rDkSHjeK090pBnkMrzxKWnrVS
ItGZY6/NAOcCUuhypMo6OtrVvhq1LYEUN2w3qrfB4c9nXFXl1PIr3LZdNT/UCyn/
ayAkTavyt+1F3dUSsinhQWLyvZCCCihAoQHTV5b7iIWThxG+a+L236Ca4ZUtDPNw
imPF2SnCQ4z4e81EP+4Ola8pEw5pjYcJEuvwaFXMbyLucKrj6MBwyOL47cE/3Duv
vgXAvUi/SP9z+oYVDJ3nhBnUPaFRTEYQq1KQIXOyV9lqTBmVAjsOAnS0eFBhT0h5
V8s1oPVityYKDy7V+s4ccIKsIbME+GswRs1flau7NJhPeR86xNGAUbqMJEFhxZUG
9NL0qPgKVJ2jWg2m4LWnDYL5BFjUFo4pJPZtMv4u5FwN09XuKWUlSoT3PlABh0E8
qgnVJ8smgExys9qzfyMr/LnCxYD+xIWoRigBRXUYbgpPJiCKGvpCwb+jsK5KRRm+
E4PcSPAuNEQ/cJb0dAwfJWk/7MDW5xHnDFj70Va7NU+CkEfqZK561y/mDolUNRG2
HZZDJn0bzvVlWQlKL5XMqY7Zyrqig4lEX8o0HNA0/Y/f9en/e1wuiazWQDDHOcdN
4zMuSNc0krpFH4CJ4WYaYt8NKvTnENMKeg0F77OnOMIRiFbBK8psquhA5t90r0bW
QsVJTItXj12T4Z/LtsVi6EQUVO4tSO+X1hDx0pnEqfmrmnBZ1JGb2vD/LCbssH9g
qnuqDlby4b2cJYQaaHcMH9d9wJIRk4PG2Zd69WFYGtt+r9iYNyNIbjEjC8Y77yNz
SV3p46sn2QSO0J84VAE9XPLHxuxHyR2HAqfx4sHUp7hgaRrsjjJXX7Mh9dFRkIgf
X6IhehTtYWX1jwkQWzZeo9bhHs38z1CtsETj9zQeE1bYcfeM2K1ZcEM1kXAaz/Tv
SxIqOc7IJTIfyRDvB8BRZYbs+qgVZhkzGfOaPVEhGpIwPdJ//f7rSPKnCH5Yc9F/
cTVg5urOZHOCoom1J3vqo5B6qWWn4HTt0Xlv49+74hvtJiV9EqgQDcye/8Xo66X3
SBs71HZvALchVYw0zYubVs5EJc9qpDru5EwT1CL706I1gg9nSia8szC5jzMIlRK+
E4mVvAl3FimkyqTmC8kxQncng1iTMDXHMVTK63/1zfD4cAhCBxYJ/3yJaWFR+VLL
7hdRZFJdv5gv+JUo4XkkVq1J5Tp8boPMuzKO8gB14nmi8QcM+wANPIe82KL0sM+C
zaGn3eAES0jMFpavFKkyc51fRo7HLgFssKI/aQeLwFNAhNBE2JDFUgGEkFK0IIhV
kXFwiFICe5KHO33xMVRFG+FGzZlRrX30qbWy1odZAuJQJf0HAYx/8GaV+EyZ3LzT
ZLcDX+OhjrlTs9dket8XWbkShcDf8gb8kHUVt7U7JVrrPIQ5dqGj5LvEhkCFQphR
RaP6vdLI3pJsUYal+Nu7lnALOyAFY+1rnML5kJcDk1h4cBaFtaqZ90U7pIfm6Ym8
/53+ew3ZEg9lXNq2gRpfCwI3sSr7BcQ3kH47YI4u2pH7+8lbk7yxhnijQYZOHD+t
4JZXCWNV06XgOYNTLuPQ7qc1eQviD0Im0HWfybqaImVimORPmTk/eHFUKwHVt3iC
M3I4jWIoK5MRuYhxtnh3vUASdu1Qfn9iNybqPweQgSVsQaA+zdGnb/MTCG2NXagV
QNu0WpnbcejSRguAKhfpvCIh5e/LG6N6HhibsQOZlBLH01/Ux2IfwgF6sX9uXjwB
Ofm7sA11JGp1wqBUDOz1we0ZOaceHpDI0YfruBlH4Y7O+5CSgXiOcl9l8u5Q2uNj
/qJWybCg7BkLfyE4BI1sMc/167LV+/5+uHsJ5dX8gyY7ShUmUule+CdJ0Fx2ZSTC
VnRxdutKNBwwMqIEKLH9oj+ODs3Q88Nd+dICSMCcSuod9ukb8riNnt/RxyRrjri8
L2ZoJ1BNThOO46gdm4Gr8/Fgbasna8909KPCf+NT40KU3cfUB35oZUhWffY8L71k
n+rzwa358ZIIyDRj/uOcTTTIKlVNcNx50MbcLY/uZFtkTfHS+ZG1AvMKcPH8nAu4
Nre7lvq2/C+hFleKX3g+BpHGVGEVjd99ESjtqbGQJZ9FQ0aHsJnXMrLT2DhRyXU4
sSSXo+Jx0/I1li5rwq5+ayRm7q2hDluGC9prZmxr+yKoh7plU1b7SNDdJZ/oMPCv
ZEsDTGeTZO5aM44k6XQ0WNZ/TiA24tU03CSd7LIPoUF27BsjGu8i5EJZpOJTooaK
IRdXjkrv/y5NsKgEUc69YU1/nZlLZEDcDJKUQrnL48tAHJtNrT78uQdFH1jGGH12
xk8HCLoW+RERNaNigpq3bcAApx2Nps0MyikZKzuAji/8/XBuCo95I61hmEdUWqDv
m5MbhezVHsOBGhCN9oFR2CI3DPpstYyRMS6VLyFbPJx0tAoYRSKzzu5onlP0U/g3
NDnEgjGt7dEgVMbz+ykpBMB9TWK60EQO2PKZxLeVS/vquQeZ7UCH398IyJ8OxPuy
q+IJv7WpMpBKqZM72GW+/6AUxNRFqMGAjNnx3ycNtFhdWZZvNTlsH5ODKBg4QGeE
VD4a6gxr82cE8Eb8muuirGXOSBbLYrA4jlXg8pBLgZ5mj6ekiM+7/XkAhA0MuXon
qOQUyB/uhMnfY3b9GHwLQaF8oZWO1fMc9tZ0rBavKIpoDKKcOU3q3lR6Eh7cpG1A
sgqgu+uF9WjMSEvois8gcdxV2QQbPDxgOnYp9gjyA7w0xDAM6tTUpLey25ufGfeC
8fyRNHPdUYui2M4WkS6LmuO4rVJG/cZ5dgYM7wYEtww/O6WRaSture85lg01ar+L
chaFtAKyhDXC0Xc9jrvqbKinLcU0Fd40QJKg3DjkBYRUS/1Xsr2nFMc38+yqALCP
YpWWI2p09MmYtXEN6hU1/POsnKVsQ/D3jHYutvQ2j/82/U2yj98N+L9xe1cIsqlr
zJxh3l7vEnbL2XE3s475Y+xfHsKtEtLfhS7wnIt5bJb9ssw0246sw1jVaJovNHsh
IP+QFy2TICyCtUib/pcuB+JPfmghWQMDgg1upzyGdXgo+FERD5u6POclGq/9QrXy
ur2c/OFyxrAl8fHanWZ1PesVePL3kXDIV95xeSHykY/7PENaJfDR3usmIK5ixFhm
ZbW4vIyJRqQF4LXtAeInhQan3h2OAarlug0ksDOR8ehr0762LoGX0yKFVbR+EMus
q3rZGqf/J5/pnjJ6I+YZS9+smCnwjLAJnCmsqZpXHg9nnZciG2oUEw+iYb6wlorg
aEGeYuR/9m/rbtHxTYXj/RD4SyKsO4UOTgCPrlJRFUgnvrc/eQoJQ9mrOAVa/w4K
N+HpAzfyMs9pKav4y+lG4WvOcAF30S+Gl/JkrRMcj1XiSEgKaqdt8CO36q+CIgFw
WcH0e4QwYe2CivL9/Z+0rzCPh4KDm5M89F79+sYOStcK5UDA9fF/NNjG5T1gj9vH
DCOU1gR/6ckT9H6PETyh2TCN1rvZOa+LRVYAx0kD5Aoi2RyZMz7q9Njm8S6kbb/h
OdahY4Ecd0MbvZFON2IlnwyEea3q0rYTXz5VNtEnDNs3Is2IYDqkTPF8QWDc86//
8G1uSj2uHDjNUb8L9wPKeAXkvbgF4Sm1fxRCOtf1/aNXEOxSxV5q5ftzlTog8Pf2
F+4CppkyZTBE7tX7gbn5lPpQziDCH44KrM5fXKJMLCpAO1a0YRkylOUoMjgqJvwB
8zeBsxuweShqPFBGXkI/hYovGy2Xepw4Zp1lCRBHeYRZNQbJvp0RZ0DIK5Rt2x+w
52T0A2+AKXTuvc6OVLKqXx+HxSxb2upRTvBOkUHlL4Fx7KB3Z+14JgjieylgHPaC
fYdGS9uloa092YQWPZj5HUFVycWQ8FZbEexb1uO00/l3z7e9dQ4QJTioYPzZz7SG
GkCRyHQylftcA4p0uK3La1odVBMiBMvlJYqylzX4JERwUq9qYSDNHgUuPlUS90d6
SlIF5w51q604lgMnClmovC7IPBpIvLLSG+8WmG/VseubVDZDJyDwOIVV3dtTr1vS
yLJ8BBmK4UfxtAyobR2xLSQUyXN3hZPUT6F3fw1MiE2O5yIUAnF81Jtqirz4ECT1
HGe7+FDOo7FL/gN27aV/KmDUznXCz6O93jeaoKqa6d1OhjX4GY+8J71I/D5/QTCJ
Bwz3RusAUKLrQSzX8CE0NrPmXL3MTZWo1GPIGoW6CQGdLR53RxFcwqiIf5C5W9K3
BExkFJTElP6F2KXBN233oPhqfH8tQpV8SJlvpQlPe0BCHaD60VpfkE+CC9oqq1dK
G/jJF0WPuR7Z1SMzAvFKOmzh2kYdCwEernAMTjefuIGx/IXKpITvUJdjONxQxDo+
h6i5k7im7sypIKMY7kPly9AmITnTnb3mo9+J3j7WFLzn8dW1/qpVxQ6oOvXpvTFd
NF8/Vonm3/2F5Ghge2T2EX6u9of1wROzpnsnpeBpfcAOpWZFYBx5dja8tf1O+Hm0
G0UQXxpNrAFSSx5krXgdRDk6DFEhEjJAdmp8Pc5gCINbaXpdvm3FjNrwFuMyZEr4
MvemM9brOk5dEQ0SvVa3T0HKwGfTJqntKSJYEJqyyeO658ystP/AqzhGxE3WJyI6
hE4/jitHpReefeULfESSSoHmH8c2GdXL1WDVKtaVdX9yv3jnHQt8ZemwqL7LGpgT
2UIKBQVKq6WOID8yff5+vHJDJwZQJRDhOmaySdPHGrPy7L712xubPAnVUWMrO4+Y
Mm3DM195xNhDaD69Jp3BJZTRV4B+Fzxl4gu2eZAYFHhVwsiEEHk1KfH/CTg38Dsa
fYo3WxCgUsr1ddStZpIuOfMEdE7KlDQMZ+JsjYGeYf8yJ0uanM9DvPRmWt/bTpKD
SU91F3038yS9fCqL0PXRjU11F2jI968OMASLRAu9yXKEIl5gDNXfYb4UthtNU7fW
tf8AucUruhSUVqJ2nJFihFaPiQMrPOvriCljNxvhRPNnJh1G3qeQ+ovZW8z/NmE5
Bo7e8ULTa97mytlpn6+R89sjo3C+zaatKpWINYzgC0urNsTU7EvhLygZKBeOIv36
1qB4u2p766izoL2qwCAwBbi87bZrTczsr/vG6t+QZZeJeZOlhPwTtoMcRiB5oVPo
/o+GJBJJZboIe0Cq4GgmHulVSHwI5iNiyo2WKbwHYoAbQm2YC4ljhFcqNszokkba
CUcgJ7GbI8XwF/7uGnGuXu5rE0Di54+IC6dKmd/QfYi7HxWUPBnUzp5AejCIO+To
+qBZmWNmipZtTpGadjx8ZJOcFGR5a592sjHbwjEKueKC/0SjYD3aengHY2O7pVDi
T/YQqceX0v1iMhgufWVqPiY4kUuRgYeNweaZ6mFHfik+6actQxy2MfOt6LJyAFyF
SOUV+yfShoF9EKJma0Xe1iarUX1cLJ1nubA2gQe//mjEKn1bdHwDhUD417U5W1aZ
h4vrTHfneqhyZuaatT+vlW24svbcKchF4HKXS7EDSy0oYdC32HiumjM1HtAP+8sb
lnuDy9SisCcVRBCgpr8jNGYg2b9e61U7kVXmFzYZTK4LRjXc8uuSnHntCWo/6zkI
xn4D5EmowZBxwDOqO/MAFTCCvBH6V+FnLAf+qRtwIXnGNYx3BErz6E3idkgc/02+
YAgOMj0t2yo+x7NNL6Ek4TFwavZ6StGwXMbmQ5DU0XMQZ34GgiPKnwE4FMGwMduq
0SWxwvuCXlptzAqaVJOqhry+Ixia+QzONUkNGRaiQIaGtYOkh/QQ8SKIIJVEzH5b
xM7aYb0wuH8deBsGZcH21Vc+Kt0L1I3XGO4HYWb+qhrhXEKhA2MjI0ilO252Sk3n
gbN77xTGlJQYAKN1LzHsMByVp8UaPD/iTbW6SD4Zymo98NvufVruJBEMw+XPOIPc
8pJFDllgCRJRtkh2JevvqLHV3Il8j2LtQx+zYw3hC64MHpCmtJsT8/6xray//UDz
QNsjyI9vtMachRcU2QJgfkWPYdBqLTboVHkjizAxiAKSkK1G13MyJWeFkd5D+vbT
nJZyj8C7vd+n2IBLHsqyCT7wHtMfCN9NCtr24nu+vFa1qp5SixvdoduJamiVzZEn
Ob3lx+STtVe0E8XjpCNTd1jvwkV2WQIuigfsM0Tu15z3e3Bzo/C7QLDNeGVEmvBn
tXaT+fXQ4cqvUkIi5znHOLM0YT48PQePlHt3ddBEdrio9WdOkLO8TkCe6+KLBlnB
jTQ1qYtpAIummbHYI6VOb88MvAAMb37eYVerDWpj7GHWLTVV9heOfHBbJXacIkbC
vPhjdSapyqZGUulEPyZTtMtoTRwwsgFzmcaFjrWT1AM+FBDgXseZYxFEN5ydLPqK
M7cjW5rnUy0/v0yVI+C3j/hAA6M77BZCe0rjTgnqSHDaJMvTukL9l3FXobca+TbE
luUHCXRJdLhrh8y4HIuUVu+iK14OuZ86/k/w2Ox2zloFvmk9uFIbf28tB+QTgGEP
giDFHkEw+TLkrw7rLxzkY0/gu2GLTsQHnQJ/dMp2lYrTEnoyoNLbtufyFXxC6Gqs
eVirtUMPht8YIrJFMX+SVS7XUszi1j5b7eJSCt9X+gZvBbOMmtSxzCom+USErDDm
WQ++xmSXrZllPSATk08Bi0RQAOQy23FmyiQIHOzrE8wXREUjIJhBS8VeyNghR5eT
Vd653iFEbufCm3f8hmQk24cx2k97vmrUUi/9RIHr09dUR6gPQ38ebG2oye9sk2tD
01Qr00zJfrd0c010JnC5a11/GZfCSWhjZPqB7XBr6h5vWPY4I9MNSWE5b1PGeL0B
jrURB/GWE/r5/Oic24N6hA300taQaSJHgH5nl7Qo48nsoBnSqV0onHcq+oaXC1pe
SMqS7WwlBUl71+PN1DEc8U8DZA9Ud/9QtVy3LH1pExz9GGLY0srpwluCVrTwOfU7
TXeVv58z7EZrQsWYvAxjJx6AN9GKgY5jOu5IsSeliXtc2zEX5i5iEjg+qzFxGOow
ziyDA+wNsqYRMEhRHSAG3EeENp0WPGtTiTIjpI3WEvT/2t0LWHdEeNcsziGMB9Vs
6CkzOrt7q/M4juSb98PCc008Vbzsh68TUWCNZvF7eGwsxe2GI3FZHVxb1KoWO4Hv
MI4VdfVHiu0HEmuQQMhY4xJ4fK9KteKipeLj33P7IqzsvoRujxHQRBGylVpfgTTd
N0Ex9wq9rQQBY5qVb7d43euW8luazh8xZrwFCx4iKc/pMztB5aTqxSQ8555sVHft
Mky9L4ygYWcE60yy4nQipF3tjuZ7gY0dQqVUHhI/qFZT4nO6Qlc4CooiVQlDJSik
ANvF1I4zIdsQWkmpdkN4ognpcinzJ4vSGGCcJ0dKkGwp575XbCmcL9yr1AY5/UYj
rXAqiUBtkqSuTQ4npJWWnadCnNciG+pHjG2/Z2v9scA64GtUtaVADj9uRymyq9j0
1pg4S6kk1FuPbX4DjE01a+haZSbmfr6sJls3Zi8dBYTP9YpwQyhkp2wNuLvyBTxS
oxmaqdJgZilHwS4Ynxah4fCBe40yPuGb5Nfw2n0RdAAF/ITa79ogszo/6dNi6avc
GQQd1JomfAzlpOazlm2TBUQ24OvB6xuj9ByWLGI6yKn5cPBzD7+cDs4UYTcJ/Swn
EYHkpmuC2N7sfAAwVDnFvT97wyjLmCqluVE74bz1qw7NoyBe45vgW4TV0jiRUyBw
TVtkdBjYnswZNdLhYgTpy0SOtghS2RFdqpWy5X6pS6KiUbnXETkiFbFbXd9RC3N2
JszhlR5SRc9O3syVRzqNTiC7kMmA/vNI0UzqINCX9sP35pJK21HNmT6FMErOaqWb
V+Xsdh39eAUmMpTFWDYn9/77NXcoyHiMWHGqVqgZ1cmUBbkKGWRE7kROqWYhVnZQ
GaAYknXBiwZrEOAEXF7jMb4L2E9nQEJ2Raf/PS8eykEtYRzP5ogz2iUQydNu3pf8
q0Azy1I9HV4A8nM+Q3Ln06e/piQ9QmUDUJHVyskREUX6LQ0XYbjzGxy52pUFeIEF
QXG0IjEsTXpQMbIL9pJbp7qQJdUkxPLFZMbJwIMl1TPgY6UU3Ftz7YOXBFby/qfU
k1mqseSMN2D7Pu++eRV2NqO5/HZhD69BfqjAw/77h6YS+vmR/kq186sRInw9L6VN
kM9291AELJsNTn0SgrWDRwe3UTXfWOcwprVXwu4RZGrkIOGScNnq+u5FXjEfFXXc
x7/VlnhmZ3eeQSRFj5yi0s/TVUH2unI//WDfU0aFXei7iUrGFkIhC7o7peFCkJhZ
Lkc+PxouGa3cbTJ0sMOsA5qzI2O1rWkeGrota2Qtl2qa8rAConffeqe4xV6HZ5hR
gb0oql7aEEe215355dhn4Kl5Hd+E6RatOH7WKHtMYZ6xr/4aajB2WUQncJCb06jk
JctsVzOxAu5/cXR8/4BwQ3d91hkXR6lkcOhzejZ8K4boZgiQbWurXBgsJHgCJ4dI
0JcDigUMc1l0lrZT8qB05v0fMsFvVS4wsowubhZ/QFfvk+NQvYj+j1PO0h5BuLnE
df9VWja5BBk5U8echES3jnp5dlmaSNirX/HgI3XvPwEBDrvUl5+c/V1UhfVUQhNq
1RpiqZ62TCh7cBmUaL1QSOwMkTC/jyiGOx6g/BqnFHeW08GEJxaPyrNh75tsprN0
ByKQxxr9pRcTOyYkwY2z8C3T9gPz64bc0IgH3mPTegovzQ79/+gs961ahjG7cpax
9XOTiXOViiee0uyYxhBROx0E+7XAqKwwFSYnWuBwbiQZa1HkZOcmYVJ9ZP9+UORN
3pg+QiOhpr49Tr4cvnosqIdldAKD49lK81HcepwAycrHL93zK7HqNoslTe8IL88m
tpE8GHRsQ4+wriuIJ8PosctG1ckPQjyYUefFanAB0OSDKcfikyB7NcAZfwjoBKM0
0r8AvISIX4H323hRXXx+defJ9c4FxWEee999hxDI9oytL1PkIGqUQEFZ8vQf4kC+
ip3zh5UjU0tyUvyrqqFQVvUrf1fbr5b6DkWkpKU4gIFK6EUWjQHsx1/QmEYNviPR
BrpLkwptVrC2ewg4IgOxJ8lWWsQpWcuK9twwtUn1G9yiNDcsja1QT8QhIN2WiTUm
NLwaU9KZM3vPHVaKgi9ksXqrzouIbB57HcZrQlImmZEEHsf16B3FA9uinw4t5vtx
ccBokGJVgjdOJNaxrgsnZh5tacVyZue7sMiGqQcqK+2BNItUiljsK2PMyrp+0gRv
Rq4UVmJ0SuEEgzoedOzHTMBKCRk0LoJEPpw4gvCpk/YrOF7TyMh5UyHDGR16IhMy
C9EF2TGmGdIvVEqtpIz6vb6dnghYpSpTG7p4R9F7GU2caBMfGHhNPdygRkMeOW1P
+JinqZu15X82hM5TBjM6AKVyjR1us48Q253spGAtDMQooX9KpGO6JUmgjLQAhoGe
BU7bBclr/tnZR9oTg2yUWOXuHKXUzmaN15TepAlXkfTt7+G2QeZOy9mZ/UUZ3Ska
zUx6FIrXLJ8TLGZMbcGr/r9bc/qo3XQTJFlznrFuE++yZpkUDKnGZ7MhiVVR5t95
LM6ceHb8i/rh1q/mrT44y98nZNf8WPHwcrlBXsrVcIv+WscFevlyAkxPn0yL0kYz
VifXXWtTmz1U13N6qexK+zYTdFWFYMgjDN3f1sPDQCghqpBSOArlaHjNlyGUjnTX
7UU/Abc7U9VuhDVW7Rg4ivq+TGWJNvPInamrdKc1XdAEveJyCJStgrIoyqsRfwEC
bqON9t7u6MoKSHgwOUamGJD0rnyW69KUaVuNuRESA2TfygQdZCcxH9Wd5tEpGsJM
ICIXI2B3UpO7Skkh8ecP/vTP9zdOlg8T/JRIY/enm9qZxeakVrSPNJ5r5+JxXhmK
LCHSylMycu5vNv8FvpLDNJbQzPHVKatpm3G1vzvlsfA9BU5dDxefyOzsWUcTdBk7
dlaGQjGNpFN9EfQUO2xGMsNs9N06J+COqmeqUNkZrjHX+dlngb+Fztm+Jtn7GImi
7fNkX9YRC6jw2jRwBWZdAQllhvk3t5lubRu9ZhDHP4tItsV8E01XUSbRefwUCDKs
7NKAnDeqvG6R+ypy+aTWRNrdcgU2Icr+IwGzqQmVg7OwFEKgB0bKE7NoF0d+Av1c
yM4bFTRuKQRqhv9q20r6OQjTNYpVKyojc/6lyPnsqxMBT9UJNfDOIF0fxjF0wQqT
qGOdPDHD65PI2r/Tw9383oSH71Int7/5jfo7t9tvXZblcjxYQRHaIUrrgTdpabLx
DOWjsrAbpn+r/6YzySxyJLN2RwjyCckZhPK1RSyAp27bWFjL6UfVL2HOAmR7hXj+
KpH44q4eZi2PwZ9oeLGZ/mDLnRmT9ToLnJLdZQkG8+Sea1mVdaHr0zRmpTGrjvqq
y91yGNg8Ice99GkGxVVa/0ks/90bF1SsII8TeLJ2m3xUITB0X5FzF3BU8ZkdbOec
oBPR1IqM6Pjnfzsbjk1OryoIxjTAbXA6zBn5VTNWGI7xeUUdrZ8To5bgTAnSTMEl
MAZ9quix0B6DdWMscMrmyJsxXDTSoOBLuDrcdTxgjRfayd7b8EICBng6Q3cjr10l
7eMbnnFEIDJnuEGoK88F7AT07gaXETt//dyXYm+6JgVdUKNKLkt5gfUbiF5v1gVG
HLSxLC0gj9Ztl+FO/FuQRg1beJUCBAm17+YJY+HgV0808vP3oeKZQt8x36xIfE5G
2hDD4KW6PCkzmyI3tcl1iJh5CDMARPArcoDmmLVl936uwT2eBUfHrBSDpHp+KY+Q
k4JFxbui6MA+3vERfcbjel5YVCmwuh8dWQ3dB+RBaYq1z0izV1d3P4uaUOzDcpEA
Ggd6RbPj4bFwwF8WwRK/akCNXZKk6FVPIoLjZ6ePHx0cn3BQDz6bstU3YfS2jAxf
ZurZr+bWZCLDNb/lJRwXht3hqEN0WNXGnZQ1uuO1AV3V06So4eSpqarYgONVdHj1
FxMKL4v6gyr1/VeFzLM7tQaz4PnkO3MIr4HBsqJPmBUZA2NuAzafLH86laN+CYJ7
3VICIWKoakCy4kEKhShnZV+vuUxG+QrIc5yVT5W0Yv3WUop1Czi/Qo/KZfDuMgZ0
nN6ROPoWsBDKiLTR9EuN4o5cXIFrFeiEbMm87sKWum3pavE2Bjk4PqcYZD+ElhrL
oZrkDAWgWFtzlHPWjYwG0ENZrAVGPnkdbHEm9aqB/G+XKrXjl8VhpUZEElKFiuTO
AS903UPXBsghipNLKNF5oBZazmMIIWX4DuhLyNpSQUMIPwiDVHtntmoQ7LA1xKex
nwlqANgEMDH/q0GIBRKr35XfY/G/tyesDxnDp4K6NTPBQqrDjppEdueGiuEpF4Jq
DqPpbCTDzarDWICvjp5Ng+AGJbplpIoNQg8lGrHGNQPq3k0f1P7WkTKOe0kPormU
10lmcKvy6FmKoWICPg64ojFkIPsqDPseRX+H0u/M4oF9QRDrHRxHwCM3TAIcN8LH
5jhO2IhSymTnd+DUu4JG/3ex88JE7spD7oT0OhbpUDOIzZ6lkunMCKdbrJbB42Xz
MlQSgocyldre6PRE1e1ckW058F/ewwX921J98oA1b56+NkgJikScjTl1eTb2qS80
/t2fYgVLsbhtLGSY/LtHln+0oqJebql4D0RQoVRMHdNFshdn8Zij8Ali9LIOrQuW
QVJljreJNLU8zvrjFNVVkE6Us1wB3b0KhhL3Avz9JYSPjnX9d50MUmQ6+jkxGA0n
bWd1AVlrY53scwV+QRD5ZzXyNlNBA3jIgE2g2KvujZrjWuXGWC9unZtuZcHQzlu+
w/ecTdOgXyswaQICGdec1MhT6a5Ik2FBIcaybGsMfy/grTB8aBbWT+sWnI4bwErm
cJytNcffdH4iW/Jc6mWzU38oBt+KINwqQxn11KCTykT5rMOEvPG9iuw1RZi+BfJ4
ktNL+G0cLv0Oasm5GlZF48qtnvfvNfj4Cf8PKbBq+nRUb0nNslcjaQRykNVA8TUO
YHTmELFvVwm+q9k1Zi1NGfK9ImDu8WbWOBFShQRFqdKHvG1OMFvaJYOMKDIlZ0jf
seMe5TKnIk9nK+jIFZvrU+NiG3u9U0PpkGi9YHRQyEVTUhAU392dh12CbDcbAZiB
tBhuD2KmeKHxZTBnXwmUCY9X9LFnOB3oXPcfhE0+E6nZY57ij/C/vkFNWWOnAr9M
QGP0dWYeLp9xV13IxR+JQsE2KacAzcYHBjVfVCNDWv2BOg55wyIUnVkaU0vhM33t
BpxPN/klUMQISmNZkhnr0f5Uj5dZNTjCyQAdzJN6flFopHv5sEQHZvYl7n3U2SDh
8PAe338CV+teWgyzVIP2AlEt0D5XYiRvsujrCtg6acXulN4E0ZO4YAq5U7LMTInK
ijSWhuoCaIgmBHTbwEXiv20++HhbtLKztW7x4jFuEw54pYKqy+wftN7bFJjVF5D/
mNFYNfricLIB2KUGbwAxMPWsRMc0LshvtgsJcyrbXTCt6usjewhVB6lE7RFfZzie
78YDJ5PeMCqByzhR0Cj26JpM/9vJvQWx83ExXiuBLBDMO6SE3yC7DoRt1yXH3nLc
VJx0SQPGB3fuXPdOTOp92akrBkyFaG50Il/Eb6HbhP7+Av3jHGsD0LDtGlt1J9pG
t6BfJ9ZQ/I4uyTiO3VXDtXr2qz+xWI26mocA0V18dJAYkvSvMDKhP+HbSkD1ySLn
a0A6EEtA+yNdVQRmN9Nj0IYFISYPigLQlY6uefa6Pu1X6rR8kZ6lHGFsz8Tys+AA
Svf933ZUMPuzNDn3nOry9ILdmBiKwopIDZsRP19WURJAVL7YvLEEl+T/DEsEQsY3
qbvhVcKxGCkvlciQ/DGvivChslNFPG9/H2kMbwjYZBDWGiCNw0DwHRvTrmweKd3J
XMHSPhBHbvR4uvcrk2DlkMFnkfkCyPS6UGNCc2qG4JRKwBe4SKQs0TROMh2lq/ee
1ux2K0PU7f1TtUvOReVtlSBLN2X2FcS9P238jGZk6TdmN84nHEUN6r2rnsG5OjkR
wclBm3H+2Ts6/FWkGkgXuJSreaGZeKi+PgCpgFu8eF1VnWgiNYeWXaZRIhM8oKZ8
qNOCfJnpipOTet0dXN3WgxvbeOVL9AOTFXa9mg2NyyJ86H8xF0nvFUyQULGVj1g0
knnBl3VLR2fB7WtDa9UICIHTk16kS+rmZ2hC5Xnavm06ZWfUWGWnR+0M/6FMYhHX
24W9nYgZI8mWlA38A0telHJ1FmAPijHKeA9ngQeAJdn6fdFvywNkdBFVvnVYkUPf
a74wYgAkNzwR9J92ClaIOfyinCnbCtgquWJ3oCLRVxHEEFcnoLi24lWbb9NM/wgB
jd8BtPV+lVgYWilyCcZtI4hsYWivTYeRqJOjU/vLXFmb9htBZbRWQ3wtAFiI1CmM
Ez50grUd1KCw4rcxc98Bofa6MwcDjMYvUy6iRROgdts/eNFGVwR+2ovpY/hj0QIj
3EV4rboje6/Uecm2QIXNa3H5UoNPkhdivj2/oy+eBBdG1RFpJiA0dgRoWdRy7E1p
amdj5G2N3HgxFNHWTe6BDUZHZYlcFo873yCuI2OINGM3DcIEzKYcuE79gW89eqHa
7v/UiGRZnDpLmGBnURd5iPYVx0Xoa6v1W3iJc0Ejvo4ysBEwujpCSLUHS5vDI85L
uV+Mpqc4/QND3jJfccu9PqpWufRwtsKCGrtxVQac3NggwoeHwB72IZJqEjrcOazA
/sralW6Q8f19/EXV8fbrpPBNVABbyZFRZ2r9w3GRl00m4eRIo1vD3HnpZ4MXTvUV
W9nLI6S0qEl1aZmcYKkLSyOYKZIeD8LZ7lydk9LQrpyDHrThT+GOkke1wCqMc5cf
nAujr77YIXRsS4JlVQjAalBQ6GT/8cBnw1krrMvs68mjOAYazQCuHJPX00HruLdm
1amM1bYfYPbVYn/+Rpaa76gwTbZ+O8WW5VxqkhfWCgdEkPvKoZcnIyQTrYOXE936
QXHTAfxjMXZjAPF3zqE0qLSz4sNpT62u+MvZ5Sbrg1ZMsFT6fl8wS3RBpNDP84hl
4gOBFbplGNWlJCjYyH35hfE3XHFfWm7LHAMf4gEWaW4tAhU/WOOcxwQMbBm2prqd
ltnvVM0ZbjjpVZlqMvS4D5jZy4GtS4nBp+zMxAzUFmvrvGv0BuWs9k4Ntj6tr6q0
RSWfDFSE1p3GhF4s/Y0J1ZL6jqUtwNy4MglaYd/R2HZKkEY0f8bRB8PheVneVE2T
bvyqjlwgSPgqQ8QHERpeMs3x/FTQDxFh8LQ6WjMorJcXT/UaxQawPwqDFS5I44Bq
GR+tWf8SyiJK2d7rGMJS4oaJGaK1COGWW5jAGrmYpIt57F1H/tHV4qWuJgRr8b4E
Y1AlVZWgv/Q3D+72z2mSaEqv8NKaqxjgOaJE9kq/5XxmvQSXkeuhYC22cHvthLlG
caGUnD1QhCiSzzpY30eVilT8PfJ5lZaL7/ihQJUaP3c45SX19PUrC93aqvz6mFuQ
PduRwUjnT9nGPYbit636kHKLjkqI4COCDdCNt0q0E58E65dCH8PYk1h31kj3wnx2
vU/tpHAOeNt0z2YEuy1cxU+iMEuh0+yuCxyOFUUh/rNLppTcslEtCtnfs5gjP/a9
TkswQ60Xzd9PQy6mKpMCWe3cPVw5HGivcsSqcz81iOAoSeXziBAzNhZdqpMqmz7I
KqJghPcQoXP94UCRA8amtZKz1KvfFppvHgvOM5ebTiJTcUbuPRZtZ3qi137IDiDi
/o3IGQT8UnAmgR3ABiDQ7ceQMzg5SEItnAoLHGWfS3efoVDj+s0dTRRtlkvQOFJi
AUyzOYY9YefRHsuL7AXVJnAW5IxSrK2x+8673sFaiaHGlfO/GMwUj8uQf5F6axKW
SkvyThC3bTzRLngfOJfbBHGdx+Lpv/xEwFsZRSolqkBt76adeXADscCnWWLE8vFX
Iq08DWLRwj788YY199eiNecP3Ruv28fXj6ltqG8ehT5yiEYZwigLfX+WIs5oHsPT
jInWjy8hQfdO6lFxtbFVCiO0zBrthRreTNRWglqmOHO0fWllf0JvQ+MBstXGUYyv
xGBYUi9PvSJoYrHFTIGy2HMgihPfTu8qDcBedRt7uVTgZKgPqSN6j2TIyCIADO03
K94+1fC9JHMCRD1YWrRfrAblnW3qMhIh0QKwBH1Gmxed2OkRgmq1eSXImXHrLY6/
BGsn2h9nhUmdg6lH+tyk0dUvV4YOaA39sU5jKJmLFOEOpj0aVLvlpWziiq2SoYGe
Qo41KVGu8/uMhxCc/q7V8DfKXFw2pPGVA3oL8vUsHREwRM851gUdLBEPcmHzw+B2
PoUqMpIJad/zD1SN3IH6hGelYdlznIaFJBztWrDrveOiCHbenx8br5oVQJv8zMdn
yhmbA5VlAa6DJa9Z4b4/f2xIt2mpjm/lsLY4fakRbRhBj8N+tnU4mJLEM2hbT7tX
x4SCCVvam+yMVZsKMDT9w59cd0dA4r9ONd5n3EkahzmB/oj5uAUs5xFptZ5V9vpk
kkoIJqxIJ6b7GWkj8gH4MLbmcLfhQ/5dsBtdgiyrM7dp03kywd0IBQjeq+pwXFhR
DkMzeVKqTcEPyLTBRc/MNY04M6qB/MbjrPqltN8CUVQO0+MfvG+cWzEQ8mp8tjK1
yT24fUWwgL/+1ADiNk/8jgg4keliLmrPH+5+kN5e6TexR2rpG+twl6HT7GlVsTiT
uSv1LpUHrbbxzay2kxpnJlhyLH7cq61edx12nkvcnEw5oym399A+DxNK3RjdLn6e
oFCEI4ocAn/kc9JsVLfjeLMHVplvuVODoGoOr5oUVITYfVGIUsZopZ8ym1wRs8kl
8VIiqzfJz/tjGE2I/0n7PHjuhdi1rrcfwdutn91OAAM25QAJTNKA96jYMfIs92uj
WjFu2VmhBdlrPg9m4L72F+DzuxZojGp0WEWDNWvF7zoONP86VJ7d0aThdUCESZoF
zJK+DeLnsG+X59dxHy3l49W83Ai3wbRsxu8iePNkXcAuKdwOR3Vf0zcBV4FqL7CK
pxAzVXsYtQDOptfbGwyjqZyKdOQog1c6Uzp6l0xPmEIcnZ5/LNzvRXQ339dyUYRG
eACrMBF4AJ5D3B8mffcKRSzucum2zfsZxgMRVzKGDLjk3EX8f6ofCsZi8KsvGyev
93v0PTGB5RSD3W2yGnHpOBayn7LQT79xAv/YbhsouETKg9ZjcukcXpXa9GHahOdy
290tKNAdc6d0ovfQfPz+swHlWa6ywyAeI5dHWHmH26E8jfE5dXl0acnLsflPvBqh
v4YcZpQ/nGmlJUKxPQkd0rg9681x26HKkY2TlsUp8NVwMgY/wGa/70I8Sr49Pc+R
PcJbA9a1rCNFDduBJMbDAtsObb5V/XrElA1/AwAVbacOUWwueTs5xlwycaZwsn6C
0N5S/wJfeex4M7KDCETlDhzsfNRBYsQVpS/epB73hE6S+20VyOMs5eVM9lV7+UEA
me40XzM3NbTGOb4X5C1tUInHQIhU7gn2zDvYsW9Bh99WBNmLPzdJFLLfSEGuSzbA
TSJpwqA25kMz9771rSP6V0UGaydSLXLAohh01Ykq3BB5Evw+CjwX9dM56qVQwqgl
SY6a+FYT1lqE6umC/CqjVB9eaNvW3Sf5kd2ub1idhlALFx9crvSAXw2z4sq6C8Hr
VRLcwEErGbSTITHGYHMCykAKTql6/n36PELGjvcm/TcC8USOqKTuOvJbMNcTpySF
p4GaAGGogXsZSaFG5KVUTuXalCMRymLpjejapgdMhK66a0kIiFGrg4O+gK6XfZfy
VFJV36Xc7Im/0m0nNQAYZ8OwmIHBYVqOyMWSagfhEQatXnKG9UiSWksZMacPZpN2
hMAmKkJ0o9t8lgqAJevIH1VDd8i1yJcd6NwseqxF9DMcGr2GbX8/Sk/8JYjfy0AR
M/KfTt4ZYX0d9MkmRJnWnd+dEsLx6s4cMlpYUfax5bAHyRqMnusOuBI2+onlqj6A
lZAc4riUaA3DNrRoBJbf2+YpVwT8PGLfW9HSkXSJeMwLUGcD4toGCJXU152rHYad
eSvPYMR+sLN+5H6KCCoGojv5ef6d/6412IhDcQBeYwvO6xcduhKquYqglQaesce5
BohuvWOnuaoaNxxfQn9P+cIjP7Jgzn1JnHbWJMnkZ9EWx+DRe6QPrgkwUUsShq98
eu5EzFkPszQtuO3nmnvLlaYh6ke5fWeeMVgeRquBIPlyDyFcjNc84Jub6JNe5x9k
tfOT+uGEu74AmOWhRW80/yfMyCbkRV9vdSz0dbZvVJ8YfWn+MSLLB/iftDABL10V
seVuDsIsj9VexP7Xvg7/2jo9alA5FsBP2YHZWfpHZDNN/WFwwFxu1YrO/gNTgIbx
+Hr4aDCg9ZZN4uIeRnu5PG+PslMfBeDnRzWNiQVNeFXbeQgs53UWlKEjKhxyl/Md
QkyVBjB1jSfHLhjtMYMV+jQl0SDYLD6ZySnL4H2ZhHFk14/hVKU3jHGoFJDJ1ccT
fLoZ0N/Dh8Dhwm40ffZH64Zqg+C6MIdgcLKbZMW6zk40XWxS2FE+qOwEjEBz+WYO
iacWzKg/8Ccbl17eSuWXszzZzX7W5GXe+LkRdE3n65tf05p27yPyr0Q9rAR9RH6j
xhVwXJkiD+2HTiIRm58zOlFQiOIh/yo8TL1ZifqMEbyP+mgaijtMgnPwbaRTrzHa
8r4A4hk5RqGXb9oNPVwIpheX7/lC2a0r1etkRSSDyC1khVXVul3kB2rvPfO3Kbt9
ndqh5+1GoTaYz8AMYXRDOp3aVyKdJwlCSbvt0XAZmgHK5FQ2++ZG7IR6NQbW356K
TFPBGXhlwz/kwLjnx9HIZHxIsbSrQo+wwXNbhlVKmoW9DAaeXpkwElLCZU2BUsPK
8M7EO8wRkjwPRYlhzKep5ylhOfSAy91NJ2xt6c9/J5xJE9nNJcOLZ480TsShq2MC
vTWnqbxhI1UYa/M1PXZSJusAinltHe+gxl7qibcHHquxCokcz8P0rYXPPbm3Q1HH
a6LMZPJ+MrEKyqvsOd1wX3klj3OGrn3+T0Z+ixbM35to+DPQM4OXfeimCMHnlVXN
+ySMuiCBdGBh1XNO5Jv29u8fLJaTlG+MtwesQN1c+Cc4RjZM2nCBWkqcym6pDcYn
ACY+AcScqlyfdcLyTSTwKW4hMqCrAdsjjB3EQ5G45oys7oCx4kTS08BsKmZmlKIV
icaggn4/PqnVwOf7RKou+GKPuTyXM5BHub0Yg0BpW7Y0FUphmskVjwtfZ5Q4Qamr
Fn8fdxcljXo8sDG0XLvza7nutSfhDAxOi+xN/O1N3hnG5nIuKx5aDZeSux/AzHhy
MjIAcBjz08SyxX1vjUS+LxMEhSPFe8ROts2E55e39BEoNVr7XCZ5ddu0DVWgf9zN
50fvmAWZNBN3crSc3FVvfAL1Mhz2pp8RZ7r72jdfP1aWDRWi4SusuA69zHyJ4fSx
xg2Sxf0MRVfpWr14GTA2l0UTaiQVzf0fbD79RVtguJE090XADk90VxGVWg0Fxx2w
nJ7LDtP+V9b7OquNPTMcUH+amOI9q4SvKAefUcZk1qpx/+uOoIqvPXOKH2LuZLf/
/VneKFef6Xm1r9UTyTyMx9sFBM/efQmElLVRX7jeAUyViBivYUUnH9IbvKXKAWCd
3NifnLrwNLbYDIIgDTD84642KXCDOQmM6TQlS7uv/l7VoPPjOI2EFyZCP+d43qsL
yt9AMlkXxecWpgPgtK/SwFH5ys85aUfZm5nUKJtgbm7T5B0VLGyZjYwxXGAWwWOR
fPrGN9y9vLYm6cQsCWVXFxqTyp1VfgOc+/1fGnljZLS2tkkaw5fwWIG3sM8OjSqa
KzckWptKKAYRjBEl+1jyhIBFZX6tv+d78ZonRQ/fjiIJPsnDsTlLDrn4GpctXbw7
+YQvJNa/SBEb1vt/WvdDeRefwIgEuYKg3kPPaQswDJXaUvuZ7KLHNBqHWSi3dEoZ
Y0yERlTH7WmTUK11FMSmJZt5uyw99AAK0J5dc3qwxfooZux39USh0Hug9r8fmhW9
dLnxFbHdQCMCN1268WezPyGUNzPx8IJ/1UEqWE2Z1XPXzqKqwevlgWMeE14UwELy
oLvTTCmiX+nMTA1QIkVgBUzD6y25NdmXcBNJuYLDsWUZ6TdXJRiBf1N14DXXPSUA
XuCMk+EP9Uc9LYUEpMfeKyOwxVcXYu6ZDxJa9lY52TWI/xnh9BC3QZORgTicIhcy
36yS8Pt1gdjMbNt8cl2Pl5owAeB4QH0GfjOEXklYrm4xcntf9jeX1op9vwxbdQX6
MDT9Mf6mxR9PgQ8DNZdXWGZuamaPTjefs+N0igVhQ2bn59FlhmJrKD0R1J6bnfxN
+Ik6/c73hmQxuErytho7v9nYGGq0VINoFogCUGXSU18e0TpQ7hRRId+a41fNcVvZ
quUF9uisP58iHa5qsuj7jIYOliE5zwz0HuXzyIu9E5Y96vpIAKrjmZ+uqRn+Lcu5
ivkkJOfPQ3e6pLek1JoJuah188LUSEEZKod75Gn91pWfxuf5fZf8keCtxy2Enxn+
DfPqVq+KCihks1n+H0DmzP6My7C2/ibOOr2Nbdoh2QqjKPO254LEvZ2tmENXT9xO
WSJuqVXQW3LUCwaWdXNf/E13jyOTI7RQwjHs7dNVLW4O76N0v4xjfDk03nhxqkbc
OCrZ5EDxz4Bdy/BiAgZy/dnJI+ezjktk9JcIxb1qo0PRZHX1GpGRgqNF3W1TMxz3
5t443mC89jgUEzKeXMqJ+hKfZ0brOiT/D26z42xeGYVFxRTJNC1ayxytCVHHXpO5
kWrRi3ESUARIQms4AfX8P0fA0KWb+3k4IxKaq/q5Jd2VrSPXQjYawvY1ZqAA4apG
PXLVFwLxWMFUBLCXevYTfqaO4RvpqTBnUsibpqUS4LvIJQfefbli0VMlIVdoXKKs
N5VErc+qNHEerF/TGosvSNrX4ep6h1119rH4q7zFJOaMWSqddbUFgpuu341Gx68m
dPKnr5TM52Uqs+oycso9il8AyR0segNfNzd6epNHcIe0NAVh4Tv7SYIEDpZ344xu
ohjF7SOF+Xa6Ci1sWNkVzFwgCi1stVcA57ztAILU+e2dPiPTAGjFWjPm5vq5gbCD
0jNY1zVGBLfWmzM+vGVtRtxwFS1+QPd5m6Q8butX0R+wjc7yVg26ytq1xDkBz12M
o6pa54YrlGM2kWjr7bh932io5PlZplOS8Fl7JIrmc0T3pT0wXW85hMnHi4W0VcMo
pSVDXbidk1rrAP2YE5FvEAludtBi+eehQ7jnKquzqux/xoLsXz62JcoidMMo8Zub
UlZhd7dFVMMBojrMBzJJknH70k+UmTCDtrxN6zN08eI4+qAsCvqSjQuuwh4YAxuy
PNyT7TUn/VcPuULD13ORUELdbtpcNoh9g6gV/1I/Vmd3AaVhZBtNRoXkYZjsH3+w
rpInnUW6xlLyPX+u92PK608frX4mRw/JyEuR/jKn537Du77QEJQSCvDbDmePr/oj
FpBcg6Sz/Uj+CfpUQV6bjyCLjt1ue59RazhhtTVKQkTqPXPDHNIbq/1v6BT2G8CT
CYhbc+0NbtA6m5Y7g9LvVbxrRi+r8A3KQq3gG4CU1b4kRPlYUmPpEq6eZECsOk/H
/3iAtuGg3DwIxhZ4J6hK56gSbHzMxTdRWHmJXn6DW2ibLGMrckPyKFwLehW8JEMe
BBEmfna8YfPtlfJwUlfSFlHuhpPXmRraANJj0mnxgsRXQQJDDYs+2Bs0LKaRLLi3
Er/110D03VkDw0uX15SQW6BfwiSW712eqJOud7pGASR+qSrPW2tsM5cOQ7hq49Zy
9RWzHbbRFxqp05El+npLyFRIx7tqIZT1gkxjIgtO5JCj4xAe0PJIJnyAOytDDUgA
sZ0K1NN5IHueu4zC1TIklB9EX91z77mNaH01xehZKfKBPYDvets8ZPofaZBBrosZ
loOuG5mfUwh/I/Hf0FVGdzawrIxYCI/cPcsX17FVUmiwVv6sSMboOvqseYBwKm9Q
7GyweXMeSFyzJOMj5qU9QktjuldnMJm4CUREYR4Sc6cz6x67v9VDGXvjb5DXjJ2K
l6HAVmSW4hW1rYL7B+ISbRIx1OdkhuGqX+b8P7wEpZfAjqx+RcmGOtIMN2AKvioD
Kq0lk2Q1T6QQbV3RcyVRAZxOwuM9+rj2LpwICcqXDM1PMVqBKhOC/u3RDajkZSWR
hCLKclPox5pUaZVUtuxyculXlIprNTWVX9VucAWjNaJd9bRgKFlg+vrgOhdG4wZx
wlqmYjAKEP42EX5UsqaCfCKjGeTsixTArbKj+Dfo/rP9XqARe06zCw4QfbogUbWC
EahGMrOL0abm0C5vAYgXOivRLGVs9QhYmE+Z9gE64fo2zrAIVAqH3KKOmWT0hm9c
p2xR2HCnwGWAZPD/0/50Fpiu9ed3Be9q6H2a1eKDsWjAOMnM8OWQwFM+r3q9Kf0T
23MCLPbEKUMwd6B9OcvdE7QR7/4z6lgYUoh1ndhX65HL1bx4jl2+RoWxjhuJyPdX
2DoJkRUoAGfB8kxWLcdNCmvtK14RzezLG2e8LJMO3tLvYJRURPd6RhfQ+Cnmvm0U
L35+QT0Dh8ZGcAsIs2lPAJw4VY0ytQcLVNYOeBPTSbnD3nVnaa1hrueIA/Q3Wuu/
LXA9F4bB/bJifGgOYtIZfEMRQ2qLo7hqMc8KuNJ+hEA61oi1j1swwCElJtSSTOZl
18nAO3aa87pwnyC2VVFC0t6s/ONHwDk6On/3WsZih2zbW425IfBVP+5Aj88ywhsU
jcCcj1GlcWAsQyLfQ9RorhT9mJbWKS0y6SeS1e+Th1ocnFl4XoeH41ezKwIONmii
7Dj14iyXRNB1tFDBe38OKcyliOjD8jRcnqwBd0CqV8N+hiXbWAUy2k+65hYicZgs
LxJLaB++DSYEBchpBd7rrmEa9UIt9DLJQ3lMeNppQoNMzQU1mtmI7mAuUDO87Zlh
bYZKeAFY5PbFSARhr9DaWXcVY7lCWWUU8zjfBEuOCPe7yOemOlJCSsoAW6PHkZ5s
5Z1sY0dg9bUsmtXeznyS1gp/KAwwsk1D2ITnK9g6MiSBc8KRJGls7n5apVem0LXb
ghGNgUuLWtRvshcjuvWYP+pLqJkDLrvBID9X1WuBhGFNVlzIqj7t2FXoqPbGUQJU
uDTROBUhJgMGvSJ2sBQWQJGN4bdITuAgK5bIHYXJAKLCAem4IXLzz8U0K+rjNoGW
uotrU1JdKzpPTDWL6lmv1sInjqJ3VMFmQceuDq65rDs7TvzzM0HzdelBI90gHYe8
hm++Ph+r79d8zTf0wbYr0wXNd5Ve4h7S4nzSyWLtDG5HFMpZ42MJ13Yu65alQeU7
cJyj3xne+KU8VNF70c4efX2NaIAFu1Rx3+lQF3/ubsPwc3dS5v4LdnKJaebuOdrB
Cl4QcXVWS/Lx6a13+hSMOQf16WbFicVWOR4ZNefXUsyllv9BUXhgIfA2KvizvMut
REkd6AqpZH1S8+Ob5fMJ4EuKin+v+wKai9jHQZVjmiTHtS82C//Wp/QbwjsUnMxp
K2iHVauMMUZZcC2fMlrSQxJ19e75yI+3H/qfaMT0uqrGfEw/UBnvbkQQ1EFLrzyZ
MCfwZlYsikuhysITrnQes8rXKWsy9mE7AhJvUeN5wrmmQXBOM6rleqniJJpwM6oX
x5Td/XPCeGz8o4fbEDJxWymgEgONzEcxS0m/+ER07030p6SjKuJfEj9Xwfpm7eCo
uOxiGQFhJL7v7VHfSxpLmIOW2yLymZ9/ns+sZE0h2hA1K06GpfiSmQSe0ARd+iIP
r62JBh5Dc2/qw5VdXIdRTCdZcBIydCxgCMJCr9IYFgUpV0Z1pnDI/orcYrLgdASg
gjWWL2oasyo7T48tM/vPo5Irtr4YCDr0lPpIXTPpQ9xNMZvcn3j7fPeIgpEeNSXC
M/kk55PU3RAOC9pJ1aOP+BJ/y7DReCZTPFrBryVk35cA5OSY/p4zpGl7d9RRgzUj
+Qj4lQEEXV/lJwQOWKe8g27om13RRl0eXCvjwP0RTZZEHHT1Bob6gw339/e3LVYS
AepBeLwiQxRp2id7PozyBCQRSlY13RBPvTjVHOYHByFud/YncT0rM5k6ixZ6jeqh
uUi4Bbz/FYn9LOnqilS1GMI9LdDsV+WdKVU/tMyamiJJ3RMG+lIVrwfpPo9aVtYd
Qq8cIiYgH9LXTp+jva5EUF2qsImqKWGfaQYhJDlSya8BAFo7FEoDQgryKQ5G7PZ4
0aPincorYzXnT7ll1WYjrXmg2if7TN2nT1ARuQRBcMGIyVVqZT3DRiiym3CsV9JZ
tFET0sLLY5YHYk8G2CkcSvo7JbaZ8Dodj7NpJ/y3VKr29BiMaMoM1AiHhfCxszRf
PQBvGCQLgfSKC/8URjuwMzYU3OguL8dOFdPCLLf/6bsa82f90TGwtcI3sfiy+AD6
fRrQVUN6PlFCdJ9IxjREBnjyE6Li0DyOE+/dZ8Fvs32+czgJcP8VlVkVscjSIJ6k
ZjkVw06gC94+ZjrGF6dY10QjvfUfKbY0bJfjabpJH4yFBkRwtAFRikx9UlOFM4Ey
RvcRdEREauvBsXUayLzTR3TxkLNpmAJ8ikwWhbLawhqKGBaqORHu0UXLCwDmSQMg
ae/GfOpJJXdKyqEErWDz4aFESfLwwSyQpmUQmeA6LS4cCl2nyoqYIobKFqPueolw
sGcI9jxr5VF0Ndx99xPQE5bci8xRvC/uf69MomJXGJDHobgRSTI50ZYSId+25D6y
dPh75C3acqRheSneJkq9F8xU3Ig5VGj7xHZN9JFBmEiPLR/RF/B9cJr++jSVnvtU
G3vjcntlHCp/1c6ktE6CZlvB/YGJwRpJzp/GvTiOTSjGk+L/jYfoJqiYruJJN96F
hCqrB/xL0qkH+5LBMJ5hUhvR8Pwlf8X2/ock9BxiE8+iqDY3WUC0HUMkugKbH9kJ
1pzPY+lohiIOuwoFmRtFNpdFFOawv2iH8xhui7PTzoPA1pyNYAH94fYisXShHoaZ
RJCNTIuJYVz7BBgoFPc8gArm0fx71pbvyzXyjE27pHv4MuVsEIPY0AHXum0hxKKo
ZCv4xQiNEkpYg720KeH3RMXpOe9NIc5i7EdiytcrCL0hTMiPlLrf4unZZRQQviGN
EH/f5HujCKOdQmtJrqaUn+0Rp8AXDF1bhL6j0t9uvxbhDC7f1uI/OlzAum02RDwq
y8JC5Pnc/N7hJQXogHwihOAxWZ3/jLCLpm1BCwUMtKhp7M/LuVXR/IjbPo9Wz1/k
lUuh2as5K2SDvIIV+hvsMFC1lpPgVWpFaIxfClmo5BAFk+tS31i6NQIG1K40Wh9J
A2mVZjr/yxJnaFEELCDzVQ16GAotSZV09nAUxweuDkBjhPM77uKH4oQy38wWURUE
69QfqCNZe6yYAa/fzZ/r+RC3mUSEHFP8/+JHrBSrq67qM/3PGSFA6YXiOOBOKKHM
yOQzzFIOpT/W3WkSD0OUbI2GbISNaEu/zvqnvDELeIBcM1Af14mRIvOMHw7/CbaK
x4Ersph/i62vSavGfvHfAnTQ2qXv97qACzpa2Kl35ffbB/3rQrLb1MSDvYlrqtPd
bwZ9WH0UFEpOGVKz9A1helQkxX0bYEFNTT7Ifmw67uD7zXV2zmIVixvBhKWhbH0Y
koA3OBEUJXJl5o0zT3M6/WUyjwA6+ZwPxuWC3h7iO00Dm0Qno4XCRWjhUTOuIB9d
AndYUJrrXAmaDCST9l78svTtcGhCU30+TBlUdcviVYVWdYJ8SdZehtjqqQ+ySt0u
y9kUw2UQj9H+85jb448iH7TIvH8aMOKJUt5+U14QGqeglMfF6FLOu7THTzFBL9/u
OgfJ3MJyIyj9G51KI5eow7Gk8+5W6pqQ3r7CFfEBNaKADp67bd2vdP5wJ9/oUQXf
QxGnE3j6TE8Ip/anXIKsvhfj1oE8uJQkhbpQsQfXpbZY6/mh5SY6Kerm9W2+9p2x
c+F0wtMs8RK8aJZ4deb16/BpV7lWygwXYWp+DokgOlyqVmx2r8ipfupWbgejxJSS
kVxhok+WPzfs0c6FbvpobVQsHcI8q3YdHiZt+KHIC+QpJQXa5kK4PLsK3tQ2N6j7
bQzbqNfqhh0rtTQVtjQKo5x/uD6+HpC+jSSod9YZThSfRhTtNRBIvsPTd5FhQm7l
E7LNI4S+N3zjbkG1ILSrtZ2n6cGaN2Jck4Qpi/3Ameg0rDQpLQdFlhyUWeOAzTvu
0/0la86FJyAQ+BQOt2uVp3ej5sROHjDKs03qCP3M0edPC8alZC8PWA40MSy4jwqb
074m3c6Btt/MtN118dH8B4Aptikl3nnKNKPnCJJ39uaYgiEIIF3W0vd9BonE2Bkt
NpB6bhLOhFcFKeazrxkhqKGEE6Ya/8Y7XlPMT80VfjtI+1wlzJfmJW7kw1xINOHj
yosWnKimmtx5+F6+UClL8sK3bAFcFBIDubn8z5lWIoIPtVwRpH79t++JrEIu2KhK
VoLLCl7WiVC1itSs5ZrWp5SQAIH7O6tSv+43izafk8ynA2a9ZvXd1UA81aAZcjj5
+HP7kDzY9jqqFTkAYgO9gT7ePoNIA2OzQK8bbwadbewSqr26YKhIxGA+B3BnkNwq
ZUPH0hwfcEnz9aDYi3SsG9T0O3M9NX3FsPWKdsAq3U0SMYIOPWo697PYBO2xb38L
cVJcqKd6lfgxblwB5aHEk63N2+TzaSqrm1KZ8QEEei0yRA25g/sh1ZYUpluH6CPM
ht6MfHybGe8pcXVi5T0BljcFf4NZ1b0k3+ps8tcedCqcz+O0WwccamZVgIsG7+wq
5bTh2wBQk2qP58pbLhBibvtiQ9GmVt7uCCVnfCJKVZDN4TqXvmMAAa69gVrouRdZ
2RH4w077/SUUQZDmbM2xw3i6f4dCqBeUalWt8D3z7O0Bdw3GZoC+tk4ts3DMI7b4
7RqyDKR/g9yw5ZbsvAmDhFfQ7FNaLEAJ3PyzTFIZV3hgDfYLbfFayul6bwjliWRS
fn3JwRZ7nCPwQPr4KptUWtf6TFqYVkmY1hmOP+HNfvfKUXdkM3zCmerJsRlhlI05
OkCkY5/u3Uy0ertX07/yHtenjqyYGKTBjBs3pGne9TaBmnZVdVAoLpYAWK1kAuqn
UFzboKikQoqll7ZXnBr2pijT/bREMLUFRsBxj0wQKPdOepMLCJnBu4O47OMTEThT
l6O7eo5aVqDoDqvOOpozdryTRgYQq0xeS+Y74X6d6t7u+8w0v0Zbvz92cPBeCRuX
WWdw1fkWbcYvnddYdw4xvsWqhPxmcwIlEj170rGLSVMOLhHByjNEEyCSF3YjU7Va
eqmbH+SvCvIxqIICaIKTM2E3VBZvw9nbgklBKaqHNg7j3icNxpU5sktqtbYC/3wE
jtCv8/xLT5rNQUlvNXTkD7/zwi06xHbhDKHcA/PRMeAnP4VMo/idqx3ThqYjz1aA
TTsc92P40AsufQIv56DRSUuFDkiLmWUxJE4kH1c82/6Ls90TCx1NKkX5MzeDQoY8
eqD/sFHA7JuhTEmEoHbts/1S1gniFIPvesVHAmcMxK+sYaKTu8+Yl2S3T8l928jJ
uGbQsgE0847n9JBCoFTUAwB6+UHJWt/XMoLb7CQWuTf2XOS8C15l1Mwjz8Z4eRjF
BLTsA+VFOsQimo0+B+jBcHIJ77wlkeUqrd0ILeD9jGB/Ng46TjiVGWwHgQmSXLBi
IQuIodsJVte4Rt1HLpDwzhHvOVVztccilLcpqfBV6wX6LuHZxmJ3ojkSd/09QYHH
xjIldMId7FG5NrJhpZed7uh1xNFTMW0u/DmSN/V8vwkYBb8597TVOIYVlGK6CWBw
2/uYM3ROi2Y9pEy/ZZ3bjvQ5p7mAGCqZdpmYihBY37PYD2T17eCMz1F5KaD3jGrv
hlBZ23kkTNjVZRVTf2oyohvEtds0HUVctVqNYo4q3u40G44QOueIGCO3Iy+qQn8i
i7iQaTCsfWEqZquTNMkZK4Qoybh8lTR/Yz6Xz4nbLiM6V1DLgdBt/jJFan0BkPjW
r5QASXIqwvPFMw93RkCoND095AS0QhMA9pbHdEbK91x44PyoNPnAftgZ8gzzki9q
Qn8BVGKUMb8dK2ODQRC433w4F66QRSCl0sGpPjhlL0nY7uNs0IWBeXiUBgMzA5Mo
T6HHoRP7xnB/MYT+QjRgzAACx3MbASZVZCvk9oqmWjG5HlkT7jNhgT0nPhng+l2q
zREo4oZH53yol2auyns7/GDwpVY43MbSANUlyLpkYY/lCcbZbpuZ0awHvTmuXNRc
hohPdMIQWQfDtp7CPZL17qb6jGk23VQZS9LMHLFhHFKSYW3V40YE+DRgOhXboO6V
4LY+qDfPjVT4YqF8/OPGTWEgnn9uyB5ZtxvfsSACob7wBKRQJrYE+RmN8YA49OKE
y2b194Tjn8YLztu6Wrhj3C43LpRscL3CuDBTGfwwu+ubTcUHO3zjzd+wcSqN9bHJ
6Bd/7fOdIDTaURQ6rAYdd8uySDWCW9Lv9JE47/l6KhOWgI4gjl4s01+K4iejP/0/
sPkpCyJJCx3HPdrA8hV2+8AmDRuskScdfKMcHCOS8Dw41Hg6hGLx3RomwH2rleYr
IpWOmxFnILXtnZeIlufEE1iQcF/n3vA78decdRLapsG9nuxXT8JY+YCfUUP2zaIX
dSLC0J7zdnIkX1ckhaf3G+YqdznZtcrrTFCd6RTzQkDOr1+L9A22Mk+90zz1kfxg
6hQ5ei2ZJ3JJBFlfN+qxMXZZacgIHXwR5+CcbgoCRhZUOs4R66vHctfENK9MQ0f/
bIhO7vOYHXzh1gTf+XtBuLQBXnRVHgMS0+4vgrQX7bwWDr/uIADU9bmpkZiggNa/
Tupu5oEYlw8lP1XhP6SleoP0ygo2eY834s7/pSdm0EVqW+uGqyDA0qNLpVqTtgb2
k5/dee6uh2tA0G9zEsBqLWIPxsJEUQbaRl8CgMGBtXPvynJjQ+WPs5G6fW1hqWzu
sDYgccvD+PEsym9cF+kO331xGG7ywFTbiqfZ//cMt0enxixZxAmRvQ0gy8/mGh2U
hm/9duYgH2AdfnRgV5mFzIRBgI0YCo1kLnxjcWfAqRkw5jdjIDb/80s5OHkVpbK+
/pAkOIrTNZJPKvjuV6aELGw/ysqJKHrfeuh54cU5McWSSHEA+xTVh+QAdgwGFGtD
OSfuABlKQhazW4LrY1+8OO3rlBrEQPTZhXLkFB+CJI5LchG3fM/W3LZel8Qajo6Q
kNVjPYbnCjmu5t02TSgNNj81yVJDqYn3YfjYNwqZsXyR4F1CYKQYZtOjkecqx9/h
VpMcwIH9ELWYbP4Aw95StD1CEPVxRmRN7QIgfRA29mJzCs1HHw7UYS9lM7sLbztO
t/NTGquLL6Qc2lwyeqXLkBUZ8bz0AYb8Pq7A+nddY9Xx26viZe2Gh0A/4YYsIWuE
YegWcn6e3GX0L391ccLdXk9Brsiyie3n2sTBP2l6Wl0uCZR9hJlKcvMil92jJBKF
bheviYvsFhd7RsS3EQCUFo725WCI69ZsHnrgmiKNXK1zvsAO0/86oVQ9LW18W2uq
qNgCg6Kkfl20aZGLqqwb+g8EpYsw7dKg18Pyr4bOYu0VYUEIVXjYmHGs7TMkm4JU
j4y2ZNz7i2bRGPEYj8aIgaa7phmBJegZMCW/UDCH2QeMscFdpS2pqp2egTidKYF7
0SsuZZ2UDWewiXQ1lYbqltAG5QT6he+ZppaF4v3F5NjzqRLa+dM9jr3gHDFXik/d
BILKXRvaoy3TLwR7f3rkiRXeshwG+MprN+w+faj0QbG+h6X9ZItR1xlu84/cRZGz
/f8znAZAttO6vqN3i11mp2ECy8WWlWm97sRsy2/MnE2wQinLKuwfr+SMfV9zx/1/
G5DUjzKnwFQis18hiGzeDyL/8094XObClxTOovwKFCOB51A49qDPPZbjgitOIV2d
NJB22i4dhsTqU3LIreADDfWC89VMGZVEx83YHd3W5p7a+047DLGBE9MIBXgjsM7O
Hj7LTpJ/a4arLrM0HdYGWwiDNK1m6Smz3CKpi8JQQik49QSmzH59zCPFgC7Me3qb
T1IxYvOndETcGFvd0D2OoQi9MHoRUY2BTIlyAQGDSt45jbDicCl5pzm7ZTKRt2o4
l1Ge3UAZ7R+XhgR8Rp8ArsSJgDxUGYTYCE36GEWYJyVkhb7biotemowxPldQIBmr
AijlRnW4wYoCGfJ+ky/oRNltYPrR7uzKXOX0joR8Djjfu2EGRDIkYQqYFCy6sSqD
iyqtJxDHFPJ0Dgac8oXX6jb3Ye8Qia5Pxx8yRnMBbxLhKoPnhriSFJhFMccPpUjv
CjlI59MIkxp4Sz/dyt/W4u1DVHgTXZZMGHmS57I7hVixiOAlyme14Ewjh7vv/9kf
tkqnt3byy4a2Fqoj5njAAMY1ULEabh1PqeBxDl3QIIZRdcn4hR0qGW8h+LICNuGL
NjscHmFmZBaVe0hS0Cg6rK63/dXqdf5SD1njuTHm8jz7qIK+2FV/q8YuH0M53vMB
9fxp0b5+7ESvd4XoI3L1ArYO4WwhEqxtIKFzJg1ocRo8IyVP42oWQ0X5dOFferOi
MTrLATd5eYp4sH6w4pbFl2c0QDNHaBt7n60e2LG5Lux+lZLsn/kp04WiDO2x2fG9
FYHnZXamj6wGxPmVSNWUX2/e5Pv3YVN8lTeHj6Pup1755HCquGnzuCQZlI0GJXF1
K+oAGmifWoCyLQZNhnlVIICvD0aYdcikaSFEp5sh6rMLBOMn8QYjT/Y3qgMyhovL
9HruZMOMIC3kb0xjbO8xIrgEKl90B0tGe+pBRP5i0l2gbIBbCDrR/tnuuCCsnaqY
61Bjc0OigC1wu0sPiY3rIHbAS3vouHEWhdQYrLNx5eh2g7u9fViSOPqNLKdYr0Pg
YaUyC/GmdBl7CQRd2gDalioCRRqxXnlAzNqahVgaiKFele512TIVx+joTrNaz2lk
4b5YIx83+k81Eumga4hx1bXmErfRiGwNHHpIKvwnUrMyHyZuzPfc8bd1PFVhRCLz
h6S2DSrVQrdC55we8+P8YPi/6ypln3xuJPskeUOuFWkC/hI2pyCypcNpcoeY6b3n
yrj+Yx3IDnI84LgX8G1240SFvnxSmWj5DIraNoptUPfqGN/gtaaXBS9+71VPfElk
0JEJ2u6BLQZKljTKpNrguhKa14jtEz/R0PUBJXTbFFNC0sN7h7CFaCV9pJkMtgfS
kuh6z5OK8kcOD/aUsVcI705daa0F6V3HlLCnm+qx11inf06vY4vJMU3X50uO67mo
AsOTOCYawpcP2hgucNQSkn0oOuKe8TD8WXzTJGeO1I0Qnnu1KdV3fyoKAI5DOM9K
NNP9dBE1HwgUpKEYqJtYE8xX3xdaRFnyz9gocURU/vU623KjDBxxuUMBooMWaw//
MWq3B7hXPcKoK0O3d6UMHZVeGDmzvBJKIloq03ebXQa8x85h4tzfyoTNGnmiJnHD
BwXqQFsubrDNlKIRei8SQVW4pBNa85d4yatNLiXZ4libijGAlQ6FWIpNR1+LEz5O
XgZJT/FI7/jiOWf6Mta3Q/Jx/g0ocEoVRrfg+kSJID1LR+KTIdfIEbHze5pkHM6V
1SgHWNulZFxb6Av8RxCF9H6mDm1oDy+a0Vf03GUD4YJkDh8XtM9+kfqThWobOr16
Y+81tTjD973mn9obIFm4nuIvan53OHU8K8PsVTPlmkA/lR/0HZpSRaLnnhm/9RtB
5EI8UttTT50RJERWZcdUiv76jWuDG863KGuCjCJhxJp9Wrc8V/oXH6zDqIfhnT02
cMzpvWDc2cEBjyUS+nyWcitE1Lblyt8ELN6a5VLEcHPinF4/dNXEgF3WxxOkMzLc
woKxnQ+SSd7bEWejrflWueKIKgfVYJVAML6TyvMTeRGME4kQ/aoYuOYdi8I82lFC
EZsih9oNqmcupj9ojrOAK1MwWUawhppuV62qPy4l6jfuXtMiYtiedr7IKdyszhja
BeZWypx5byL85Csaz94in1NYQn1Lbw5trtk7EbaBuRDzuRayNcbfiIV0BFdhybJG
wCY27DlvI7HQqc3uFgrqUBwqIMh8/iBaMDGixXa7W5CuIb5PfO/iBBIRzTDdgJvp
JxBdzs+8sJoqjbQrXqffq0SJIcOKdiKveutE6fcVlXKlmGUVYS0xDImYHm23facd
TEGPn5h/htp16pY91qCg4SWX0U4AnzR4oJOw7MevGXCu00guJSJQjbBwyjneUlWx
/whF9fw9DjhgH99fPltjl2UgKydhymLRfO2uCapLCYa1521FLwd4j/YOLwy1q+C4
ugcYqYJLasxJP3DZWENc+9uOYiwi4bt83h0NqFpcrMTBW7v3AZ0AZ1LBvC7VX/kE
gZDxIetmvGCZLNxajOpGzOG0f7/OkwEsgL/p8SaUi+bS7ltOeiylXE6HR3OkW0Lr
rj8tEc3OPbQKGrEJ7b6ydMXMHFLIb74pIguvTbrUdVuA6EtYeXpBVaAN95G5V+7j
5sOJXGAei2hP3dm1yhpQ7/Q0E1H+jj9KOJS1PDR2+YiB9KA0tbaYJjhuo0r60B1B
JqdyPvAyGCLNJCpgctpeUFXa04OwLi+RXBHQVr/BJS0HpYsPWDiTCJpKz1K5s5tf
NC6/r4okjE2k2U0LOGkloIaC8AqpcIoFgtEfceMpg2lNY3NKCwJIhbu3KNfs8O8y
sitzzjAhv8LJ/gwnDW1ehJtsY5ptZMdSlGcPv0u01xGpGtxDQy6gjtaSeKkS0tdd
teXVRevFpF0gnqbNJzoUKCHNHvyNB+Nz1quelSpMWP0AF2OHrqQDW9onB0X2O48r
YUBqKP9L68Ds3Ne4wo4tOg+yX9VUGuwZOU3ZRUtYHFax9ZoNJEQX8HsgWNIFJMhX
0okrIkunka6LsXkve9FjF1QIK0nOWYyuvAXhlensv2dJnVEuzL8ZXbXPRmBcWj1m
G85mO7fGTvOqCBeSRCTXy+/TJXnyjLri8G9KpFfnyDEJax2i1VP1gIEwiaT+xa4t
mwf0AsKgZCbIiBmXbqEbUbW1iBUhmyLayLoV35VpmkIzvrQgArvR6tdLvBdj5/Rs
6o6p27HgE9EbCxuzod91FI5FUj+1MwMdu9d8RO3ko7rKOWpo+bLNiS/cJpIekNhU
Bzrdhuyh4kISN63OzO1qzy0ELWlgHMJ5+/gIX0hfA9aQTSzTCavOYBVcJjl4LkfV
oJwrHbPET/IxpPUsnh9Amg50cKtbNf+AZgvW9ghva6E3tFbv2VVPqccQddqRA2IF
LsqD5IvB5ceDpcnlV6mD7mOW47CvJEkmYvgoudBpi7161/TEaMmmcFZ8YmUnrayC
quO7xShASlfooswe0/vSYXP2dWz6Hlwhrf22OGTeJFQcw4v6Jp0sPhnT6T4Zw/O7
qSHxhFKvsQU7EPMYbe3TDcwPf/R7WFAic/BTF+DXyW88LKMnmRzEWbKqXhR/IpJy
DwyC43J/TAkkzVsw0+JSMOgZpdlRwwGrIWBBVCNdI6J8BHLMMv2m8keub7gmoNdS
vaOyzekMYylGVNE2feepiPv+Z+BqMF4OJXVKN0Y831niLtSyRZu0DNhJQiwXWlow
jJNsCAwOk2KZbeCdYfIETuBruCjnZSUA9Fp8KNnr5tCYNgLg1lyllFaD8J5+DYY5
ZMTnni/QNMLLLNHpmgcsWquAESO3OOiO3t78ucpUu5Fbcw7fiJ8t8lec0sEXUHzL
/U+yCWG6nc/+O2LYpdSNLgEHTPJ+X2nGqI0o9ZPOdjx4XMjiQc/Ud3OWe3NWwnyC
M1KgD60+x0Ji6vp6FiSOSMaXOoAGvWVASs6YanvfqIwHDVkeY0GLNJlHj3R26mqF
Oc324HNcVc5JbfLiCXn0sehAbkCfAHXVvmrVE3q2kuWt4EFHcoDpKVKRtwZKYA9X
Wi4ggbZft5oq9REqt3pCMQzV0k2uJ0CQqpqQRX3V3210tGg3bYCBrYktJwAgIetm
gOfz+2KSwdDZD+I0YfDc7lLJx3px3POlEfTgIo/Se4TI2ejIsWl0/ae1RRBr31Hq
+/Yh2rFTF/kRmSCdud6UAtHgZWBi8nE6CXXlsEFeZH/e0on8XPwjIXVyHPKi0TTe
9IB6fFyFvsSC9FweCv0loE7MWsAkm3xfdHS4hf7CWZjitu41wEekUkwPp4tLdq9s
aghBN8yfxKWbEKTAnLgqJssZMcq2l4OLJHYs3VwK356/SywQTB+H+9r34cP9y04T
e83zrq4KHOUqsmhgpJzSQBx9rery9RV4yc3TFaqzUKLIxMHQlpj4RA5CMFqMPnf3
63HlLnL8nF/J5DsMVpxxxGQPAtYr1av9QwaWrYukyZVuTZztOwg1pygvawF4ibd1
CW6ox928uZ+lANKtYSOzbL8Ynw0edtdFQQp/Nf9r9A5MfINXJXSlQEg48bb/FqG2
nEkeEVBGHe6VvG9SV3tkBBQQLhfve9gvDTtuJYwix5ftMeALOvgONis1j3XY3dc2
BE37/UdIWNPlRwwheBdk6qgSMkCLI9FIE47YZzZCAHzBFev+6gWcNFu4yb/whtQB
NPEh/iNFWDrq26u+QWbeJApDZNxoZ0ml75y+XdDdN1ElnzcKAxs9LVpRng2tVqTi
Dd+YzR5/HVN2xDceZENeNrs2+UlRely3TC6rUNNcJ98GxMAJv3o89SMTFHOuKSej
qhN3v66a8vHLTWNnSULQ/lBMyRqo6LJ0m6/jfisAslduCCmfTTXBy0wluVSNw72W
pzJH2px58xJ2PMbEKkSVHmwXTLzQq4Uc9sS3euLAnIXOXHn3vy8tBlk6jzkAU5Y5
q08SY68AkpPh57LE/FGFQ2kwq3yB67WzNp0OLJVS4kyX5Iq2wL25W9D2kQUoEHWH
OlkpXGg3iWmbbiVdYN1E1OYkcV/o8N0Ee+niPEJ53Q2TPihpoYWOV3YMrT+y7LnD
DL5dm4uZGd8Tw/trSFWnzb213Dnu3iSbo3KS+jT4IlJOatVF1OX9E58Kd68mauhX
z0LOX7HBgh3m4j+nWltKayK/6BEsU5W8M9z2H8oP3y4pUhbPCbnf289WyO7kgrZ2
snDUxRiO66N8kUr/osfdaXFMx/vHojgpyrNhJfyFFvs1XHwqClV8n2d3LZEu0sGz
Vq5xhqb04oCTZ1D+vEWi6KAJuteNvArUlsZO0OI8E9CcDwuYSnn1YWRx7708s7pe
BnQrl5ntxmrUA2z+duUqaW/U/tnGWLTQ6RV4rn+5A09E2O4MphqPqPJrIG1fyQHJ
noJvr+m9LkspDdNYwdjD5prMu1tR79/Vs873GYh/KBEBQ+4VFztLZUl4wQ20c0cQ
an+OQE7ekrxOPteYAWcLtVlgD+Jd7/r9ccQgut2//Iro7OVWeBOLso4wUN/P11mz
Y+4HKgU8opKLXKFJ+JzD74bZKRiugTwKYM3m3xNfcGdUTozNk97UrIA4cStGRJWG
io3DC+4/RSHIcyRNdL6wjTwt0OhWCwWJZ7ySFo/Ti1NXrGAeX4YHTWN/okdRrcnc
/WQ+CROJzzTtebACHQJbKM1q4CzYst5Dk2Tu4Le9rN6JGHbAngQp7Cl2DNKLQ5iP
/7ybDA2gAPiWEqwKmW85l3Ftwa5YvRcpoTPVbCzYQsJQ6MFtCI0Z56nkbSsD1VCz
1EyZlanFwdMYKbV6q/6CNIQf6ORKMk/Osuot6JEUbfFYpOjhpMtXFL0izIph+l7F
Ixt47ojqGP04nG87hnuLnknW5RO3pFi+7B1sUSU8WHT5h1rFhRTBKWxz4I8Fy5Yy
/OWn1NusgqrIG0ypUBXusqa15tTzHMudxgV5vSjNppVTKJIZOrITUEPjwnRkI8cp
PwITdTYrdz8wAs2HkjReFK7JmO/xJWoBhDOFqO31i82sijjxO3CfbzI+BJae1ehg
K22dlpfLZb8jwi8w9+czzt9NZT2X2n6wCloR5VkDnhUGZuhxe/aFKlcJgTt1gVtH
OaWg045srB/Afm7z8IRvGBxiYI+CSvjAMziGWfSHsY+XpfMIUrQOG6m8jT1aSw7r
iuvCpZtXrLxk5yuGXFvLzxzpBdJ4S+AQLuk/1a9FsOz0nYlObn2rFmQHdUnvC9jg
dXXgsIfYOmyATQiH5UmsBsnGY1merfGuGXxZ4mpVle5OhxiPq+LWpnfUvM36GfnC
Xrz01kyMRxdT6P/Sol7hBnQrpCGTHo5LA7ybpcwFMOxN9o3bIuHriud2SQxeNSRu
B0Kmnnx3+sAmharnMJKhGCxy/quiSzh+s5iRrH6XQam+LJ1WDIOZBVXlhbA1ZFEE
80/Qo7LHLGDUhO+NTp4wyen/jwgXniAVTgWwUvKD8TJ8fcPpzESFeysjGz2IZdjH
nuuDGTdlROoZUE4p9HsVStUd+zErhzOam+T0qEetYqHflK5JtTjl/ddXivpVvk9o
oJdMZfkMKFgkpIIac0QL+5jfXiLlxHT7NI01yvMNX0Mv5Las/JWaI4FHrcuZ3/iJ
hkStq9ysxH4XgSe+ooJIHVp33wGu4sybbmC9mhUwNcWUnv4N4cvN3N8nll8Wntgy
eUmDUHbbN2wA4Jce5dgz/h3XrNJZgx0kZA5n2mdWfmL7+2srbhA2iAH47aN5ELiC
vM+gdBts5IbOPvcYH1O9WK/pYC6rcpIQU8MulpmjcUr9xkn2OOTqs6krBh2R9ZoO
oKrR3MxJ0p+gbQgCbJIRS+I4vO8eULD2bbdrTGsxtP75iqATQYg3ScttWMUvLtpX
zYYPW8aPuMW9VicRCh9ma/jdyfwoQl6nUuj/arZOdxJ5Q9HfpISlOZfn1Qr0BS+3
hO76jvs/spIyRBCrUnsHNwylDSkPPMWnijhhC8OV2LiTYQYkDBqvQYzAWfdtHrLt
E/YXHwkMuhh8bSga6+b0j7/N7/KCU3MaFIPFdEDgpaoibf99uEzTz7HUOObz0Vy5
z8KSrnr5Muvp1af/MZ8537CoqU2jPsOrwZ+/3ycESyzX3yLH4dL6VdWNUWW/Is8a
BJW/J/YSvhPqjd7Hmsufrx+rxBQh4h9+RY8DDuEnobRNEtY6YXZX+2j6hd8DeTpb
7LL0m/1Sa1smxWe3v4Y/6sQCpoKAMdpR3up1ds2y2p4K7PyVWuDnqKg0PBYr/hCx
ryBwqJ0gK+vDhQIkQFyrpTulMA+OWBB2siiEsXG+mqjZnucGxRtgOka+AAfovATh
xzRwoQ8vDeiCZjlLhk/hvLjb9h0bq2TAu9gT9CzSU/z6V/77gHp4txkXQboxX6LV
Ro90Y47O6vjpU37IbxYA2+lIfYPCDTyGHapViOC+PABH5hCOa7qF/hl5OIB3gq/i
iV50HwrPzpWGjQ0dpx8ssGrVyjG0NCmt7dQzc2kgcH2t7q6/V4/mSu+EpL7aXvj2
xHY2NgPrUGG8TC11xSDnZV/B3Sph4YekoNh3li3AOwxZtILvcmDvVvqgDtAmkObJ
iJq7e0FefWcTXjPsOVu+B6ZflpnSnU7KEBEkltACXLSGAVaHXCAy4yoM8JqbSHzj
CvcYGd1144pWEb7seDGwzrcD6XLc2I1L3T5cIw89zm8xcg1Ds2jzZHZfCpUGf0ab
xPDenN4ewGmGce1K4VGWA5atJuC6vXLblVRuflk61jFPej1ryaQOq/ynLH9a2hE5
41voFHkeZLLjBvmgTK51g+Q5joE0mcvxD4b+pr81P/JXmpTASEqszgZozTzhDmgo
9RHEKsbni+vtd/XyY6JmdULq4WkcoHP1yJRzES8aKFXf2yKKweusZAclFjyF+j/n
0/ecb0VeDe7DpwpIeRcaSbXOXXQFawIqPSYXPRmbxtfW+QYTmo2/KN7kd4Vms/Fj
dzRQhMhh0oWwfWwcOclwD48kf7qsFGWSzbvfKzX/v4sR7+6woMpy2XOcz7cGjZ+q
2J87BPFzfmaVTjsOUT/Jqf856d96KCcwJbKQassEgUSQ2LA7y62f477j1EfAwp6L
fmFFtlWQrXNb3ozu2cgDVsPR9CuhmyJjOS5IRb2Rj0dn5nT6PPiTd9spCH0TRg3m
xKCnYWJOv/wkVV7YPYkPg04CB6SoLMVd2B9UYqAECLnWJrbwOJTRpMg+nvFFOREV
POiOSw8fL35Cfuti+3hU/qWw65X2bKXhBlrRDslyXNZDU+nxJ5EqNcFY0s0AX1+2
zG4TNyrFU3B+QniSgTHrQKpUkv6LpUrOyPDomeOqBPoV/VyiKnT5lDkF93Qo+UCJ
p/+QQLH8dw5byQBR5wHZAWBOhcQJH9fkTxgWe2TZzRiN8gGsb+WM32fxQN5UpxJz
pMZcz/ahGHcLMlzsDwxn173Xu99gGbcR43r9mGOiA3cE1gbbZXKnmB7ZiiqEZyVU
HnQU1ljuaS49CPlf6bDSVX0nvp7kUt8sLoaba1OWOtzbrxFfwM0fQ5znjxsqsRv1
Fx07wWzr9HSQDtxQKQdvoCZa9HhHQLIrQH+gi4EhAeRZB+zkZGhFgGE6xLvphiI9
m/d8OrtSa73XYL20NVKqY3luyYfc0KlCzXOm5v92fZW9oZoykEopEzzu7UfDWwW5
vemvdX1MHpVqQojJBugEluSC+YMG3fPaf1lOuz8r0t8GzVPVP1GEKL+HzoTbEhtb
OV02Kp7pLi5zHJNap97vLYObtHk/HmbhUPYBEcn7w2ixdjJe8n9OEg1aVh723sJI
vWY05xYTDakbihmuykdEChjnQ6CNOhmcFAr/NFwBcQ/6L2wcmo0GzDxFA7m7qoFG
OrFPjkt/ECZ97pwXvEqhh+s2nq0A5/217ie8MkoBrnTq03BPDtyWI9yeP8MZVail
3JOtfZgxg7HxUY4y2ZBDA4AVddGNV5cbO5nqP29bVwhGMMKBScPgtcTlNHQZqZ/E
98lH1NsQ4l9a9IZinQxDQHbQzPxeYeadffkH61jvEIEpNl4TKoa7iP+9qKdE9TUs
eeFIETd9ynv5IT/hgfzHOx3knRl+s3cx6Y1UGOlQpKo8TOnZj1daSyHhk0zQGwlB
xyh2zjaBLNIhOyfQynyji84Cmoy4VH2+dD0rXaStFI0Qw3i44JYRdQbIB4+DIeWz
nUaPJKZp79MJjWcKulBpbe5PdJxLNISw43O3kvr6d16Jt4F8F+QE7tYTCehY4/jA
EqxwiWSQAoa69qPcj5cMvwQc3dgX1nlRWbh4JotNYtLXeYkQB2NEQi+pdFcNaD8p
S71PYxmik1Z2FXYeLAbw8FpaIv3qEr3eo5PCLCVlXtoDnpN8+c1Cnw9ABGaj7eoQ
rfowCXm7Pu+v1lwPKFPfZDTvxOGurAQclebhu2rVSuZH+7vQ6pgqAJUtTBwTAVou
g7rxSVd2agp2NEGNNqcOpuJNkfrF4MpcGmAl2v+zBBRzm5WIXuNJXGOFfX+b9tj6
8F0uW1vmmOaULTH9uePQBr0lBzYcMmvIB7p9aLJLr60+3j7Yn+O88oe3Fn6ARELR
8jNU5EZpaVv/aMw2861ULcGbn/sFo5OckglFYNq/o8JKlLS+0CDv7zhXhxYbiFE2
qVsu7jMlGPbB1YXUCfcmkv02uRJV024zCv/sW5OL/mUBna/8XXAtEMgPhrMgLA28
PbjsLcazuljVm3CFvoBclBSlDrGoOECA3ihUBo5Zr+t983HDPjQP3AkhyZI+8B4u
07u8bG4dWZnoG98C8jPsKgeZJeiZW6Kqb2ysaXjeGUAobHmupi4XsuURenDv7mCh
Yhf5Wd5Q8x+0x3n+GPBI6qOUyNOihIzAn5Nw4pceffEsFQe8ERHFed/C63RPgqHy
R8+1+CHnuRqaANCY96pQIcdXEIiLVEBtsQZmQQgmVC2DC6WFGo6224NmzgjF2PUI
OUzz4h/Z/LZlUgRYAPXMocYiTFup8WgafxRmZU1798jMDVqPI9fFRfNsY7/TSUVb
NOfTVDx6Nsabao8vrhty+XYDL04NY65Cu30ah5Bnwrs7fMRUGwQ0qsHFNXuWVBnJ
P+fkfYUBHkOyf+S6TPkrPtmXCwKlhQrz1B2mGdQBmOEcGjgMX/X2aIoJU/pSBcqP
Qt5ZDgEryxlZ3jr4B1BarfV0walso/PR5adDXViOGi+z9mUI1dOxuD3KcxJFc0B3
hcAxXW80kiS0+OsXLc+xB9npcSWp2qba36szjgjcMWJlVkOzE5VBHGByBM3RXZmh
twiYVeBpwGkF/2ekgWu/T3g+8skmmiNpvPZnGWiXSPXjcrf++fnpkJPNFJcDmPtE
/B655aoHWZJmDtXCMWFi2Oyrsiy3x9dpVdPMAgcTnxy8WjFK5pKlUzxPGyKU5K1P
mzmqEfuszLeQKB3FOr/Xx21g8QcmJb6JWQz+G6PJcVfDVoFi1fK7p9tQhyB9xhY+
0qkBqnh2NesLqxp0OMQKl8kj0HF4toezhwiHtFIXlbip7Rx41cOtAalchIxzMXN+
mKjAcRJCA/D4rr9R7aU2iGhaq+HMosnuEE3CvglUte/kMoSGtqoUaX485BLwKIV/
X3cBO3aka0f52FuC6js/kdYOfV6q2J1hWbvT2qHv9i6YDle2bV/W5JQ7EmILzivH
nLsKPvA5NbVgfGw9ECzJtLFeuWjxerOskhEVJ5oyDMZ41hjLFiTKW/ArtkNoO4m7
kF499MIJSHvxfmFvxEk4A13Z8x44ue1XxyRZlsLvamdJGvzNw+vJiIbAAoGa6b3E
toB36Ezu0JhCK9mKD5saxgF6ySH9SsTxZH9DldxZAyimXqqgPwUrOgZhTQcqAaov
LHLywt2BECQRl6AKm2oGWdhY7mEEKRmbWWl8cA13FC235CUJXqO5WVSGh6DMmj3N
PRwIMgpuT7dgmM6iNNjxqn5hUCEavR/DpfjbMiwdeg1uGnC70St2PVYBOae9ym2h
GfD1od0ZGdgZDfR5i0QIu9q+kMdvXq2E+y/qQuKeBtVvZu9Gd57oAnxaF2lSsiaV
Ygk5FnOucrztSjAMdkD/mh2BiFJcFBzJLZeLpm2kdgpBwqjZzN5XUgfdhLK0tgyo
2OLLXZ2FNd7tZSX81U4rls2IeMoPBw8FgV3z72hwPH5WZxNw2Zk+9I2LkvCuSlfT
1MNgOJt7vFehYSEFfCGnOvwPjca+EqKJEgLE2kCakZ16qrwmaAK64p9KnO+ynuOZ
uE4zV9aJvbinqLekl7oY1mEMDBp9mlose3ZHL0maT4a0BuNVrQZ5jq4nuRGYQZZK
Ly3eNCQlRkY3f5Cnk8Qtw6ifGnKi6FzzTigAW3d0TZumJ6gzXXkMBg/2hJ/n6OEd
0lnleCWdhMD9ZF/IZu7/GmvitaBLMRWCQ7tnKhz3fnZEGPtFs8YgmF/O9Vtn1v1p
UHAvcMBT0B/sn8dHnQOOmVKRp0wS2Br3/qEt6BzYLqYF5O8AN1hBF7jwEcB3cBr/
9uSKQryhOB5xBAo0r2rp7hA+IjmSJzqa6z/tOMCommwcngKXCiFfbe4PEmbS6k+B
srMZQ44MZW6slGvk1KnwCnf3v9MrIMW/3Um/LbmDHi4xF3h3a0bZiaY5C8AD+tNY
fxgr27FB07vxS0LVWmfKm7EzeHLDw9dJHS++CuBrPQ9JdgGbWH9djD7J6/+Q4t6y
H9Gj5xAmjOHq4mjXTStkBQadgmqBhY6XzwtF6dmw7hvq+QzmMQKyVT/z5lvPZxsa
bxaKV5ZtrCo5OA33FzyLbgquBAl5BvvJfLsVIIFOMzh+9yPW8Foy/F7sTKYIthOP
ZSTlve2elsyF0Iiq+7yTzbLKPZut0yT+WgZSQT8B1dSk4yQfG05Oml9gX0AShPvI
AWAHVXX++H1IoC0nhePuEEmkn71tYOALqLFVs1lgjFhJQPell7HLHuntpIABVW5m
jSycUpP2oxL3QgUCTSmjAscCNJYQFodXMx8+5ePTgnI/Eyxqz3H3YTs2rVBacNX+
5C9WqMnRV2XLctPqkBRyxSM0sMp0pgmLZqu6PXoAQZpm8dO5f4zhzJsZoFjhPYte
/0bYr9StnG6fFN3247bgmh6xXZF9kAgjRftrKi41YJQBcRqsJZH6c8wSSZkLau0a
8Cq3ySAedDFB/6H/Wn48lq5fDh54P6Vt3KPPC4GznGTnQrHCyIL1qt2cY4ubIalZ
hP/V27vrSC46Dmf54Q5NuQcPYb8TUNxhNf+Ab/svWB1+UydqqjPPi5fpv0wpe5oH
ti3ozuo+ivbuQLMRa7XBXcCgrVkmJ558AK5FfwhdMaeoZrUChB7j7OaYLejhaMT8
wPwy2n+3D0gmxhAob49NJJnaOQnf7uFlnk3i6e5WZ81RvzVv4Ryd+Ig0paeyIKrm
Nq2okBCK/aQkFDSIqZ0LSoKt+INgfC41DHCpup47ru6KwU/Id4PFjgRSN8TWsOvf
OwsJC5n7DTRAotkh7deVOkhpKCZe4XB+wCcN0I0iT70AHsY+q/uqErGKuH0aHl7S
waLht/+YKZSgN1UvY1GIyG8a40srJRn5Nm6zDFYDMJcl7etO6c1kf9aePLZqXrJy
s9pghCRBu9eNtqO13gT+v4yE07wxLVpyf/BuJGUH4EsvTL7fryC0vkw0RROBOiic
7cfND0WHvz5z+IIcnAe/oAGZiqe8cHEkXq4jSy2OKDo0L5iOWmhfkhuhwa+3P/FS
6gyAGPVM0x5w/EnPe570k0vkpZcUM8359azfybz246eWPMiIpOgp11mdb4iic/2I
1cAylsZ9WxWG9aUH8uDGe4DS5UhkHkcd8Az/ZzCSyiqyrVt/dQoZ6UL4X0SNp3yn
x9LwKTywPl13YHJpxRhXgOFLWetTy+R6+yEV9SQ1Bekeg5xYObgJqjevgCLoGoHW
npCzywrok2qwyoeVP/vpWhNtE+HL4vjlCx9U2hxb3zOcZgPV4WUsfkqqhTOFktUq
hZLWpZ033F+3yjUJ760+P5nzyUP6zVUpyof/NO0za5WyoAjEnzTWgtAyjaJOwniq
5g5QkXXwHcYLy3Ua8QRYlWbJQpI7uqrZChqlHaWGknhc+5nqLfdY5qUskDCQLAra
Sk9pEs6YrrtJMzidXXlW4J8RvPexGFZcdsn/DWW+Rk5OT5cpBv6AWAyQABzIc/nn
2JK2HdmZvFTIoP/aiYM2nCive5x2hG/oLS4tVC0q0drTi6QRFOm3dBGOlAtjBehL
skMl3U3nWo+9zMe2+ibtyya2eq4W7Vd6rJ73ZyrAAS9sKXdXOKqU2tbPFOcwZnr8
zrz/D18a0xhJ89R1J5jlmZYIDJSAD8pvocNZQgYGBK7LgWTixHSk+kWemZoADUrH
Q2V3vw14bN0R/bD/NdnTCOj5YNqtFjKHB+cbV57ff/GV5SFbLvSnyvlPjnt2wJz1
Y+6fW82KwTEqztMXk8XIGWcTGopMkeNRjh5wHmd9A0Df+QuD0au2ITXJHvEpqTqe
1KyKgTs7ARSnFCJ5fRZxMN8suEJUmTer3m9M+a9F0+/HabtQdyLIbvXCS/Xwf1px
r4ZSruQaa8kdILwx6PuJ0+sSa6gj4c932VlOaRFYequqhErjf9jssKXyRk933U7q
60H7+ayXM68fPwkjr90p2mNxbI0ml5UTLBDM+qxFc3I/y5KUhV1XdMQ+2vvfAFK5
2bLLkfNJRNgCGuzx1TCJ4tN6WeoIk/ZDeFM3y/jEogdHhFRU4Cd3V03u9ZR820Aj
9nGyb8Pxi1W+JDLCedvae73C8Rf41XrgJZBheI/AGV/OqOg9Oo2Gu2wjlXwUHObI
l5JeZFWGs6Fub/Z5QgxuSazYrfFq8hX6tQh/od8qoKr8SpaQuOZR7iBLsUHKquZT
gqLHovc4cAXBMOLEn7OgIOu6ya7N9oKcHtjxmTHehoLogMq+z+e5NM1L4Typ8hxm
I/B+kbrMjgYwrYPGyEoT/RdR1L5e/GrV0g7PwFfASrSw24FYBrhAh1a7j8NCdlWQ
DkknTi2tIZuRkpMKZ7yFgiyQHWsGMsGEufMYrBELdOP+XWjaw15Xi7RDd6Z6g6nS
IXCuLS0SG3LC5VsFYyliFWklg4j8AY5BN4sgYlZbYbBOcZKppGQU4VydH0cA6x6s
/rncftL99yCwhNeCsTCuJRBKHKUHxdBJ5X8z0IsCQ3qUX0nSGWJh+v/CmztoN8Mh
WcUxBmDXJvsh218AQj2OXuATQzFng2GLSzo3g544VSxcxDVQ59x0plfr91XDqaCQ
3aqJwIvsWDE+7yaC0Ktu977WdhzAwTXUvnb/f8psDGj7/XGO+04uaDaFV57OJvjv
b/jn/hL3uVvyVVFsqLubrcxSh2qCsrRBl6KNTmtoZnurho5FkWcw5gtXvIgXxe0n
hQ0f/PgsCjMm8nqK0Ly8TwqOY6Xl885ScHmVRrMsAECSMoTCRdIWppR8882TwW4z
ZuXV0KU5GwpRS/Ndm59xLHNRT5ljFT8VL3qJV6i3I3aPr0IFxozNaWs8yKblqznk
QZhWSj8JI4D+38NTlG1vMVvEwb9jWMTlcfmUul4My0X8eOehPBqE6ds15Q5LJzbp
8ECvpc4wKoR3JkYoYpoI/n2SVpJeWJk7zN4mU2IYcy45X64Y1cDyVlCskkDBcB2Y
eQX1s9AHIvn8Q58aBWtLXSlH3RE2g9X2INlHqjstZTRx6hYGFkr/wDzyR7dn8JjH
6LSJyH/vYfVJKqAQuf+vm1T2VN/1VL+KXApOaw8nNlv0Xqkvk8PnEA0bm3yAuwJ5
QWuvn+EQsLTkJld+qpL9F9p8SmuvnYUAcDVlP7pCoFq0L+HMZgjn6OqjCVTtG5+k
ciI26MvWODQj+TwUXJKdNSPG30d9DSRMrI9DMFypg3WBIjSaNZltqv4xOAO1QSwF
cRIoOEnVrt/Ve+DnwQcBc2nciMZoZyQP7u0gmYDauQNFvX/GlRwxnGBztOPb/btE
pBWGDb38bRbMacXHMff+vfsFsTuGxflY1VO/7wIIYTiA7rBgGT/3cR+dEYbAK+UU
w8qT6amgYb8VTwCmplPXxGwKeBbzlnOmNxhuwrZAILTzRdcg6LVq+9Vr1D+vrwOb
6BqOz4l9L5rfwRQ9zLSnG1ApD+JpGgzCHpmD9+2EoM0kXLz2mRdnbHuSxhPD881m
2jqSHqTFipqp0EzoQ3dTQ4tc6ioMDeXi1Ap+b0cpa2Tj1MD/uBXMeAYjOg6JjZyU
pRwcdF3ysgLj5cIVtq19jz1w+3bjJqvbAfWjIbPJ2SQdVhn31kfywm/61kyje4ia
xCIudzKgFal0CHPO8zavkYRZVKCcKmb7/kXl4w8D9xPWRRxdTZhOn3x02a+GIiPL
DVfy3RcnTxbRXlXdx/eYE0Ysbbsv4xyFfYo10zKoLs4h2utyTECS/L6VjIw4NiaJ
88UO+eqaojw64k+QeFPOhcTtcgy1I2/dYtWQb9VdZmDOFAGVLw6IXN4ojl0pGa0u
6iAZYAzJu7wXXLwV5qkODtk1WOIJUojdomroN7dDz2mpibrGLkd2yPqBjr4qwq1/
D4DPrmDdJZzgZwwHYP25xmD7XmkoQE90a569q5nGrB62mF5PdbKQqiTboPIFylP7
E68ZG1XZnUcLC4C5R9R2CtJegUxiF9XwG0SBwZG5uWyvbRp7rCzP09+bSvfMMeHR
5UXdChr75dXe8kUoAXMBb+EYLzbtC0xVmKAGPmRSij5SQP18s2JEKACU7jcjla1O
N8155PmGJ4IS/PXY4Q+tJp2NvGjDcDu9Es6yilDVdhf67A8rjocw/ZvooxCbn7u2
eAZgTfvhmD+tqQcuY9mCmDm26ipR9ee+yebmF7ZNIs1k3tJkg7YCGtuAY1mVIG8Q
g9BZ4tscx+tKZVLcowp8UyDlbNoiPU6yj/XfPRQmf2pWCxTtcbarl1fE2xsFs18y
L+gLxO5R216gI+oV0JOymI2hzKw9ou8byFeoGqxJ1zi/8t/pPxkfvxsd/U9d/HhW
GSRL/1Aw1Sn8tu1Zkh82NuOugJWITRd18yl/4EQrSH7bpxnBhGmpNd9vMY/EvSAi
87qUYN70K9YrKg6TtrLQtvu9Ww4SGjcFkA10Q2z2ZHEgLAkuODHvhpfo6pG4VIV1
AKtO+ltJXf9AX3L5cNKcb34ZhgBBNKyp+B+d93wyYgENuIyYb8i5rRF+vXclgIr0
jlTrde9SaOr9BF2qvEHJlWuHgNANfCEEWQWc37ieLshk5oQ2fAHWEf4q0ciy4XS0
pWyp+5M0nCHoauAwmuKlvZSxiBd8js3Tj8Uii/1HPJQuUSj0412vfxsfvmaVp79i
oWNIvKtdvkydWyoIUzwwMgtYFdrh4zjGzVUf+xX/ASSvCp3PXjdOxYwqDBS7qlXP
ZQwlh0gc+ztT9pJxO8696iowxjkmelzmxNzMYiYnIS3HPgttCVvliu9pZRSNQFBh
LudFR1Hp+OnsfQS/aeW14O8yncoyM+QZoorbZfNEFe3LdnPKgwSTcAQYfqxeyqvg
PlQVfGWH7ujQbdCzt+kqHkZujCAUm/ujj6mBpxFZ4biMrbh7gcWoOBwU16QDm9KA
ID8IgextBbcGVM4pUU4UCEgAztF6V9kv05rDyRpirqqnsPfWI/Z84DwwFtG3lg92
cS1N8NECPpaaFahiSCTYLq25rw6ia3VinBoZgpcC5nAtl4QYb/+BQ41tx/CuYnhv
Ma8/osIIGXbIvBfC4CQSjTD5ZcRZDcBzrEVmI3oWuzJhgBlNfkgkfhU0FkwLxSxt
Ebq117GRG5ip16ZMy3iEXCbsmlv1QatnyHzbd/0HP8ElAxHkFLtZ5tdJti7PhZtM
mSfyXLgL1CDS/OkhSOPuK3BzFQjF+E2iGB4fYyxmY34s5M2Q+EN/KSG8XSzQ4n2F
qCjimYo1z1vjg7u0XgKkTb7DJ9viHCJz8DyjKzcUprNYXz9RbmEBaINZ5fnFIjZT
G6oFfOMr8M/AqdoUW7Fy1HXJXwB0gIJnbKJsEe2ewHDC6k7X7GE50U1KAj2A1sgg
MaC7EZgbS/xtgUSD9E7WeLfypWHf45IXzogwHKOQnZnYPeZ3U3OEhtO4kgvJVnV2
6nUXcE+e4Ac7qvaUlWp6jf1JusE/Y9yf7GWknz8XK6CgvZ5VdR2gXBL4GVHQmqtl
I3ExtXGbWCIJxMIT8Z88052PinVTZjQFa5M3lbP/Y4+s5WuuQ84hvoCGoqexsI8K
bTCeIoAcosuf6UFIfPu0MMsJvSUggDhhnpgLgjvUxkOcoga/8QL1eVtjdSwvjYdr
nitiH08BwYjuhEhcZOktdSTmZa4pe5QAcVHGyehlAr0HwlVF301edCfzkDsR+Gd0
PC7ny6CUfpyKPWUintLaLzOJTzIvOxIvKrtDyaUJuvfu0SnDbXSNBeFTVg+jFIpv
/Lngu9DxFAGmoZG+2vuHbw67IBGExwBEM/lWQV0nNwY6oBPfTLC5wFnpf/YRiN3j
yEX7rgY/fPGAU/slFxF029EGOf07NgDcvJPom1qJ8+iEvLsIcoSznQBmGM1avMPj
DGZBmQiOoYY+a3OM1aSe5EHc8GD242rgW1R/JwmnrdrTf0c+smUWRWJb2dorGRv6
qfQrdc8WLpW5VmoioWpMv78Tv6CayCzurAyKbU5HAXSiRjVw/yH9RxzTJj3YMvOq
RVAqalL6yCCP7a+UmxxBbn16Jh9iXr4eXmwbqcv4ZbmydB39cP3Q8K8KHiyZSOqQ
XfLYq8SLAauMwXvjbb/EbUin1CSs25dlikmwcRUbKzNhH9QAUILuylaSfVIn+iqn
tx+sDIUHOvt1kdca92ifUw==
`pragma protect end_protected

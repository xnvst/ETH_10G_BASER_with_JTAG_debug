��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?�T�RH��϶��i���z��%2�8�L�f�j{�0��c&�x���(��we��ɩuD���b�#ׅ[n3&�ZQ	L*��Z�����h�m��xl5յ��7P�o�������AX�g��ttJ��L�@w����q��/�S�� {�@?�3d��+�7fs粤v,��`�}*�}F*�@0Ǉ#[P�5��đ'���Cj�ƈ��^ʶ�Q�)��n�k�����Y(^h?��j3��B�y�ِ��eU��|P1n������v�mWK� �p�m���5����o�):��'��w����f�ؓ�K���DY�|UO��;f'G��Oe��mu��J�B���Wh�>�n����f��,Q/��4	)�g #��a�c<-3+z|O6u,7մyG��Q�͎X�,�L�-�0(����*&�+�G�~�V���3sғ괬��Q>��l3!�H
D�o{��601�wD�hi��Y����	riP"�q`��!��ˋ�D��c��Z�(Qv��"�L�}��a�s�J4A(���D5���	8rMЉЍK�~ŝz���={��T�tz������
rTw�e�V��v����Ǘ�_e�=���V�wQ՟�4.�!��|�B�r�i�ց���������r�@��h�`��c�I���W����ZܙO��Z�{?���JHq���+!�@���E�Ӯ������Fx�qq͢/�}�!��N���'��q�j��_"��#��&�2v��%T��D�����; Z���i:z�X4L�����4~��Zw��t���]^ԣb˺w�}@FN*-\A[T��f����Qnb,���@��<�o���X4��,� _��_L�=�j�O�R �8�Q��v��	ީ�X�7�B4 ���\�5�Wa~���V��(l3VC�����U$kX���z��O��gS�� �i��G,�Mŋ��@���R���zu���������u� N������;�9cLwL�.Gg��X�-�H?���M��[SǇ��	d��֚A�WI���i�PN=[-�˓.�	�X�P�����bm�%u3��Iu#��텔�	s_�s��23u��+X�(ڿ�!Wf�M����鳘 ��)��y/N��y��paVb6�M^�Lul�[�\jI�s���/6���m�b\�j��}=�BTX�4r	բ�v��
��l�ۣTT���	NO�����lL��I��6��Ȍj�w-9��mL�5��P�l���$�y�C�n�4�x��Ɗ!�w�bU�\d���ia���V4 %�j���oĚ�dEm����C߯@�ߡ;��awk�O��X~�P+��9���do7��I'��&�(�ʎ=���^�n���;�k��[��3��fRB����^�n����� ��1���UԺȹm[Rg�6��t��|\^Vrc���T��s�W��Q	�� �Ș�4�ˍ�4�ˑ]V�DTN�7?0��NB�mu������t�B����%{7����;���r9>N�G_���(\�{�V��7�qr�I������q�r�ӝ>����h�d��'�%�se8Z���>O�~��nƽ;��������*'͛2s<ub�����׊M{~���rl~̰-"��9w�&*k���|J/M��ˢ��Lc�W'���$��/XTP�rv�(¥���S�����y�8���b-4.#��D�Q������7�l�9�
 ���3�m����t���"�`��cڙ��'p�z�N��J����c~�9��/�N��u���%���Bw8ׇ��"��Վ<{/�!�7=U �v��tD>�k�J�8��~������;�w���܀����jׇ%b�.�a���*��TN�·�H���-%���c�s4iVE� ��0��}gEe���B�*A�֘�Bl�)1��S�:�`]�j{	�`"/g�H��j�iʾ �܂N�f���ay {�����˩��r�/%AM�2�'����1����Q�7�,2�Y���p٧nĊ�$���o�l�By\���;�;K}R��l��F��ALyv�8������Q���#����m��e��r3���'.�UU����1 Z�D�U��ֵ�Oq8ZQK�pQ��s��\�ҝ����WX���v[�n��F4$��MxۨdJh�ޗ��6� *6Z���8`t���v�X$��̴9�7�7�8���=3�s
8Tq�\r�Li�H�� ti���yY����߷Td{�հ�&��-G��/�\B�
�>_Ls�C���4�aFb�6�u��}8�`�`l��=�#�61��OT�mnժ�3�K��|�U��ʹ�Y>O��P���!u^p˱i����h����t�LO�v����K҆c(�Iܘ��̭��QUB�1"��ԏd��u]F�OX#����:s-T>�<�Cut��[�B� EЇ~� S�G`\��h
���+��eG�kY�X]�kA?���sK(�/OW?'5��^���X�S�s
����R�յ�Y?�� rKS�k.v�^�}0�D�'�֡t�d�`6g���1-sW�zղ��nr�'�G2w��~�n�����Zdq��>��CR�QF釴�h{h�gl���Ms�F�|�|��ѩ/Ns̤p��x3��Ki����&�Y${S�&42��вa�.�J�Ճ��H��0ʩ��֎W]{��n��"Sb�k��uK���h��S�A�����-�H�.�?�C5��{3��v��T[�A@^0Њ��(Ս�ڻf�.�^��[|�|�g�-ա��ޟ
TŇ1+�Tj�)a���:QQ���n�S������${�x��Q��p�*b�*&T��* ���b�F�ݹ.l�	������c�DG_Z�,��Kr]���kcy����^��^�4�,�6j�nEnR�>�۞ژQfj�8��`4��x�lh=��`����:���נ��=RS��\")��K� %�NRaTC�|���R�����p��f���g<���m4�1m��o��gEgZ�=�.ˆΟ�`�WP@Yrp�b�[��eR�EӼ��=��pt��M>�U��o*aڗ��"�4 0��,�3>9*�*��J�Q4"�,��NW?TL_��J�F�`4�"Orf�1'�y)/�C	�=lg�D}�.�Cc��.l;(�,)4��(�Ӱ�)O<�ri$�R�mn'�$|��7���q ��S�l���c&��B���y��!�Km�*&������x�'_��
,m�����qT��х�$ɉ����L�����o�؆�}�T�����-X,B��J��)CN��ots�,��Ԗ�PжD�����?z2���_q+��xyu�^��hY����.��붊ZXj��R���x��ӒL;�o�>֝rr�UO�I#"�u�^��d
+V�u���-E'a�v������eP2%����!s����fH7K*��۫�?I2��씑= #������T�f�;P���9̓c�з����|���/�B �b�x����{&}��G���B*5-�a�ڮܦ;t$<�|�Ǻ��NQ�d�������c/���ծbx}o�Y�.��P�������sa���>61huG�%As�?��2X5+��A��tp�~C/ ���*K�:l�VH�+IӲ�_��{N\ӯ�?s���Ҟ̤�/�D���[��t+����̑`i~KB�R��'�ڍy��_mw�q ڸ݇��V;e�'#�8�~��Q'��z�r�@����1�fq�R������Dq�*�\�Gs6��Ѧ{�o����S:�i�fu��{�b�Yc����c?[Nq?Q�y(���;dE�œk��\n�ސ>����/�9�FӃ@uhRHP�#��[8�����u	_K 8�?7�%��-,=C�y�Z+*9byM� �=���,ӣ�lj��]~�.�����q
��u��эKց�"�E������en� 	ǰ@=T��r����4�pc�?!�W�HvcWgόF?.�§(��� W�*-t�%Ö�x/�ެɉ7�/��k�@5��l!������EV?ߨ\�y�t�{�wcl������ss�y�U E�2��m����\̃uQZ��>2N�7囵��G��n�iU�������5���"'V���$�܉�����H��Hf�n�G�݄
�����R�N5�Z��ls/�6�{k�a�5���OȘ&�������ّ�v�70������bYYw���0<鉗��dt�5��3���D��x��;!9�I�p>*����������s����!�\�o�X��c�5Cp�;W X�P/F�<-��\�t�v����q�w���~]F}+}���"�b�w׍w_���ܷ��E�����h�/�Ʉkn�'��#t���;=��(��tZ�����O���V�,_��M	~��4��������.��9�$���v��9J5��;�t���LP�=����[S Ф�"g�s���.�0j�P�^�^�8l��k,g����>�?�������P��>�C�Q ) ��E�gcW�3{�`�"䉴�TJ VB�!a�	(mD�Z�̘����z]�F�|�Q,-�44蒗P��K�LZOe���="s�SHpI��#�����}��W���F� `L�b�uMbK�	f�+�~���L`Z`�D\�J/^0b�|u��`K��r4�2�&�)�����#�`���!�����V�A�^S+G1;-9���of������sq�蛧�@݂�f���Yd�<wd���mMyX$�[J

��kTu���h<�6�����m���"GuFD��#D?w��l=�L�M�I�ï��߾r|�X�ӥ\�V��q��h6�z��t7�b�5`*~��\P���f��N�7w�N@�1��' |�`A4�?h��vc������$�!9f���gu�x +Bg��-a�̶X#�����ߟ���?�~���x7s�5��&�s�@bb�. ��7"y�5��K��"%�u?��+��cx��-�0�=d�5Z ��K�����������/��5��\$"�_���1I}���e�r\���r��5��!UC�
��_��[K��My��f��,��E=#w�W�s�E<����tľ��4k��.F����Ы7u���S�G��i������B�Z�C�&g8����v	.�l2qC�@��ye�Ç���z@f��<��s\�pwk�3�1��Oe�#��e~�^��-�j����VB��D�P5,���2wX=�9�d�����(�Iq�8F�	Iu����[i7�o�#��q�{unw�9�Q/�C:���R%���}�}	�_�ڿW���d�p�P�hbo:��^V��.\���e���w�y��v�EPUv�R\Q���^	��:��?D'Et�s��Ҟ��z$o�Ӡ�|k�e�Ki���*�����K�{ʑ�d��UM�����\~�O��^�mlP�'�������TF���8�ZV�D���> <#G�6����>��l *�걀u��
�|��ghY){z���/����X��.�޲(�:0s.�ͺ�{���SA�#c C��Բ�E4�-[�]�5%3�*��3�N^���b���L[��Ǽ����oM?��⎞��eL�~4r(�:�.�b����1J�@���6~�N���c��j�^%@��;�����-\"�8��{|Wt���eсԉ,+�_�Ț��x��O�hn�3���v�#��m< �I��>|��04g�zG"�܃c�"��O���@�?�K)^�AC���,���S�U-Z�EO55�q=���E�b�%��7�x x;�w���u��[%�)���O]i������}��
m ��Q�w8��QXx(��{��wY�陿�ڐ��?R�\u�\Y@V����b�5�9uՠ6c���eQ?3�t`��������53��&���C��&}������w���z�Gxk��>�]g,�eh1y����*�n@� �!��J�Ӥ���R�ձP-n�k���E��+�@���=TM�	���0#��~�
�
��	���A��Y,?+`~�e�ɴ�q��|��;J0l�'��X �m�/�6��n�n9��M�Wz��k>Qm.���5Ы�F�@�W��K}:_aXQ�{m��g��%8g4��^����H��D�n��X���|�i����b�7ʔB��L�J���f�b��Jc��I�J`ȣ!(\z~�T?����gƕE�?hg
��\��"�'� �[G�Z�%{d�P�������������4�?��jdr����{	�1j#c�qG�#����i����np�	�)�7 ��@��$���7��٦�����][Z��9�/��{X2���0/B``�N��F�����f�ʲ��1{���l����ͱ��W&`��:�-i�lo���m�K3�L�w��[��6��!@�Z?�lmX��S�;�����C�x��6 ��7��Z5n�����x�n��}���t��Q�n~�K�*���j��ty�P��e'�����H�5������BN�̭����6q~:0ʼ��q�ֽ�ٽ��)���=T�OȞ� ���<���ɪ��G�����3��,ZY��>�\
�o��;�(ʽ7m)�d�a�)�R�&���ӁG\ǁՐ���r��,xY�L����6��	�C����2��~�\y��@�&K9J��2��/�+f�~�p$�6
x�}���D6g��4�H�<,J0�� :6��%��o�	��2ܶ�_nB��h2ȩ�� x�a��1�H<LkXM��Ja� �#��M,��F�"�>�s�j�I˩/>&�u�Ð;��>;��˘�@��1�n��(oS#�J�6�n�\Q���3��&���<]L��T:�v\:��) �7?�;����B؅�YŦ��S���`�rS�������(��!�`��gϣ�JS����T�gu�^2�����δ��1}i|)(!���MI��f�Lкg� ��(�\�n'2ɽF(-�)�|�٣׬X��1rft�!��'�0���U4���R�Ŵ!Me_����^����LF����g�℄h)�OF$��.ϕV�LD�N
K�1l�k��A��m��`�	��uG�_���=��K����W��5Z���4J��U�1= ����C	�#�R_�ݴ�8#�����&�>������D&�|�(Kԭ����ն�U,'ݐ*6{�ٸ��ӥ}x5(���1���1���ʛITV�l�xa��T��P���J��-�A:;n�˭?^%����YV��N���������4�E�� ��@7����yW�1�ٮ�/9�R����N�=	�b��l���������R(�����/�n�^�аt�,�S\��H1s;[D~C��bl�B�Ax�Hw\nqr���mG�RN�|�)�k�`�K:��ZY��<�J%���B�$�+�yy�+ HVF��TyWdr�2�j�m� hQ�b �~�Δ1@�����TOlXMԜ����Q�Mb$�٣[���������:�s �W�INm26�kkJ/�uf����{zZ��:r¹�,|�n�+���!����*�@�Jn����_�~�h�7�ll�h�zm�j�ڔ��	��'����3��p�Gq��f{�\�o�hq����� �:쏶�5���Q�B/����o�ds��w6��HO�N)����/�RNS&�+��L���H���]z�N8���)kqg~5�N�$:�_�MB�Kr���u���v��AO�[x���K��m�e"S�b־T̘☼k8�K5���޸�?�Ǽ���\Q����[��fls�t=:C���y�� �3��LM�R���W(�j�mf߬�sc
��쪦d�5%�!m[� �����>�-���3�}
�$�?��,�vQ�����aW2��O~��"�秫��e&�%����E#�������9�1K+4��5U2Y��l����6����t��`�d��5�>�������X�v=�D��R���dgkT�@����|� p�e�ƺ�7� #{�����Y@������*`>Kr�8�-_�y�5/V�7I氳�,�����yx���s�LS�W����5�w�9�"�R�qg�}��y�	�7�9�ИHe�/%
�r���1&.�ú����u(�Ưn�eh��������~b�R��OӔx@�����0�?�Z
��d��6?��;��!u`��f7cf���=W��)���$�������9�r��0<����?" �c�)'o���*.Lt��a��_yD�;Dq��E���C���6�t�9�!�sR%�9�F$���1����5's�eg�p"ly��~N�E>�j� ��1S$M�0�!.���=���h���'�*���C;��e&7����_Q�z簏a8J�� �uB@��ZH��8���YR��1r��r�,sae�,§r��R�{��1�nJ ޢ�уJ<ó6�8�U_xtT���o�|(ޝut鱧!5/.徒J�JV&_̫Jm�WI�,z��
��|��걆�:D�WxZգ����V�����3о	d*�!l���S*�Q!C	4d��`M�WT��M�'����@&[b)]��p���#s��$�v-���`L��-��%�I��b�L�ڤ������4�hV��lW.v�P��g��v�?:��*y6L=`%E�����Z��=OC��>�)����ji6�vB.۶!|�&��B���3�+��!r��tvdU��@ʳ��wC+R�=�Q�æ�)�K�=���y�΋? �3S��$1����G�W�È�q*$ƬO�}{P&�c"�-�(���p��N�XN��z��5�cV�Z����ഝ]
��!K�u�O'9�5T�ܫ9�G��![黙��g��1fڐdI@�]�EL'fWo;����?u���hV��M�1ͅ�y&��o����\V6UX֕�d��p���Y'���xc��Q2U�������Vಝ��^B�;��b��|&e_,�|� �G�i}���Ԝv��p�ww<���ndv��p������q��y^J��!6�Uh�$���*�]��.Lϻ��=3��8���Y��?"���?XUlO�VP���-M�ׄ8qU�G���׽���:!F<�Gb�Μ�n��D��D%�f�ժ� �j��N8�4��2|OI^Lw�8��W	X ��`�����I����	�K���A�ӂ�jz`���u��T8&%��f
J�Y�+'��h� �� �"�0�u��6���|�]L¹*`-�Kt {w��*ܦ��,/N������30���`����_�z
������͏_��S��B�
	�����B�W�*8����Z&���o-�̎<A+��.vk_oɩ[
BیcN�m�_���1���^ɼs�����Y}�����c������k�%��x<��N���ԑ��S��N�gu7Kb�6���O�����S�8'�\_M�W@M����9�s.�Zhc�6�:�(u���+�D��Vw�{���[���nTe��7x�>���Ƌ���y��ጜ5d��꟫$
sw2��.ֳl_̏X��FФ��HB�#~Ϛ$I&�"#���������@BDW��n,���R���0!��c#�9n�U��3N��7���Xg�:Z��0X���7�x��6C��Yh�k�v�<�o�5����H�@�ߝ��QI���̤}����)�	��9��c�Ԋ�+ū�t�v�!xU�[��CVm� �ά��Χ��s�k��	ա'K��n��Hm��� 50�锜HG[�z(ME��#��v��ƃ��i�w��ѩu��GF���}v�!���
ݎ�,��,�ԙy�6�G"���'����E�����Pq'%���#�@���<�X�u������/�fd�IZx98�)֢)C�Mܪi�����4��s�[EvHx��cpRz��^����0�f#u�x�_�	tH�@d��sM�����c�T-��l��]FL"�0z$��U���]��N�C�M��Y��i��Q�����Z�8co����$P)Å�~�*6�EF�nwԙ� ����$��^abf���ڊ��^6ut�m�����9�Gnq�w#$��V��weޓ���l+�h�f�Ȁ�+�%&`���Ѱ���+W�p�����l�\�k�6��¿���d��Y����
2��T��
JO�9޺��ΓS�_n)���
�/p�;sj�Z�k�*f����&�~����{Z���Ȟ+RA�v鄊�Ve
Z�n�Ib��#6I��C������;��}{n�����k��Kʉ6"��<|z��W�N`����>}���)E;�PK	��"���:YT��(������VJ?`�M��ӎҡ <�Cͻ4�l���ZЌDy1+Fg�|���� \�ad׻ʺGT͗8$G�ͻ�����]zD-�&�#h*k��qlA���������D:����e�Hn�g�"�f���NH\ �f��PF8�Zu�&���.N^�nN?�I�7.@�Z%6���*?�r1�T�����h��k�����(���^�~� l����j�1m6��܉J�5,*B�,g[c��1�q��&w�.A��0NG
v��@[���p�ǝ)��Z}���%���7^X�>4)��t������箮jJQ@��O�^�A-��1*�D=�>�+C�&Ϭ؞��KE���a��s��e��0<}="�G ��%��rg�u�5q�-��}�H4�4��
�Aވ���"lv~���13o�hϚԟw��)��� Sc=���掅��`���LXla!��g.�-�Nóu���_QH�W-���P(B��W_�f��/�2̴��F��[�!��Z*;��#K��
�lxM7ǻ�Q���.��]��.ag�W�|��1H�p���ţ��E��'���½�Z�#4��,�M��<�i0��O�@O�����/�����D�C�|��	�#)�?�t���Ȃ�����[���bo��"P�;����[x��]������	���ߠgv�����!�ew'�O��6��;���|�������R��X����N��C��W��h�1���w����=�^Whe�#[s+-�N���5h���B�ݖ>IɆj]]T|�euH[�b++g��81|�7pJ׌lZ�����r�S���.<���WУB�/��t�DUɲ�E��Hٺ��f��D���lC��!�����*�*�K%��������=)�v �{�a�Ҏ�r�k�Z�����Q�T�J�>S�6єL���$�kkpxw��Ot���&tݾޭi�lk���%B#>�6
�I�|��ߐ���Fq=*����xU�Ej��6���ȍ����A�Q�]�Lx��{XK�����������w�u[+*F��s����&�R�V�8�ŋ���Z:�e�`���M	
��X�f+a�ߏ]'ܟ��0K>ɧe����gY�6k�A�Ů d�/I�^�}��4�Z�yG=��7(@����"ئ�IN)�"@��Æ�3�k�"�}E�ĕN�_X�rZ�g� H��݊�b�k��謙r��W�����z�~�P�g�[aȺ�m9v�^弒��Z���c[��qEPQ�Z�����d�C��{!p���])3�t�vOeq��V}����~���8�;�3���M�ڮx���xV���v+�'q��
���oB�@
�9x��J]�L�Q�XNcr�ѻ᥆�dA��=yo��q�ׂw4��LF��Aֳ��%ځ���V������HY0���Ŗ�ʮ&*�V�����ѵ��:V���D��g�h�IJ�L�ɦ��9�b�#-��܋T�q��Q)�����tv��o�G�f���Z���߲�}���mB|������l�s��Q�x��9y�k���wD8z��l��t��t�>�5�nc�	Œ'(�P-���5�L[�Flc�����dMw�9;Cp�GZ�aA�@�X��~���|!��4�M �vA�}���H��s&��c�u�>�[!͡��r��ž��fw�.>^�5�.�n9<WjA�[�"@vD���-^��D�п��.���g�I�Ľ���7s�p6��) F/JR���5����
�m��6�ӱ����.�/2�Sv��v�sp6}�'-�I1oa��:����l$�vWV�)��h]̪27C�2J�L�Vd�q��ݲ�S�z.x2�4�����[�&׷�J�����\�}���謣��z��p�!��Z+(�B!�&q[ņz���B�a��*���A?<[�S� ]`�K��X-����4Vf���q�V������KXb=�n&~9���)�]��էe%�"�+���B��s,Db-?���X��������9P�\,���YV���7��Jro�q�u�v��ȋH���*�r���pE�?�u�i���9S�.��$�A����QR�8[��[�sȑ,h�"��L���C��Щ��h��`4��,�Tٽ9��/�/�q/�1�H�H����3>�_e���� V����I���/�Ŝn7���ڸ��%�
�U�،&�Y�v&��_�����w*�.�fm��N�b:3R����\�X��p�e��Нeڲ��P�t�3?xë��0�	Z�,[8S��U%�R�����(������~����{&ёHS��v͎�h���������sf+�����Z<�L�����7����K����~��y�}�	��U6^�H��̇�,��9��3�O�Ż��*r�,ˡ*:�r_:l�i<�CXST1�'���S����_��$H��Pk$#~�zD��#���В���qQ�v�k����^cP�{8K�{�uU`�al�����M��\��r���Ϗ#��Q����i�u�u�b���N������'�Gk�O�#$�� ��������'���%�E����H�m`�{����0�Z�y��4@1X��Y�x`a,�b�H4nv�c�m���əc�w"Ð�*���%�&��JEOu���!�.}P���L�D$�ѥt�< �qo5KDZ�	�2��.����цg�*�ý�ht�Tn�)|������@�}���1œ�.w����/B�T�h�`�$M#O�b:���4/��ą9{��
��$z-P(�u"���c4����������tb��~�[�n߶Yn�V<��� �.�a�s1�Е9Su)I~�h����sو��d���HKƕ=�
��PnnQr���:�"j�ߗ�Zji&hV�����b�<4�l��`�)��O�&u&����17g��+�-�RG`+R�/��F���ơ�������ouxUN��
*�s�g�7l�c1_`�bV��j��߽	�R�#�-=z�
`ƦG!2(���j�>����`��}�S�󒲱��^P xIC�Mᕮvͬx@���֤����WV=Y\�~���8�9��JI�g`ү���ߐi�R�q�c�Ԛ���U;꽽�k:�.��:�H�3��Q����GO�����Z}�A]B�trȚ�m�<`D!���4!�#;��"��@�������Ϗ�Ft|Mc7	��k���Dfl�N0X��Us�\��"�)�<�a%w#���C&/�㬵�t�bpS�E���w�KM�Ś����j��Q�$�}��r벁�"P�8��Մ,L��E�mu��3�vVn�.	�� ;|�����n�����~�
�H�n���D����b����(I��(���<��/a�c"�%���B��7���1'��^φ���94�ADdT�I�;�4���16ݒjT�( \Y.�A���s]��t���;b�>qs_����(��)�:�9Y`6�Sa���ũ�6+*A|�E��1�nN��&)�q��#�#}J
~�u6E���\�@��E�1�>]�~��R�x�J��1'@���w	q`d��ʲ���K_�^U��1�1hð��|Mw��\W+�ěMh��$N��-w�UVyz�J3s�+���+�b==�1x��(�P�'��R�/J ^\�rf^*���؅�Y99��1T�@T�j��2D���̢'�=[��\�Y��S�|`9�94	&y$?�ED�T[K�4&n�:������rt�\�c@�ryZ�C��&�e���mct<2!D�4ЗX���C�Zq���I�L�A);����F~�Ơ1�����̕#l�SמK~���|N�����z�J�'��Bi�
'������ƃj��G�����Řs�����ThP����"\�R�}&��]�親�5[l`��	�� ��k�"���b�e!�p�� J�K�q�k��s���;�[� �[��B�6M_��[6���� SM�Q|	<�'�[^nh���e�v��Q����]*�5ȹ���b
dJ>P�����ە/���PAP���O��8�V�`��C���<�6�6vŋ���ku(z�����R�ۨ�(,x��&?[�r�_p�d���g�i�\�UY�,o����F	s�qE�6+�mg�%��$��V��u�L%I��u� �(]�7{��&c���w&e��U��wZ@�m�w���ۋ�B�\�F�/?+r]G�[\��lg?�E?p���䐯�p,]P�M�4���nI�S��Cb�����m��F�Y���rM�	�K��.��>eQx�B4���'�o}��u X��ׂ\�~�#��͋.����b��ߠ���!0$G�b���u�Չ�;F�ރ�7����"��q$CĜJR�����:�gUp��FVޛ�@x�*"�0q��~�8���B�ׂ�a�u+������ϕ������?����-��,x�!t��i'�*�7��5�7��G!%Zp;��^�6濝��瓏~y]�%N�K�r��J��2c��<�$�~C$�: ˉ��B�����4	[Z-\�抵���B-U2Æ4���]]a&��X��T>��N�C��Y��I�����Ye�0����u�i��[;Z{�&����.�	�O3����T�:�C.�j��D��y�un=23��;Ï�� �s�>�n��v�Ȕ�k�L�k�{����+�
ţouLַ�Lt�!UN-FOi8K���汞�P�!x[8v8�I��
��}1�&�]i��8�5.)SFϸ.�E |���+R"|��ʒ�Ϧ���4-	A	"��%�",�|HT�ن��C�qI�L��+���P���u~�,e`	�����iR�=���40fQ
Ba�!�@�&l>׃��d���
59�AY���+��?�P^��T��)W�w��Oԭ^'aF��p�ey�KWQ�t9܀p	�h޺��6.��l1Rӷ{"4{l˔=9⛖�����l%��KH���ldv|�3�[�)�[l����ě=�:�#�Fα~^���7�g-Su���h�6��n��X�s��Vo?��7X�bQ��1�6�['�dw�%9�6	�Ző��Wa�.��g_����X=D�t�τ�t^�@!	������&������=�24&��0�-*+�"7us�����P�*���O��	H0wn;������1�hT��3E5�: w@��G��w�|+��҇lD���^Zs�l�lD6�o��0�� &=��l�_�J�$!����.�b�?c��A���4!��ׁ���n�z�1���g���<N�7������6c'�0�8�����R.����-�r���V��W#���]ye�X�h�Ƶ��S�7��G԰M�T�%�x8�\���aF�bw ��Z:��W��y�m��b&^���&n+�&���nFa��K"�D�]�� �,�K.�Xj������t����+n�:n����B9���@)�pV<�����W5"�U��6���G#Cτ2~�V�_qPa�;uM�!�'��k�hL��c��^q�a�7u�fL�hB��y8a�Ąi�C:�V �5�f�_y@<e���O~ZH��g��]
��N���g ��=�ry��Y���kA��𸔵�>�b����c�ʝ�%Hz�@0�$+&݉>����0�1r�_=Yl ��v���9�n��D��Z�L�㢾�9�E���:���v?*��C��9��X�!������ �� }��V�T!`؜b�K�ȤJ4=gԣ���@ܓ�vr8�,��/)U�px��Hx���?�ie��>V��}c�x݊6�y��c����<7.{U�9�	8���<����T`����Rw�HQA�r���ۿ09��l6c��QT�K������;O-��ux�� �����{�O��K]�U���+��S1����Q:�EhcmGd�$&_�G'ףR�rfw.�d��wBV!�Yϱ��l��X�/�:�`H�Es�yd��x�K z���W�yn۰�� ��m�^�N����hO�!p-��������Ǭ%�r������ҘJ��d���LK��V�>�&��cF���jW�J��}��t=x:4lm>�3f�{�Fϊ�-�l�V��Pv!pS��19��p�=�Xq����I��/�X�~M 3�W�(� �t,��%}m.k�]��r�v+lh񈃙� .�7��N'�#�"�����d�wxv��-kP�ؙ]�W,�++�\����;�^�M�84��Qs on`/W*E���4�Ur�6HZ�]_�W-I�=Ca j3n�-)a��:Uc���v0�������0���ڝ|V�":˳�����G��k�	̷�2�Ӟ.�_C+)J�#�]�:�@��I1�G ht?*5/��3m.#b�9�TG@�hv��|8�!Ls�o�{W�^8e�^ qTZ��D� ۾�JN��fg�I��3�n��g�R�K�b�8�os5���"��q�a�>cw�'��L)[��:V�Xz�8 �������8�K"��XwK��Ѭ��.��͈��?���z9W6��q�ئ!o��n�bO��d]��kE%����5kM�>��Vt�e/�����E��w��E��t=��������:}FE帡gn �$ۊ��blW�� �F�@���Xa�d�7w8��������N'N˄Q����il׋LjN]cƸd��4����r7r���� Iߌ�T�[i)��;vN5��m�x���\#�%�� �<V��s	y�q|ۿ��9�(� 1۸����(�g�Μ��*�\���j���8Gぶ��ED4GE�'����D����lQ��� ���3/�Nlr����JD|�yK��=!�HNT��"Kp�V�=4�FזtF�b2�i�x�p�~	o�M��U@+-A�ÿ���
��˓>�#��{g�z����/\|}
�M�,+,�W�a�l�m���L�3H�G�6y�tY%Y�c0lw��*F�)P�Q"Yx���;��*T��zS�̗}v����l��1-R6nS�J�� �H;��ͪ�D��@�%���Ea��I)@���{=�O�j����?M~.s�&Z�8Z�t�3��0	<����9������^��+��1���!����]��bֿ�\rZ�X.c��@�P�Piy�S�}��Z�;D\#^g;��L�d`:h(���M@�l|�蓯ԗֆU��	_�/�r��*_ ��@�ֳ_M��4y�f�(�L<�;ٍ�p����ط�5���ă�|��;�n�#ÆW\��w�� #�^�W���������JIh����So�>�c�����ͪUj�H�6�U��j{̹��I��/�q�5S5�B�yƗʗ�n�!��kQ��o�DQ.˩��o���dm��Q���`�쏯��Q���R)��a�Y	V���jP����Z�a�d�>y��Q�����0�9��+��|~ULa��׉��,��.�|�C�ˈ���,�|��7����ɐ,�d��k��Qtձ��\[EC������������r��}NR���� ۉ��A��֪����Ia~�����Ü��W��� k�����0�PϣM޲?TJ@rq�P��&x�*8�;��2�LP�-f�?�ײ0����,V��O��#vN1�Yw�r���k�Q���g���|��S�Vg4.��nYݦ��C���`5����Zr:��e2���7�ɦz�=�mh:����F�'5���Xoe:�0<V�����T�v?x&��`�=<{*z�t2���;`=��b_�G�q(n2��g��J�"������I	�Z�8�M99�R���g�����W,�����g}���?�Z�jޗ�(��ZM~��0����%V�;mߗ!ğ�G�0Y��lRu8���^�\�QR���@����n_���yH��]�#}��fϠ&I����w>�3 ���>z�"Ө�}���bl˅���Z�&5*����mG���n�n����4�k�����:�w	��,eoi�_��ib4�}�8��&�m�)3�G��2����7��'�v�p�N�)67,�
A���1����X�� l���$������م�k	tUր��to���_zc�W��(܃�Y��}*%>h�f�	��tP�g�4��kU��]3+ק�i�_��&��^���Q��k^oI���]��:��~�J��K�!�Rsҕ1�8��2�U��ײ�6]0R�$Џl��"}� ��:f����`N"��Rc�^%/�bl�Mv��@�e�
9UC	�oÒBK0F�3"Z��@֩��br�������N�Q���9a*�j�������t���ƀ�K����A:?��a-hcѧI�˹��$S��[Si�ך�$��.��-/LC=�e� #��K̫���Ef���Z�4s��m@��r}EZ-��h]������*-�TC)�ٵH��7����&�
;��w�,[����0�/��s����uJ�e1��t�WБ~(j��4�)'z��\�A*�їĸ�z&�I��`pf���F����}�a�:�|��ԟ�����,��q�5L������]��z4�M{��́}�W#Ә��<�.$�l���D�a���s�����IA�����=��X?G��N��i�h�����/٢��ˈ_P�Ŝ��A¼���B8^w|BW�i��{1[�Á^�^�bA�݁	��٤,�����6ؒ9pt6y�o	7��(ڗ��1OO�K���C\��ҋ�Z(�t�5�-X��o}�M����1��Uyy颚��S��D����
ߨ�QI�V2~R�f�Q)��i!�[��D=͵��ԡ,��Q�b���s�� �J�+������}��?�����N&fۈ��(�S�>vy4�Pb����C�!5B3/��:�O!���b�+�"){�`�}�'���1��K�Rv Dƞa[��X�D�.������ a�N�O��+.����(���s��\�r��Bª`�T5�����J�]s��TM�Ts�*�JYa�e���V:��ͥ�5^�\0g�Q/{Q!�b������V�����6C�Gy|���q��d�Ѕ@F�	�3"���~�f��>���!>�m�������Ix���eo�����J����	��`*�t�]1/ǂ�3ԓ?ݚ�u�:#5�tQ�E���s���I�L��(OT7$��OGc1�<��^N��3k�p.~P���_�z�λ��m��{�45�t�VrU_��$zxuj��ҝ���l/������<s����Iޖ��͎��D�S̲|K<�p'�r�r���dzu
c�m�i�r_tq�Ŵ����|S�
��i��*f �Y�,e�Q�i�*V)6��v�O~��gtݔ&�A�/��O�j�AW���bn�w/�a]�ELDVW�(�2��F�#�s�[ӄ9}�vo��x�J���!{h�G�]�tJ{�7ߣ��qPāb���5ϊ�:���(���n A�j$�~n�X�d�gv*x� �w��@���k��?ߵ�R����+ak�u~O���-���1ۃ�TϝT�#�c۽}WAγ����X����nb�6�hlKQ�ǥm�@��Z��`{z'π�ܦ��kʼ�I�3n�h/u�ڥ���"!S�&u����!窷��4��m�-�?��q�K���Pܧb�Y]:��)z1�w�đ%'���f�f�ޛTc�K��&�{�ԣ]��d�"��y�~���2�`I����p��6}�t�K��o���L�N3����?��8ĕ�(� Z�q^r�f3{U��%{\Q�U�Jꆪ�������pPޣ�ʗ/�s�n/�EU�R���k
$��q��ݓ�f�0z��#���b71~ɍ�{�g���G��lW3J|�_|M�X�3�f�u��4a��w �5�PH�O�����FG!.�M�4�t�ʃ�0Ր0�0<�KO[\�sY�b�m�����������A�Pa��T�^ڝG�������wᡓ�Rȯ,J�5�����a:q�lB!�9�?3�~��m%�8m�w&��v��X��K�X�a���\���&
t�K�a|޼n�R��EZ�d9��W96`2���5Q�iV  d
����uD���s�=�ܻ��4��q��l�.G�cJ��/�،�[ߒcDr�M��NRU�3�g��C�r�4Z��s������o���9��m�'����},UZ�����Z}�}��_���0��9�j�}7�A�T��=7rS�=h��%�}'M<��S��}�jQ>�vM���7���� ���R�G�T�މC3�q��ZXu�&��b�� �U����*�J�!��p�hRM�����e�|���$�X���O�(�}G�x@� w �s=͍IV�(�ol{��:������6m+H"g����q�?)��?��V)�4$oq��������Ӹ���-&;�Θh�p�ڞ�[e�HQU�Qb��qՇ��7�7���+�O����PT�B��+2���܇���ygN�A����z���%�"I#�#O8g�_�^�~@r�>\�N���V���Ve~4n?Y��S�'�O��Q��a�s�D�!��?_�� ��ѵ�½/a�-�;6�n��~E�;th!��0��������~m�x���n;ȥ�)��M�G��-u�σ�O<ۘJ�3�N���ɵ�W��A��������%nG#%g��3o�5f\AA�rG��l65d?5e�\D¢�'3Ȅņ�(���AS���=�;��4��6�F�I���2*��&�{u�׻b �֫
���34��l"�D_[[��9��{�{גy�D��YM�t'�B��U�Ey�< ���d�ԃ��I=-�G�z��(�5�Qrq��� �����7�`�`�3��-�ێ �o�"�a�a=.a�ck�r�ILEEڮ�5#+9	��<d���,4�J�za�o�/ӄ���g��f� =A��Y��q�0-V!���B���nc����	fKv:�}��D���g t(^�L�xjWG)����x���9���Z>'(e��4˗�`<'�n_Y�����_Q��P���M�����k����/�w�Tk�}�(hM�?R�6t_>�s�.�sD:7|�������&T��ԶTvZ&�B��E���S�)m/��g�t��w} �ӿI�ϱ/{f�&��$C��\m���,��h�e�������"���v�p��$:���t�P��;��dY�{��M�㭀���0Ǫ(xd(7�&��پ$&�� �
�N�d<�*�)%\N��6��"o��_���[F�j��y��"��<ۃ�+כ�\�c��ٿ��5�CR���-^<5Im����i�▣�Ĳ(�
�ަ(�N[���y`߾4�]e�S3~l/��lp�z1H�B����ϱ�d��:��drq��(�C��5�{R�)�L*�!��R4+��SJ�G�>��Ҭ��=�� �/	&o�=�J�ʅ^	qxgL��\`�˽�	8�k�h��iPaKoI�r��@�`���Ń޷g����)���=��Ke��jk���N��>����Atױպ._Bcw-�Q��q��h���F>L���3T��@?u7��9�Z��Ѡ,cS6vօ�;����Y}7�4T��f�Z�!/�"ڏ��D��*n�[¿ƻ���AL�?߲h�ޠ;C�xXd�"��ߖr@��Ѹ�M�������!˙�Q���N�G[�i|� .�]^���$m�!H+��-��^����M�x�O��ǚ�	��!ԭ��Z��̈�Z�V?U/�iQGEJt�f�HR�T�S�q�SikA	-�W~?ݑ��x�ѥ�O�S��/����uZ]��FUM�F|t����y�x�i�(�0�,��(;���y]�S�E�n��G���]A�u��ڵc��Ʃu H+xΚ��|N�q�E#��>��;1�Wz����j�w�&���}g����i2�%�k�<�1V��&S��ج��Ӆ"�;��?�!�~��0��ђ�5x�v9�=?"�9�$��zn����K�[
(!��vH�
���tP�Yb���I���rL��s>'ĩyL�eY�PM(�*bDx1Ϟ��O��T����ݍ�i��h�@W~)�˵#|J��<�9� 	&pV4���(�A��ۦ�+��w�ώ��%��&��wa{�g��=(��g���dԙ.�r�.3Ksb�����KD*6�'��==�7`az�9�i4f�o�L��sڪ�	�I�8c�Sr�e)�E� 6&�2��7Q���)��M�&�Y?�7�l�
��5�s?ً�����ڕ��!}~�D�T��Y݇� N��j�[ �u�W�u��x�i��zYKt��P%���ɶ�I�͞�a��0���3����mw^C��bAP�;Ǣm�
�a�M5��׎����j���l�J�U`��g��8zj�6c׾p��t�L@�?y�^8A<u���L%����[vY��Ъ��-�sŋ%_����&9���fg��c�����uԂ;�<5x�YĂ�6R�Y����������ly�q[���Z��!��A�~��3h�Ir��Ak�<�N�W-߿�"^�!l�'r*�ej�blY�}40q(����X!����.?���cG^�:7���Q���28u#���p�#�\���C��zm���S�$��X��$�t�FK~L�o�S��K<�m;Z����r�(s�׃MCd�ѡ�V[P��'USE�dO���Ύr���o��,�{�|Ȏ9>�o��q^�x( ���}�yk�+o�P@s��:ؗ�?�bL��k����D˴��@�j �c����&�'������6G6���l�Y���*��p�k�ӂ�����&)�A@)U���v�s�w>���P+�D�7���DL��0/���Te"%�7ˈc��: 6L�dzq�� >^Z|Q~H`3K��p`b��b.��~jUg���Y���J	�[���Z�%$�-L���M�cu�~���ѮI�����(�۟� ƹf��,�i"�	�M, �*�Q�$�!�qJ�8��c3����to����-���:�0e0���7�sm4XFYJXI��ĊXl�=#�^�^ǽ�9L����2��`���ӑr���m�z}���E�D�Z!٪�؊#A��lb�S^ x��Ю�е9={�X0wV�H�1#3����,qyq��k)j���D	��b߲�b]������'�a~N1%���9IH ������in'�͝���u˂�؋k���7�?�|~R&E[��d��E�|l;�`Y�*Q5u!��~=�fr9���"('!�z+%���/�ޝ����U���F���8B����b��=<f��g|�Ia�k�9���k��xh���_H�s������f ���Y^�%�3�2"D"��cX�^���4¡(a���tI~�7�yv9����eD�������3E����qf�Ҧ(-��;��\���[/SE��i�ܫKK�� ^.���h0��D�n��[Ui���(��#��.��G���T.��/��m�A�tO�[�7�2K�3f_=M�;�H�i7I�L�
ԩCk�%
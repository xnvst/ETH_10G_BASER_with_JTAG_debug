// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
AoZyOc2ZPuAxDdrW874PjQ0mGKJgGbV5X/pQtISR4anWQVNNuQM472G4omdtXvyZ3OnpTorNQ2kx
utOVe4V8EVF0LT3gdU2zXAkrWaebBshWt/x3eZNhfOz2zHD7R5na6NwpcZ+UUj2wcrbjeiq522M7
xvTNDPysyxUGQABdjxCrxTaxy6jYE53oEq43w0KEN8z9B4vB2z36BchNOIbC3Osbf91GiKE+ubg3
wI4SHuwynovl7o0L/3ge9QUfRFN8pe2cXcydfHc7CPHHDdeJU4J8UR3DSwJNCKOCvHrew9KzKqJ/
30uoxsHHwWBSry5tPJpXAaHaYdb5wxELMrORxQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
bRYUZhEdg1DrDpyOqWEmKZuZIUSxw8yEVQ/jf8cT6uFncQQBHiw9xuv134HPl/V2PwR3Hemp9bv/
Xauaiw++4xl2nBgnPMWucbWxgV1rqoBdt7hilCAdifMP6spuLqPYMQba2dV4UqIvM5RYWA2wl5ov
fdB+MKgi2JL4StM52IrLqDynItF+MPUWX/frWbgt621cfPb7MjNZJNi3OoOIkDuqWYGmwr7hxxci
BXRShoFACgrxM7h2tt/Le1P/exK/3TGFyr42wD+5PWJRmweP3PoSc2DfekdvsMR8MzC2rqwnvFf5
kzZb6y+4vWf03uncAjJMVtXTAabI84rFnZZlaFIRe7Ak2UvZG1naJRqKBncLFtfBLPTOuvOgi/HG
mgulAClMqEKE4fTUtxov3IbnHxEsOurzPOu+4HGyLcjiH9es50Sc73uTNZxGrhWmP3c3p66YB5AL
XYs6fIMbURQEgq/Q+ex3shB7Qk47seAgAjMrzSYsLJhoHcmshgLtjp+M7OOTeSEjqwJza5buXKZp
zbjnw5jq1nQaYa/w4H3nauyqq3t3lKZFul1GMnt/PTmPxUQJfXrYvyz5dnwqR44YB/1reQUchDlc
E5oKkB1+VT3JQE7GYzWZR8MJPD7baYotyblkm605H6PjJd4n6tMGZOqwjdkKn1g0vfaYN4R5cG5/
XlU0JeF3+xmHjurd9UUTzNxz+hK964dnGoPz+xCykcO8PdsgOO8Vx2sPTQqxmsCLVVBKQ914oFCP
DZkz8I1tVJlSHGCsaEe0BQQaEMa/s2qPQbfnKNxsww8VBjFf17FxdSHA09UiQ1YLn1H9cBpDAAuN
/ifx5bUwvCkn4c0MKXaq6YW7YdmwN1gJeylQ3CTn9ZDlbpHPFl41rtcofPrE7UwP6PMuqZTTqefS
bn09uxz/pN3dLfMjfpK6kz8/TvVzsHrrFYKNPyXrZ7SieEK4C2vSXA/I7S1Gh+gs0+3HBfBPMpZw
LeuCdR+PjBRG2JNNRJSKOBUXQSB+ofWm/6jaNC0LGl4wSkZvCSuaOGUfxqTr+HqkA2OA2rYfU7u0
ikc4UTSnzerwZU02/4MECRA+97AO2DPPbc08PWpxoL/m8K0LBP4FuMYSQksJXw0LTCv5I0bjVbuB
yvf2i+6GHxKnoweZOgBCRgsmTVvGjNClGvCaqXYUF2EKVeikdyIusEcUkmxvkfJCqj1UDKqJRjrv
t92Bt1yrkeY2hmjcaxeEsSydU467/BheLqv8wuBI0ZVnfwk9fU+gYEpNB3FSCwjoQCTCFM5itv0m
5hhqs5AoltbJ/kRF0rZiqYoJ5bOzGTTeNNwe+XBEunBnrVwqxH32GxFhBw+sliDWa15UG5KXZV2Z
uxADiVY65wgOvs8MOm5BsVe+EhiDqx3BoY7cryz1p02V/u282klDA1XoPskHqh/NzWDtwU2s+a0M
A2gHRqHEMm3Rm5JjBhEd9zcmmVOWiWxH1rW2t0cdG9eA+lpgkZAFo+n7ci6kQtzBlLxcpYPctwHc
6rj4YrZPdEctvA6LQZfg/J9AwgPwwIiiIJVIUNsPVXeQQWqoVUztXReanb0hslH8KO8A7iSWT1JI
0rOHfxIpYaoVhPMXAcrVO7FyBuN5YcUu5pwPvnmnXrR0QmqGHPfYTcuoRgRcZSaAr0Ulm/T7zSPy
KmZavmxL9CeBESw1JBnL1aPq+Pjz/bE6A/0GwqjIQR1Ue61Vh6rEPJcnGhXWq/bXVcSyN1fjWzdy
DxONHYoMhv+sGO8WMKHnM1I9/eTebtCv+7ad2uQeiAI0BgC7UZjlC34GOe6R4yN0k5i3Sv0XGxn1
vhbyp3CjMT/uLTM2ayB9oOUAWAa4bkJP/Fl9QRe+BcwIqMBNkidZw6FMJQ+xC5KNIreFvZUXya6d
qOFf5BNWT/ZwBERPE107K0zqnYdworwH5g2vJD8xYO0kuMs3dCeDkl3qqiKHv9hoNrjXVUqJxf4+
SR/oIPIL+FsbCUqTwjEHLyzkb6ytRBVs+eCvtXaPgLRiDIEVj05L6Zs3Crbv6mJ+ow1QRX6IWQTq
Z+/S1fr1l7Lb7GlX4LE5rsGTEOPDjt1Ha8Tte1Agb/NjogOB7vo3tuMi38vRRVs6ln7kbO90qduG
j322j13oU+Z+RDKGTyD75VMPeRydIm+jqIdT2SmiahMrh/hXOAxB9ObGLGBARJ2iaLIqvgPbwGA7
ib0dzQwI7Q+pmkzxtC88R0SzM6uWwKTkiU1Xvk1zRjkBKKQ2Gk62WJbLotoB6gRR5XDKp8fxDbxa
0DmqDMgToZdH2c5h/OIOUMbQp19eBrfh+stKm++9Vv2MUKqh2d7Q4faBeSFcarHFQ6+Nq/vH7E2S
aJNcwkGULbhdg/xVCCXFo1X4oE/MDV9JD6an9AUERmMnH8WHlCU/2vYFuF0Yp83k72O3w241xKNA
OvhMJlCeFAnS2b5S9xtjsPtXXR6OYygDxpOtzcooYN6nF+NJwZm30tl3TmetkufWzczNCi8O2CMN
I+CE62gHWu+ZJ8ZiwztrYM1f4yKREGp9KHI7LqMKAUp/paQwnIl0D7cekj5rb8YRfUX71NBsxU9W
les64D/lxmHBjf2tpox2yUWoOZoF38JVuFC1OLLo1Hl4NHVM5OoArggnRv0MGmyltjQSxEN966jj
2Iejo2oj/9jIiiLK/17e3+HJ9H1Q8O3s4tuOucc+M37YomdE+z73CuwgPrBGKc0MW9NPzvjft5Oq
wtR3v8toMFAJRLXeryARhJTYkvuNjn2ebDeKC9kbCyD/wKuDPbFTs8DbLS9pTe7sU3FkrpQ7UT57
XFtLWh92dcRWoNLjNKzkbTKziU8h9JQ8YXxDh3BAA/R1v0Y0zhUdjCUy++RZ2X44v3rP+Etc4qWV
bGGU5uarzKk9PK4eOzopunN/UzbCT3AAauXZF0lncwVNwLnID5pWiBnTYCPr2lEwvFNpjP6WfqJL
+uKI7bP4noqO98gltbg99lydhhmm3BX+o9CUWe9UZ49hZKCP2kJqr2zbn7QHUrKmfBz4v6C+KjJz
4SDIItVaGlUWNGRnvqKhuAE2x1GZtu7031Xa7Nt+yp/9b/CnLdD5YIMx0J22ygrGwYIZoRuQa3oG
3iBTGhUNkrz7hZIeffe1XyV8DUw5gbbcB4iaYVXCXu6I/t7HYSbmsTJJdt+y6H0y8vJwC2nTd6uV
VTwd97ouCv+U0+lB7x3jarHn9fT0RJoMJ+z93PR9GjmDWEyWI6u2+5yRwT3g0s8Wktrm147Z9YFj
8lPe2zBdRc8gB1jSWf0acydSN45qq/fUsMmLb3SN7RUNzm6LT2k+5GiUSNb7sYhO6oEnsej+/FS3
Sx8orauGi1NHAWDUbZdJ+nQ2EqEWSHF89CCbf2m/UclxnqL3AiGiZzFF3fK5+xLm6/QjwEhVPDKQ
7iiJWy/FMRxK25Bc8nuu2Q6HIjYgNqXbu/nVxqVRh1GJvBLNsfHaEFjYCvKbPpPhWBzLE+V3AFyu
18yyz3yyJhOa6MJXmIzWHkFUxv2eGgk9QfmeQkQVfwi7wpmcRpnnscRTOC7ImF/n4qhjcERKSukE
HhKxQg3pqzy8ngD1CNd0EcBSr149jAiA/DudhrZb2UUV8/h1gR1+A6aq4O0AjnMLNv6RzazksA7B
RXRQWxn4tkyBWZgd8NwhnpEnxJ1B0LUbXORBeDTNk1/QNR8KMWv+GSggtIR3XtXNsCwHE78Pop3+
Y69IAv2Eo6yYS5oHi1/bVRms00pqS2JT6ry+LKM/YejTLLYMAt+FdyKg7flN2T0InM+t1ro4tjOt
bG2QiGtgFlsHEN5gOYY/G+jmtCzXJmALpopKiC2LRAeATlfD7cB2q2g+XtxJit2wPkpvgr2DiiQn
D1C99EtzMXb5xXANnsID9XyuPS+Lpb+HmeqhNXS/Fg81SoP+EhYt3CIHpQLjBS6RU/4SZ8/bKfv8
rhNhXTKHXKKVOkvmZDc3qL0qx/QOU9J0cldf5pEDM/o+LNms+FFNB+iRrUM5lw7NngU60NB9JGfK
UrAHEoUGPqyhisYTtetdrBlFDAlNF4lw+3seXZN1QekgIJFnTPpzb/H/Cx5rCXaeJQlOZ0mEL50c
DMTeMoKifj70/4nFXRmGTwifvFIIn9CIEDbtTwP+umlf2ORamlyfwXjpe7WYZUm32RKO80vOY8Io
fY/3xjNXV8R/XPjZqTLRUEbpDzxZRAc3e8ULWCx3PXHfsYbQ09G79nU20Mdq6OKq2InA7rRv1d71
T1A12COip1bPW1VUCT9mqz/lh7SbpYShg43xbFt2+mcN0VbI/QGSy3iptuAzpL/YLzAFOQxTtbfX
pKPke6xiq9w/H+pGXjW9FVcIEOndp3rRA66Udr8NjSYaL/IWpdGT0im1bWczLZAO5fIIoORo79ec
StAS9Tk58ByqxFYiuY8W181LlaFsyDwdzcHHDOF8FWBwZuvFmLKF237UkX+rj/SPG+czv5pR5Ttt
Ekd/hMrTtAs7JjBYgDL6KraWJVOdZ0C06aM+gtivs05LoZineFxX4n/2OBlHAgt9fH7h5hIbNtEa
Gc2Ku5574eC+5Rm41ZCic2rF1Wyzskvt2LJBbDjg0IFsv/MVWOwRxIMkQEbfF42BDV05cdhqchuC
k2b2cp5jsWIu4P+OonHnAvrmgQYbqdZ0C+6gy2bB2a2p//HLfuK1Ps7/QhXtkpPdoCw3Ix8GSAqj
K8hVHlxJPU/o2Lv6YTDk5+F5RsCMuwtJB3v+7RB5JORCNfabzzgafvYTpY1D++7Kc7/QTfMwI2Vu
os1h2kAkFPNZOni9lf0aqNyvcGRjLSv7yFYijAi30gK61RzwUPAklDyx8c9eebyX7WJvnhKHBW3s
ZA8jWrP5JlRlVqtlBU2ZQrziMn6VMiKMwfvbRvDe5/KED465wpyLZo4lCRoDBLZoWFbZlU47HIbl
bXAdRho27xZdU2lbf0+bDMatbkALUc2QbpxZJPtshMSJ85LdxQqWtpwFV7yYyS5kQiof4cLnKGwf
xvA4avI6UkFWEWeNTmm8uRifcBtC8uvNA1ihMrNygB1YstxYeayWQo1zx86et4cGWn9mYm8UFbHO
AA+LwAusBUnuKZnXPH1jZ9E8CuWY8Qx/Dt0X3zMiINk1qBFIE8e9wodd4e18v6Vp2xZiZHPp7V0e
n5wib6Q1Zn/sQuq0L7t0VRG8H0Sz9GRfnCMEr8prVNS+M0UT4FAit0lcAw4QwqyFMJz9VQtRzdv5
t7EqBMOIegaH65zPfM0epXZh8znxfoSJalzN0LBFJXRCpWutmlG72wc8drgGSDQmK0JbOkH3Q0qi
BPCZ+c50gm3qQ/mH8meFXxVOgrVd5bKcL4BDRfR9pym8v6twTvOeiPumf0vYvykYDNGAHl+8iDfV
qE6lCeyRrGBIVrxPNpQOa4PGuru+KZOW92AGRM16pEemLrFhpGVd5uGCqJaVuB8vETfC1j/KVbtd
LTBVWZsdngibpzKDMnN9Elb9GRI2qp5RLu4TjWx/8umXUqh7Bm/H90i86L7CcYie8vYMEtprScJ0
qnAf/X2fZSTQYdp5W/OJqAuSXqdz6kUFnzlozi+2Lvz0ou4EOYTVAqjVxsebRZlxlleg0CGX6D9i
T8jcZTa7cug6yJM7upok8ZHJZtFgkypyuJEyzNiETNa+Y89ErN+K75aIQR0n5k7sqDqoMM6GgVER
k9OrHVFAWDkESxdL6MS7MDF2UApqOW57WDT4+JQhcYqPwOukFsgFyUvlTx6dWO8e1ABjKbDMT5iD
7RtupyvVPUlbBIIPu5cJ1xs/Ed/zEzNKxImBae+LBumvDacB6pDBP87RfmLbt55OIAkgDxtPilsE
wJI7SKKFbjd9KZnC+x6dPw1FL7LtQLhl1Ey8gBXytGteJ7rzHl36EAIZbYi6YAAJkk2AS2SQ8s0V
4HveqRrD/NSa3hk4VzbDY2Fhx8rSON6InLXa+I+E0CSS5VxsVVKDf6tCNHiK7OXY8KeX/8+6XyA4
A7vEQhXmmDI/Ec8HWpJXJ+F2Z09KbSUvR51eZxNkA38T3QQzWgaixIHL9utW4+rSUR7wngCrqoIQ
oRhqR2yn1YrNX23k/GFBKlz8Xeeu1EZzCPEILzJVieHE+WGutBKbnf2d0PlLCfoq8a41CuISmEw+
cahWu8A2x9+zMPjjerhbxxBkc6xrj6SV0M2HHlwkSnLk2aMCjp6QQn/NUlYsU4Uu6wrietEGQzJS
xZDJLXQSy1jeaGsPWZbHnDRkIY5THpUiP8YxPUWt1aoONX8NOMWMQJwsWsprH/pLZEFYFaXb2bcW
oMuMwVASkRKmp1GKxKibOhNfQbImBscYEvX+kifQfrV7tawvZ+z7nOniWPHmG96Ev4RxlSUquK0I
B5pVNH2PImuMSN3Oyg86twC2lGN83jcn/SCoYaCEFtjbdrglmPzFOjhGeFHr5NkpdYKkvED74S/P
VOoDVghk7Y0NjIrpJDR2eLzhylnpsj6jRMe0JTz7Kv6cbLlJevMxAEkXlaWbGsfqJosxh2lTDmRH
JGhkOG10fijaExFlYyySohSNKfzFg+w6npVH2Z8Dlfk1R6IzixZNo7ts+pqzxka7BxhOz1unjqbf
yqmgL0Z5kw6JiQnOIWnIP5+ZIkVwHsuvGnP1O3O3nTGTVOPwaxBmsyQYxvsMCsO+IJEkXU5LUzd4
6zFTZZOTTxcqbxZ+/ETCsnkQoJzsSX7Zo4DXnXvLi4adkuLZgTL4DWfLCeQ6H/qR4su626gxNUmu
vrjshrVONlJX0Id5z8MRIy9vpWe8Xn3n4RvAhfBR7wGCDsqiDvD0c/9VJza2m1VWh1moDdyZdwFs
ahBVzI6VQRQOXsmJHrkX8AL2506oWG7ZEP7cXhKf/4aDEhDOdaSBuYlpW+xcWuS3wk9EKPcUBu3a
W9Ld9wlBr6NB61goY7/CBYAwljvxm3CIDVSOaH1L0OsHXYwJvR7d/HYmZGArcIyofRIqX/zoZU54
6oaKeydE2FCLmd7wADyg88wBnCxZAuTOnGYVuNwtA0DjDCo1ULgA/R2G/Wr8aa15h8uytPSs3VT5
tET38kcH7oCsw7cQ+2Vg5ckU3T8AaHzRuLF97s+Gle57Cu/Hj2UMV727xElvDCmkLQenOQuTw2GX
1uo30KLKKejNpV7/T+nGEL6fFM1ip5jot7pnIEh1KXSSBiCAO+wXVF+IAo6/RKBsUSsAz7r68Y++
apibAsr8NuvreZmyeN1ecT4X1xvmMu0/6x2JrV510t/0m/zOoj0EIjjqUaRQyg2M1pPIr2JRy43M
4k+4Pi8QnMJuHqrNb1EXGiFo12Sxs8fQ9JE+XTJYqX4xugIliWslDitl8W8ckHHzukFZsKw81/B6
BqYEw6YOmZnZUose266L/qhwRs7/YonoCG1zEO3KwLLLnlH9QIUl14APxfBNMSClow1VX6Br2/mo
rEQwRBstrLDTO/X+u50t8ZDuTlRRjw25muDwcZcVDAW5V4JYEnL90iSm4u1QjsAi23jI0nNGUxtA
ShQFn7EeHIzy+0iHXrhQcaaLbGqheEesVMJqZssgAGRQ2PcbrXuLdjb5LSwo7tPuZ4K8Uj65y60V
ndNR+/MFpKh67/4LbsPq9VeHNbqVkTlY/pnXY8i5PGL3dt54S8n49m088LFKIEB82CLGZ/CC2lhl
vbedNpj5GRP1IANC7fjpVNrXFNEL2tlS+mywz/tnx/r1DNynGfHQSYS7efMWS9+6nZvEuk3FUTjI
OD1zaJx+h+al6MkbW81qsg31wNupe2oGgVmnEbKzN+x+MkBeYEW/Gq9Dn7HrDR84MG6CKKRA1BNa
og45dCQqqwplpfwr6q20+xfheK5Md9uE58Lk5PXBLzOwSW+BT8PTy7E3KHgQ50waZdLa4pqmj6LI
fuMFxmYZWvNgvUUlo+I365nRnxw1Y1LnHVYqbO9A9n41FppCgFRYMi9whbiyNnaOVIUFqaWI6m4r
6P3Z/3F/LjQb6cTiR/Nee3HJEI8P2tgqzgtXI7TqcS1xPzA1+PAh574KbR3vIzT3/EcG3Bh08yxk
ShVYrychsQ54YltP8cUP3i817BFNLT5VmdVO37l+a+VTsjuXBKiKqN78NvyObIkG9d0/TDu7s7BW
+66bytHwc7FH4basU54C0jopeA/4a/sS3yJyVxAmqhAiraNtq0WzK/jg9PAT+pM5mQzHGf7LMnyv
yXiT6UHihIj7ZU/1VRJ2BScZGoIHhJzpGtCLmTHmhH8i/GbAEZrxVNZmviyfApVM+y/mLxDEVTl/
hJ8bq/Ig+Je3imHvoFIoQ6L4eb5AawvmEAnJEWjbcb2piK8zAP35NGI9jzcVEGCWYVkM5Zkfnpkj
peLN1qxZHRV/6qXcCg5rR1jZyfsllWFMBZuXrQDG6fA01EsNkQRfIQh+b4J07GV/vkI6QUjBOSDC
n8szMRJFVeUNDtfI7A5F2i/CLmQ72XTwtyAmisNuPNYFvpiDmivgO3vJP8Vdm7u49C+N1ZZmb+6Q
5WfXLp0XztQZmK/9Kd9hlJvzp6jq+ONCbgsbxcJ33+qwIj594uXjWJqWrdxiFXJ6US30RObI98Fh
nkLJg1Udx3oatlY6KYz9hHHCYUz5ehYcH8IMve1KX4Pn5RVlhlKHw0LxVjhh7zXhPEsolAYN34Vn
tdwbKYERY/ABMLytcUWwmNGqJw5ghCLRnK+QRPnONjoqbiAjsmjUw0JoJo41VL2y1VOj+ufM5ePh
54h0rycoJmzQ5DVW/oc1k8FNOVXRXY3oiamOyyLpxcrmprdgm3Z1ZClHKOm04Fe4rdiHc3kosrFV
G/YP6LAcEDaIcUZ6t1++MpqNkT8GKG4pLqreFq2B07jzjjWvJ4c3j+qnMlqzZovGL7L2yF4u2wY/
XMzl2/YdEXNVYcAKtfv8Aj/WNrbCfcPzfDSbxi2X2M9YwxTWYLpTotQlwvKNt7e8JuwkW0l6EkdD
AHsyhq9ap3cGVjK/T0jf+6WSysibm7yQL7cP1vwG3s3zgR+4zWCDA4xzO/XUSNC+e5W9u5Is7jov
rSaU3oSADRu9M0W8/FYUBGsnyI3TqWMsaFKjv55R7AXZLXkwY+GkIn1M4HHXSgF69zHctkVLoPlN
7OiDiOVuMcPDwv3jjx+oHOAFkWW9/MOc6VdEv7pAUEGHLAYokgrvRAG88ozhZi56fYhpZ0bkihNz
VLtaIZRLqQ7Uce2lAvn5NCSo27cLMkzoXu+JywZA24LIG0d+XpRJrgIfgg+IYjgcWUYQXCWvUY3w
kdF3+DzNnC685SyKTqo+3fvKxBHEXYHX2UtqnmYSS2gb6SmYxk6dr3hAQPYgaPA2NIFCzE4uyrbb
K2tfuAaoMWGkIkFPUkoFB+Lw1+kY2+ekFZOamLbj5zlAev6wv4/hm4V4ueLprJbo2RYCh4axciFB
y0E+m6NINAqoRMv94bhBom/7C1hHBSPzEjvbcOVMQqUDGHzcrZDpxd/l9wrIBrudE+d/sXmRKs5L
pEH1hCRwzKMUA39Evu8EyuyBazIcbhvFfWR4qm4mGjEPjdVydeS/cFhSpIW5rG/s6e+aTKSgGr+t
dydrWEeyPeIIIiw//IIq73IBmh5CzHIKff51zk6fh2BjgjbzYpYnHzzCScND3/RgeRFQuyf18IZv
FLFAoUYuc0DksHGI45qSWoSdxmmUXpJN1HNgiFJW58NAqk34mikRam+Jv3QNRtIPW5Coyjwl4e3m
NDouR9g5wcTd7935poVQ8NlLkAzYriwAbS84exbk3BitIcOsUN5QgMfyUEGQ5/A63BfdcgffFvXS
7YRE3hdbvy7Uq/5jusaMGPHF3SbPJnDQGArt2ySbLrv+jqp5Pbkri1lO8GpFSQQFCPFQa1ueT7gr
XIuPGvN+gkePPlKI5FvzQnwz0bDq9BzsPO+TfUCEVny3Y9+dhpjin0xlfTdu89IezwRFulZ2H9fS
kLLaD4MHUag5liRGhAMARZlaBx+UqWZgxiJ+OFDpBuTtumMt/OtXvFgKrvNZcchUy32+ewiu28AH
ghafTeOZOoFLOY19nt0ADMIzmdvayz8g75EVxRUaRPOmuSL/pzNip0H4zw1VbEJO9fMP2683Wy00
Pp//yNeDk0VijCJDHTZ50m5OrZhSLJvx2rNIMBunGwHxF2OdKLnpr2jhU+sycSW/yYq1XIBbmSY0
otsgXZ2IFh2keKpyFOloG5nwwlod0oDzCAgPGxqzY5WwQVwct782iQAbPbxFpPsO/1VYqlBD+WU6
f0ex7ldkDnxHbXuHXkJTsW0tv0KfRo9Ah9x+zVlEaSWiVGFjLO9cMihbr39LWR3gdHislYhXISye
h6lgqP67pDu+PBYVAvdzqY7p+Xy8DUm4hP8rJaJ0j+5+aoXz+XVbyoMlVOtxIyAAcIB3gDxCPf7C
ZbOt8TLsAeu5ZlGsNazlfYhaCxtOqpGsUtuZ+YmoELBQ1xCusURtYDxRhlk2Cu1EUyVN66XFn+mX
zVyzNBgexAnETMipW8Tpc4D4DTPXODvpARFygAAdlNgrAGhmhqF5r7Rq+EY7sPvy7vDacs2CTE6D
SKpKcMoqrP804+0ReRcac+Cs4lnhOFvJGWQR1LLTbZBMWaDTQc6zEkQewKmt4ezbrF/wSIE2GPb1
BdC2gXZFQpwDrV/bWkLl9PIY+drSyckx9C8MjuFLkbsS8bSX3jWsUqletmyEtZEKy4AP77zr+a7z
WiohyuQ3t6pau54qaOqce0NN4wBszBxus8g7zwNgTYACUqi5sxDleuu1w+KfxGSsUlzWvjcZz8Eo
ztgILca56edI9Ff2D2qY3y38tt/JOSaN0ecGKMq/pWB5eBg5t4yNi3lvjyS0BaIZ89iLl7H4Exw/
thmPrN3heU3sr/wsxxrnJtcLiXScjX0bJJnQGG3AJvy5xS5t9SJ+mmL7EoHclSeTjm4DBwRNOzRx
TwWbVeCmYXquvfVwOn85R6d4KFhEKX/GmiyB6U2Kb0e3kMdA6Pc8xPVsPiy9uBfQdEb0wiqOIkOp
eiYvLNVOXahuWxebmMi5yhXE+dhBhJrxBH8UdJEdEsSB1T1uqanNVfbAYru2vkvQvTNaa8gHF2ZV
vKVZp8Ak/Oa3SFHgv7kQ6w/p0UjCf/UhIyxVNYvn1hZTqNyGUnIswXaxauAUwMEHRa3zbJFY/j34
3HYmbzNpUSzOc/RTcVdwcFQ4tkElDZSMsDc5MvRFhpbzWDUQsvwbddXld8+uTYVF0rv1kjHOFyk6
d5y4w1NrEx+CO+PapoWSgBX9mi3xL5fQKQbzkJahmis4rjGhAdrLPvvKjM4+4yDbYJMZA80KlrLT
G3c0/HFLtxXNNKu71f5SZEZVDXpvCgRbq03aufBxnSpHqxmZVkgoRVX7XXZOVYhw37Tu6p0UHu7d
3pQFxQeTGp6j8EUqseP0wauue5OjX4P/c8ijQ61HNisZIkS4KvGYsw5I01tttTFJmNMc2dQ+Ove8
sDUJUU+IrRFoiEORJO0h4Zpg4ap/1AiwHOKLNixwO7UCTLzBk7ZIrzk8ow7m07SEK8UJaQlY6iD6
tqbp+UIjxbrmG/HnbXfac18lRhQOk3IunLPraFy3Hq9U8dO2rw3R/v2ppzZhOfRW3/8A/vbZLwXb
uqwr1HMVXkZtugTfjyU6IoY983pTNc21EWxVvjcjhhs+3vZr7LCL9rPoD6Ceh4YNxg2+YCe1J9eM
rXcrMrK9AofNCwK97q0hyWNj1ut2J32GitK/bAC0BCch17ils878Skl0Vvs681OZRsF84mygHrww
9EVo3v6ToroHxOz3jkf7+4EVMZUyM8p2CrCQHD7SRuJTXZ3tnqjb5Zdv6gVTiHhtBeIL4cDRNlQW
XAbORgz/ntsa8cb76GjmOt0MaBy3r208LczzxLMr4qXV21O01nLsF9v8kQX4COEHo/yuYfSfUM11
4vCxUdoX1ji6aDZV1ZEq6MoNmf8ZzEPh2Mn363SC8o2QH6sDY+g6yJ1XXMSruQ4crVUpvi8oV4PU
/3VLt7qkBQfs5myWdJpQZGbkOLD067mo7b81hgcRbFToBHKy+ppSBzg1g6Qt6/diY0KS8dyuT6z+
cfwUtXp0boGnk6b4wCSvYprODnqQoj9uGQ+LCylw+5EpgwqEm8kO1CxLh1U+e/+lkMRaM9aRUKg7
QwDq06Uw4tQM+xhbUFQQxk6oOIQI3DEVk5XXGKhFYZpAp6QFaVr/NLIpVHqB6Dx5iaPppzzZc8ef
/ZdwciW66w/Rl8bHcMegcEmPc0IWMmo5L+lKqgzV1dIURBaE9PoDB9R3g6X80jzLDojX0qDwGu36
v6X8RVcAJSm8r6cPZYlB4svh4evuRwO85JPWJOb9nKU8RO/EqGudT1gzw9sx40LL2fzFZ5Wa2hb9
VUlWl78rm3Or29nvvp+G9Y83mijYr8CvgpPGJnTTf+WPd0DjfTMuEy/9RD1nm/xJgK5V31xGY+XP
awV5IF+2z2P40hjtgZPfYuQ419gmiyPUd+AqXZ2R3d14KclIuJlUOmGH1BUuAuGtUbmdKLeiTiJy
byuwtKbMKGvsoV8Wk9uSZK8RW1IaXFNl4TOGOmjPYu+jJI+q+phn996jWlWH+p6uC6gxbYak6Lyt
Ry497PwdF1WX47Y7Cuvhv+mcDv3sUwn5TV7BKgS7lRb101KwAKCsQ/gwz9vogeB+ONGTVB+ECpOD
chnEpBONPBEUBeM+uoFlG2dPLBX1oL+Eb/QSve8QjJBgQDqmau1Tm2ooRv9+z1mOP9j7Sb3ctvxl
M+XzvlLZytU=
`pragma protect end_protected

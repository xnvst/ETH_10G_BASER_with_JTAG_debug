// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:25 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mJZN6Yz/Mw87BWNOsrAHaIFcwnsYDJSpaFd7B8p7riVkcSlkNDkgAWUxJRq9Z+8R
sr6Mwqbdae/AXKp52dksidkE9Z3lSviRpAJJy3vdbkHIVrqh+hL6tBDr+OHoHfH9
E8D4o5mnIwgb6JJLFFpTGpfoZ76r4UC5FKTmcnUlIiM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22512)
Rah0LPVHhPm4G3NQmxbjFxCro/SoRP7DaQhXkIMrvK/8dfT7XBLt9G7NnRypRqJZ
t9XrHQI2d0qtXW3I47zhn8JOxZIg1WYJ7dxoUlri6hwj4a+0j7NnjfxQU80MSgvG
B/ubdsWnuZjQr2EOrL4nLhmi5ZB1Vy/QmgzU4ebuiKR2PkXhoUrnb4eU5kemBcVQ
jDOQJdnWcIY03VNLvImyqRfEuME9pvH6ybD8HyHZ2n1bntL/Pn+jQCUn52K0yzEs
1I307mjfm7s4qLdbXBYoZVbVryUxeC2+H/mt7DbUcLdmtrLhSBBI6aq11c0pv8si
nfv1KMkYjrYBXWwuiKyfLWxb1Uu3vZwU8CbHKeVUpThc6Nte7SHSgTY4l5S1pidx
exCi5SJksLnLLhOcjPpeXRVYukNIp5RTRDNV3Ta375yvuBx7G/DSL09Qu2m4Rcir
+AEXNGdBzavjpl3dGNxdTZiuGIAqQL2CicK8ekkXI5Xvee0tSCrp0UVI1usBKtD2
Kp+7FCjxArbPS5CARJ/yvOTeIciQLspre8Bi+Y19nKX9OwwDgyYoNGxr2vQhb0Q8
4PM459p8nfxPGGX9yvT4/huoGECqUrtiZUueFeP//75WJH7zHgetLmvXF+3bJHEK
JRQa5Cav6/teN3fDcoM7pZWQhM1sI7Tr+dnQOOI5GaOqUOlTeBTbQfUWAJV0OtHv
5twF38pQgR2qH26yzRR9oBQRDW/NJnvNEjDCah7ACUg3arzAvRCoGcB15JyAS2c4
wwlPxnyaagAJGc119BeuT69xpOfyC0pybCrHui+O6g30c+bNGl+Hq9uc4kqlk8FL
51zb846NXaxGviVNfhtukeOlzsyiUBrvi27cum+d9RBoOmfVQgSAwPJ2fxH56TBe
m6kNIQ0ycs0+6XQWlvd3jac1iWbL2MwG2hzr5rNduXTHPzjiSQyUvFz97X95qqdX
s/3uLb4ityGxFZuK10y57Stokskp5l5dB61L10wNm45NnJ3mDEGA2KUMIcM2iBt0
oOi4k11JI/6v9a3xrYgbqDuZwpPBGTYank75C3HVA0WVUOVlwPqiH08XJIseyUT1
vlCkLF8p5w+LvJVfumXDMYCtdicbhlP26l2tVrEJocb4q+RKBU9Rwp+RUeQayUBH
ouYxfiURiWB9zVXZf9Q0EcPzLy0WCxjvQhWyDcqp1XWrlj/+41IdrdTo0cV8Qv0i
RHQyAwW+tm+kkKpl60HghAysdHtkbFXoFEdfoAEuha887ktKTGUgEiy3to3vjV7W
6YqIOoiR7eIqfx4LDIM8IHhO6wLw0Q91KwSpxkUF3xMm5mIBGaBkDu8GoAQDZ0Zv
JHiri409UlcS9hVmx/+rlEEx4A0R2wAb9ysbo4pzTkI1dvLif0ySAhZNc0Q2Cr+U
ZQ8eml56UbohRw9HiANUROjj5jY2v73gLXu3icvfDhTC8QIwqQr+lfFQMT/n8u38
rFqCk6ozpT9YFc/VAvVka/FlDXzELqnKhp+MnN7FOwKuT27vsh+2wNANv6j4Wiwm
0lo/55P7G2VvdJeov9WzRf83vvxB9fnpUexr1FO4vAiG3meTRBekDYzsWuozXgHG
GAfL/Dqf8T0J8He18cfQkvONiprNzPAXKHpE1Gg0yRTaSyXd30OxCLiPBubngtSc
txWGV/xyYyG21DkjUpDGMZ/F7W9NOsg7fyhuLduGInLecRnLeghr6aW0LImCbrLw
Qf+Yu9K7DIs2VD0aWtDvTR2cNVwTdufKAsvabldYMIAnASIQrxxPUGTv8h3Ibob6
U1KY4xY+oAkudGuVn4O32LJrWKXVRBySkUkfp1mEa/0OUXTNNZgGxSFpbN94rOTm
q4/E2g/XAJl5B5LOKtUHy4TIUVpxiGwvYv3tgDOzXoPD2fwXr6G1vm6D+l4aownE
t4UJPGKyFBn3Csb+TSQRP7vSMIUuC71F0r2wPR1mLpkwQYNG8mZnLoImAsSw8DI9
PFiPRbTeCwn6IjKhNnef1ukIZsPPNAgtsoDuTLwU8JvrCitL8wqh4HnZNPqudnS/
hWuypHCv/ZdKlh333Kx/0Ni1n3hr1dSgykqKsRNb+hHTbcEAWNJOE5vLL1Z+v3TF
BQRIjd92CJ9d4n9i+nt6C3i3e52+ZOAeJ7ZiDIzh6xHo0mA5Ok0NQi8HUqEAIjSo
vyf49uLGOKbledJtEah89shfijlLZtGgre3WNssxajgYgajDrzcjBhh9j82or/UD
RwhBqigiySB20boNcjwgRle8P4rcGhiEOF/Go3+liZGMZGL8M5wh3h2OzS2DgmfT
YW26bw9DnzuOAM7mLnf3/XBQVGa8uFePvP6rsDBz4M7xFn7HL0xQwYpP2+iAtkKF
x+czTrP1VBjlidpB7p8kKoZpYKl9FlUwlodBV1/Wd6rC+Uv4mvkd9NcpKH6JTOil
d+VeaIWcHai/M0/Hls9t6m/1BMuDzkPoDFtQXylWVDIlwiPq6/BgIXvxIRjA6AV8
hGl0sgAn1CzqdCDpLmAeVS7RbOxFlO+WTSwpLq0lLWJMRw/HFNnNK7MPBfSQB4YU
yIihufIucKigaqlrtUluZLVWCfZUJ9khayr+z1cGfGQ8SyqPAPAtd235hgtK5n/Q
nS/GBFMfJdZ5Nsyl5Zu6v7QwatXMUjHHqWLhtrEQOpvkqxvb/8aNGuauhh/DVU/9
1MsvQfmPaUMKsWOZsC4qBQwk4s1w4OYHB8CaGtgtrVhbe5XAQJQ07Z3G24/kQ21c
jx23JLLl0MGfAEEbLj0HQADf0nITfRTA10B8rbrpcFGL7dj62mnKw7vqCE5sT1n9
qOMTYzNj185mjKFZfWsU/ZsFB6wjC0H+wA11jwkrBjvpPR2cV3J/tNCqlDUap+uP
QeNwZHT5pcwie0eWj/wEOZZUs0fYRpWv7RSKH/lZyTIj7k5P3Dw337rXd1V8eBu4
ZmZrh4A2hQpJbTlTTIJQY3wo8EmwMRtesdysiuTRJdSeiULa7Gx2kQ1gVpjR6az6
m/Ztfrou4NL6QdMZ+6GVoAHhTDTucaIDZSIf1TnKktAxUM1evhpvFlA1oxSLOeHR
Xb6vD4+Z7xfEEgbiafYYAwanLt0A45BivURy/8804iHvFpbHCP051tu5KVq0ygPB
bAGDA0S5g/6NJCsdcZp+W0U1VxTwNU0ZwZKpEXGuuqEBpEEcf4HdVD+29AzqlQrS
HHmc4VmiETNhb7O8H2NeOohATz4TvOvCJm5yvhm+E1iUCTmLZ3uJek7/aCxc+ZDw
C43mE2HiAlPH1xe2kYfqacR6nLRqeuBxd35aJHkbJVSAJwUSpG7VMdlETgxRL4jQ
WE7L6/F9G2yPOQwo+lZmvNtJmjxaN9hgAGcJNPYBqhflc+HpZUn5a7ULH7aUmTj8
0DnAvjVXhgAVOZFgLuFmyxdCTKZ8ME3/X/UjjwqU40qH9cEUrMLhPGxbui3r8WGh
g6fneFldsawC8bCuNwLmMNuTK6TXC2ApGs3+nUq5xIybgsqyGdNzUsnxFW3plvdg
GfQqdVOYCvy+ZjpzhZDk12n3vWaNfc0flJ0OtV4qqPs0jh9yqlRKqgok6u+78Epf
exaF4mroNEMIi0//DaNxcPbREfD3CA8jkQOWYTNEFMz7tFycCW5Ucqn2K1glLBje
9vjMXczqJDicEv1nao4B5CkWqA4pDpHwK4H30fRTgHCgK/Rj/lYXbwsO0+f0Y8Sv
ryhRoCu8mhBxibh+YoHU94hXfrvmnV2plBi4zXplquniaLWVH8BdZxB/6L2iQ/ue
BEXXOfOo+lRq/ylo/DUtS5SjLON4CQPtD+0a5QjpLHkOM6c6s1/l9hxB4j5t4VT6
aBPGzhyHDa+lELBhFyqzDa/g1/gspXT5P6Rsc++LwDzGFdl8i/i9P780NV+Iepoe
4P5vXKx3ACZASTqQvO+HyW7++tJQ2jQ4QskAD0zs2zTrOntgIP76SZEQpns/qxt9
B8tggleiEbyGVqyRSNAdTrQ/x+frxoME2PM4eJiZVfkkzyQnt/Ns4ByqGiSTneDG
sYaUvCsDjpKLzOVm/vNhPG5eKM09gTtagjsjE6/sItM06O2Sv0+SvHHA9aGdMhI9
7p9rXwrRlEdu5YCd9t4QWz2ekMTTtEhbzuL2B9+0EFvORPHC7aFBK61rW/5NKIUR
VWz0MTHsIQ27qtH6wM7Ij4/GZSdE1xiRBNfxdBE14IoNH+V23m35ns8+FCQWW5D4
+Z1u+85xkXg7GxHR8Isog4+n1W3HgUlbsna0dYNGlWgdQwpNYN9bZfAHboAMuSTS
CEIbgGuy90ihxdPD84e8vbyMMRyzGrQXxNEX3JlH8MrWaAvpedtFQw9fZVAayO2O
G8qaMe9ZllIyNotqfgGamnauEL15HmgImn6nxLtvy1R5nVzgbPCfTWt8OmDjMxQp
7p245eOYFvlfGv/m3XPgY/BQvNwTH6RaJsh6A7rZDfr9HjkGcKwpRuz5fL66uCBQ
tt/duZTZ1rGa+bAXsdRD8RKA3MRUW1FECahtWQJXfrDS45tGzOFlljvjSgKz/ea9
QiC4yAf3i4oWMSWtyNf1ykW0kNztxi8I335DzHTMmNhBhfIma2q2OHbLoFLQ93t8
ULBK275vwm/Qv0D+AWUMcVcDEro+hKus/ieAkg0QhBmzDmT0FN5ZzJVPftStCSH9
ROWBnFoAo5mQX+YjiGc0OV7lPhYUSgt1gqskiF20qDY/v0/+lMDu5rmCCZJX/7m/
CSfthtK2raKax20Krp1Wnx1K0C37EJmWamw9VDYTMj0xULdDRlQE8G8nAysDvK4B
B9L0oefBrY8GUMBiF7SfG194esGMrDhW2kqbX/lI/AD5ps+Ex62lbfztoogxE1UP
FOQ+W+mgGK751iVLzD2GbUwiNBtaB506sYuQndFM629fh79j7dL2ZbRWdFXbDI/V
/ae/cgdLPnRYpkOXfmOgJRbvGI13DZHFl3czS6HpSciyxPtaYOruCwLCr46WDDAS
/pn5mrWQryLxgO2wo6v0WikdzUhg1GINPkHqcmcsXVRVLiJJVV/N2rfgPYxSYT9J
nFOFaBCi1giljlZICfUdGsmlV4UCzsNQ3vxdg71vLHoiVenmLZSpZR1xN4OMPC1Y
KVgIQh2HIPrS2JT++Zo/ulry5p4eqvUjrmPCcQPGamcKiJz/W1RaQpr/6auQgWxl
KJxGvcAmG/vaGHSRjLOEIuQxevus34/J4QPrHLooWD7kwXqnyzl8VwfKM95at+Ja
TFaOi/AVd+YWJAN5LovshGPR1q2J3G4dVZbSZoQfDqR1xpWwGSYupTiwgAli95a9
BmiXV57qsdm1GfSxUNFcofanMb9ILOTsyqfjWRPCYC6zYhL+DHzwipJyt/alz6lP
Jpwep62L8ygdhWL3VAoB7G+vfqkJqcZJAHB15Tb0md4JCA3fETAeQrjMOITkt44x
oNB2jZKBk79cv0IbxyJKhdnxJ05JCyF8BtxSPohpQDoYGx1dAuAZHnSsOdA/zZQx
60Z9dkxKRo07LLSl7QW4zrB2zwQbHJoz7IhRPMxfPIkTsogLNSrXFCk6acepUcH3
2udYOh7XTLanIEBzvrXFtY+Jw1hoHDlHGk8c06wCzFSiRNUhJVHeNS6ODrVCTzui
SJyTgAuPZgC3yRWesrsmTgHpK5FkDi7rjdq3p9bDsCQldOYFzhFYtXr+sXpH8nKE
1pK+MnOtSotsbErh4Spq0iUmAemPoOD58N43NbUyl6Q3xkT3TOzzYF1LgRV12kKE
HfNX5uSpF42Kp7eJdq5zCToCvHfHaXYY7cro9iy3wnLIbSR+1rm10mfVCeaWLXoA
rDROXkkmXchSVK/CQyRnOPP7yCl2c340RUN6GnidRqdQcgaUnB4zju7qqDCtSmND
nz7/B4E3dhRM8vvhwavqVjOIrLUEuPSX8WDFOkj2pWund6Fi4fFCgiS+aXUuhi32
gimDBQJBtECQnZYj/NhAhL+XPI6oAndStsdLuWaPWblWhGvT5bSyn4ZH6zCYspIg
QniASf2NFYFPJ+qMJxxQ2ROwb4FKsvZgHHe3MyAN/EEC78mRH3gbCtsMaEyfAHyJ
XE5+AOeiiCZU/q9fzUsrSGSYWoHQQIgL5HCgaNraARLQsI2+qCcj/zJqLVTFf10p
0VStjZKKycEjxGzQiiwjvHZorF97Qcw0f11X0BR7+sTLyASnX8ig5K0Ur/QsiXIf
Lh4NgMGCcBUpnX8bK2nWcAn1P3mX2XL0nvoiM52lHUr4zIr6I7eClDLoG8GqfKdS
M3LLOJGmgUVHku7vjtcR6s0ogUmQBsKF6t4XvzlccZXU9AOcXRm/3wL6BEqJwhC+
nf4bsnEtRM8AXhAqgT61TGe3G5MzBOFwonkEbSnVeHLxcg1S7PYZjUByxJMFnhVK
zfzNZJ6xTN+6JNS7S1WLGMUL1avBYILOuDHimZXoBKd+wxjZH0QJxq8eFr0X/SSU
cdm5UeCAs29RN9V676+bb8yI9jJdgf1O5ND+5BDFsqbyi03qkgqgs5YRtSgzjMx+
YKBL4LgRG7kkvjNlTmlwys5zAlhCaRz1HfY8qZuFJScT7XXcqrSLfWQF4a77XECl
Ggml2jKUObNMKSu1s4Zef8muUD8/uO6TPOo2ic/juOo6W7U6CjCRCtCRW7VhQnKk
8bbRSXmpzyCq7fwBi/JlvXJ3y282i62Jgh2yk4csy3BDSyuqHdysp8goeMLF/6At
TCHWflaiTZrwHANlgJSu4yd///f4vnLXPX6gfpfIO4d3X/oUDGVqG/aUWTMJw3IP
5Q1Y4Er2v3/q1WjVrh4C1AitcPa5Yd6XD92Ecjwht/yuhUzfDq3ykRCJCwxnCGkn
6eNO9vbyEtq0EcSiNmZodWiBukEvbci3AobG13T5NsDEEqGkSTldoBdAq6W2rOBn
/3zVnf0u1f0uuHhBtIOuj+hQz0G2VGG6m1eI1n8iGsO8OKBKC87MTBogqsjk3/KQ
xFgpILxYTvlO4MGgAgDsUwShfFnejfpYakP6dQYKK+AZQQHdh5T93iZVJE9e0Cdu
UAxedJF2jp26pM7SBqhKinckeu1Ui2+/AnGpVjYGglY7Q8rOxvUrCILDJRBdTCak
C5/84nYyALMfIJWGDipaF0MToPQfa4LLtigdq5FIrDltaxsCoqrPkSI1JipR1DlY
JmU8Du/O442nVMvG+wM7IVkso9y9+GSP9UWg0FKLXB2tdHL0u7msFJePQYnKwyHi
D0+TIbee1ABU43Mu5BN3wlAG7bjNQyeBvTdM5bqqy8CvOnlwRcORg7jlQJ6oiJMX
ANkKOuNXvipE0Je/TNFxe/rKE5U+EAqJjwNEknEwbW6Xf4VNrn+38RCn3W6T7oPD
kVX83ZJmvomDhiy4n9r9Z68zeMVY+j/obooD4oc247aDAPXHNwC1Q91z7pRSmHMn
jIMbv4lZeCG8E6iiaWdSco2/VEUY18YuSjlGEn6IaTb1ZCtidBXq1vAIIggp4DUo
1VOrEMTZhpxs0jkgkUZEZHIqZxcbqmYr1aT/G5KCWzbRJbsQTKRXgIukqOs+tdEV
IOG2MvjCEH0M4kme/Aq7g4qa9aPxS9ZApWFVJVOq8imjhPrxFkBI9Wzc7otw/jqo
dKbGNGDg6fyOsfcTufeN8S3VCU724mQ1R59QMnc4DDAXNtFvNceuN01C7+DkGU5+
XYuq86X30piV3tXqtkHu5IwMXUWK+SCX47yestRJNVdGIdpL03kUwqIOC9Tdk45z
VFFQb2i7oPB5capK7/atsy2rxLMjmDQJo9BUgJ/uvppHG1y7qiiGotSQjzfd5an4
/cHH/+Is5nkSqe6anVirBxhfhYSr2KpEVVhH6SZQx3Cr4IQUON0K3x8Qj9BqX3hF
r1hjsFnb3YcK6+ejBRTZhSeR6I3Te8c7Hax8dftDzjEkbyU8vwWznNzgzYYb6+hg
ru+1/+Ofc6I7UOkPQ2EDfOnzTKaBkPQ+Sa171/IEqoxJ0jokHVnjrdzxPmFFWwf4
Cyz8A+BTWfRajAge+nKKIwDYWm8DD7ht6SvQR21DT6FF4GNYFIL5aJR5KWORoKmK
zeragUfxDZvzeOvVn+3U3TTv9B507zcp1vNk9jtbpoaMRIpdSjRzlkrW9WUjIBzl
mVGSrfxZaB55+eF9SbOMQp+r9OIT+tzvz/Fptjfj7FfHg17XJh8+P/fQYfhPI84c
biFL62mllVqkHt4pl39AMTorP2a8u1KFS8HnK5KhwbItyYzA7ScaU3BL0+dH/cyf
9jlh0XNGGUHMnWF2r5nkKRHN+T5EVaU7PwXPbXkcFzVsY5vgmDLgiX1JZBnURQPE
ACbuJIvw8wtX4cUX43ya0yeZytcBH18KAbKeakzkBOVaZSjF4bZOYaisif+0ejZt
LYhLc8nW1B+7hrnIlQoN0vXlijuyC3hHU738KwTyExhsIoNLg3dLdObn0mwYV/gK
OWUN5BvEGkOROGAPDJKw/w2RteFvHfOwygzI3qA3nI1zhTIiiAeIFxbVPeJZ6z3B
zBfLdAA4gpMvHiWpk6Tr2CB2T3LDRlQgBAXDKTqawnbvN539FtA1TtpN+cAqvP5/
ya+Yemz/eQdGKW6glpDqQrbTXLYpJaiWubDkc6jWBUu+zx+ehLeSKuJ5Z9ognJ8k
eyJy18fysXatv9sCe816X6LZ16SJ7xw75jTtcYrgZlacqtRA28/Qs2xKiY8rvT7q
tafI4isY8eh7rReUGbxEvANxr6DLJSpZ68TqIL1IyfcawLGJnyFtIjwR6q8s6vuo
r68vfFtOl3BVR/1HP0VPbRIeB6UO9A1gecWA8b67UMC7gBOSutuYBXLG0qhTBOFf
kcs6IAD2j0tTzFVzv/3b+BJH0M9JcD7l4prKLjpItdYR/0qIMbMSMv1n5dP0PLOM
R1GiTD+UK6EIOK3+xDdm8qnB8WghyH7tJaxzPnzbpKOgvIWzBqzOkS0ogHBM+ut1
D0UkAHG/eI8ON658A6s6u793CaHm6V7eManiQo8z5aCiSwy9Puf+FHqKdyMMCra1
mLMrxUKdy7EwPlVQi2yqUci1gaavz8VOjaQWoHfAMLTmuZ9ZvT8Wg0sW0Qy/Q531
OxrqY/s58hrkgNKeJDwbmxKXh3zH5jjAHXFYzz98rqOjtSO3eKGOuJeax/fMfZkm
h2vVRDmbSNsticLN08hjd+4o6bfbfh1d3NMcrdLGd/ROReOQrtpyExhsNYMIWunf
dfQXDqIgK9zZasQmMvEOjKB8+UbLyNa9Yo3212PzHUYOyWaMh7TuvgIUlcLpCobm
/z6dj7ym5F149+Hutu3WPZgZXcMtbu/EnlrRCLInwNhyU7rBP8/3mERjMen8bCq2
jXa9ncUXQ76BSRn4zTj/U5QCUG2YlmJ68vMR03rKaXSadFU7UAB3bKMw5VGIzj6K
Tqy09qJYpDwgHqJ+1pIhTTaUrok8BlFPLFmaT9fu5MCtHuVn2QY/LnkMUtuHSwzI
ii45Sa5WSV85le9qF50l3uHn6vLqMmsuRJ8scHQXsBZdkAB7mGwfiktnOHP3JwG3
UEXy1LEs3evuWHxaRGIrDrsfaJub5lY7fRhtb+tGdUyVYF+iXr51dDsmWL+1OADc
Nwtio8wYl6epUvejmzw6Mka1CVM+NHOn1EWS9OZDhbOWrujR+BorXryCVUW0hmq9
ugC8EYfssSbYvsqQY6nazTltL/7qyfEs8DfRehFaUCPClrAnb/oc1tZWiPXysQWW
n1QoOQXKSGYJs+lF1WPmKFcb02hQgCheZVcOXPN6nB2pWIpsENYArgTAsnLaqInB
JUHFcGFHT4u64OsGk53lQi9JacogSgSPzRNWfEaWTogGiaSWBtSsi/q8/U4opoeC
S7IoelDCd4BBq9CzdE4ml6md3592MD2KfZtsfiBLhCk9YGaFUHnoUE6Umq0ZsNfF
cywONiEgp1NMrHSHMMtG2xB4jVxKR68bRktjDtIDqtuSwTS55stKMnYumSmiIped
PZXliSNaXxYiDUZVJA5T08lzlZ5W0Wa0nHlh3XDdiuB+DN+5aHzCfTNlHKIUkEn1
IhQ1U0GwGqSUj1ZvXAnYdQszNicG0XIbG8AacH0/SnT09TeED7sDO7r3W3w5jL2T
DzU0byDRgRSGUDtFvXsODcprkZcVfS38qSJuleQgxsHPTVIubAjkqbZxFlJoUAd9
8f2ovSpwFky8oYCdreo4ZmI3V293wMW86ByGhugKUl2kZbQ1eE61UiG6s4alXoE1
FsqKrPgLHZ1b8IfG4RqnymWEDmbNLbs8FF+b/s8iFLgo/JjfiQeow3QPA4QNROq4
gQQti1iZMY9zHAk5DvV4jNAPJzSrWJD3qh8QWIvghOOc5L+quAovZuDM3f5GZOHn
Q/5hFKprHoOZ/uwO36XKgRYmYlvcGuwJp33Ymksrt0qG5GfO6qsT56tQqrAoXFLL
ONw1EOvwxkmDGrFbwvVfJT/YUSOvtM04ApTSgoypSxjYkfBuiU+EN0cnQVrE79rr
H/356fTUUMczwehO1b/WGq9ZQlV+0FOdbA05X5R0VnD5ZVKy57RdtldXROSwDhDp
jTZxLZ/Xg7fV2nFP+ACgLIqPsfk5AxftTq2hc3vlm9bHvjkbfDEVyjRAf4QaQrDE
F2i4v+f5hLCq0KCuVFKSM7Y+L5yvKwLhU68Wf55q/1tpjMO7j3DS4Tqo6RHZp+L3
6DGfCWicYHkyyy6vXTZq0iZrfiTwMw91LzUG2xR/jZn5goZ/jZyWBTEiZ6tCgxqR
VPOSVUzun6iNQEWmG+Y1rK2FQMZDAO67jW4Yc4L50uGWsFg3EfSybMc5lk2dph0L
85jB97ebqRiOKCzdgdQZkEaoSy7cKltq9ltje5EnryI2PVqirGk60YYGYmSR9+DZ
nyiVe67E7VZIF7SPgUP+jGNXkcBTcBiCjy652Ks2smc5E1D8xxgI/N25dc479uyV
CxpsSjJQ7ET1OFhBamvcGVjdPcCAB61AifeCBhEVCWZRZYpAAlzBZXKbYTOaFmO1
jM1D1ZuRt604H/EL7DPWqreD2aLKvgR0fZtaDFtBn1Rae30xkhj5hw2AEG44seLL
F4yEzNgL2k2YQU6+lfOuu9sRopCYhTT1IInJlsczxokUb7YfU108uxtq3Hqut34H
2ez5dKcGbnpicx4Do3mrrare4iNDHS2Wl1isTvJ3iuMDca/t1JzMOxJPlpJEhS/h
9lcO3sDSYglJ+m4XcKRfTMmRWnnH1QoU/RPBGQbLjk4dPGbcbqkLIfSRkRm8Az7J
o+k3Yv6kYuFKrc88CyHFtA2bD0RCn8YCOY4bqt2b8GJgK4n0bYsEvrvjErrQc7cv
4z+4QJ5N/pinYGcNVQxDYpc7fu3UZ7nI9XvXYM3vdOCsLjhNryfl6Cck3hCxesSv
JE8nBbpCfxjDO22OLEcKVomneMxePPvWdZIdLZ/hvXy9BYEh+Z76K18k3AVhW1po
hUqJCU+HRFC6SB4jyJqLyAYrqHOVqM+6p1UK/jOC9t4mvFpFbdM+dK314NMgHB9P
WntCq8cSh9h8PLC4pwX7mbGKRvwtnArkzQD3nni7DZHKvCf64oDhwpLMeS4IuEu8
rdUMvkVB/mU2tpcCp+Zu0i3UthImVkllLDxTDfEjoT5nkKfRF/RUs7neWTNQ1zGE
/MhbM8tRKzqBgjNqEnWQ+C/Lip4v/bqVlxcoMKWgJ6+qgwWZqyGtnK69jyrlFduN
6uX4PaWJGS4J/GDcq5QuN7IVpLH62qxlLzeRi/EGf5zeU5S/I82urFd34fHlVGei
Kpve1twUWMPppFagSeChJB4aBH9nkcPZIeZRRmMkrDOv7LgDdC7aipl+CsQllpCh
mEjzKvyNR0QVdPFcXo0n0ETKDaOvqaVPu8WvAHGFIvlm4D0aTu3TMdGaAilWOfIL
aRZz3ibVMSIEtYvDhhztyJPRt3QOVhglqdH72e8K0ypQeckk4qk64QdF5eTtZ47q
pCjSWL+tDGFlFzitKoi1O5XdCQw9Tzkl4dQ3T8icbgZrA6S5F1fMx//I1dCbUONW
mkxTNNRrZqCCucpip7IWKGg3xt1x91KaTPyuAvOz2Mz8I0I7Jb56sWgQCMm4JhTC
3jlW+vKj6MS8E8J0nIqM268h/5o5VYUyBh37vGwNTjSO0nxmLve/+UkQoX2nALnD
DP+e/QEz/8fX4VZAkLSAahxpFl0mAGmPo1vs3c0zj4CTvItLcRt2Ze8v6Hoz99sW
Wy53BsLfsJ2ZKJI7qSmCm/JHvnF1uWvLiGsb4AQn03EiUuhShH8TkjCuH2sU5RnB
VGs246z5yNreau7DmEgpXMTjmRNcrNfl5guji1UAzSIIntFeQFwt7OmkChz+1lJL
A4xbR+SbgEdJCICu2aKCVyLKAMVhViDwRmUfq+iRvCQyogoeSybuU68QWs2hQiu9
/Sz1mGmHwuYkYgSNGIj5eNyGnABz70vX4dKkv8YHwazQcN/KPhnG3yXZ5DVxG3ap
Ue7t7ZT/e0KoowFb/o0ZqI2lmDX9kBsvnCwfgbNFGGYQ1zkgEZr1St/B5ISdOuhg
N129OXk5qLT39zS6SJQOFDK7o03Czj9Z/W8Ci4NqYr5DKGVO7FD2s7WITD8j1GBB
4nYeaVOQzxWIBaVGqD/9JKAHAW+rD1pOmVIhd263woKboSDcLXLj+SLmOBzDsEx8
Viq8JGaiGsEUHf5ydwAQpSaRUK6TbrOf9DlHrt5HyGM3/KevHqpJoM2gwXG0CHys
cMDguFODZmanUoV9ZVdpas/FJ5BLJDjEJBYEOSmE4UqmoJtv0EfHzaVw44pgjiOA
Su86g/KQaJAz+ZcmmAVvPOiDwIlHfzxKlzu0C9df/P1MfDlFzhXKd9H7ZTzMc2Zp
KhmoCUuKLzct5ZbEndO/zNqBkxid/xRd1PnS2leUKwPDo3ddM+CUlT7h5FAIypW1
TRTvdRYXgdZHLUu3Q/ZJE868gdIA98keGD5W1uiXNUk0wmgRHLvWjCVzE+xpYreu
wHuFS07oUFUWI8sA6m60SAK7Uymxb2S8RyB+EUg53w4sz4FEb7BQFuLMo+p7MdHI
Nc/ecsETpwuFJQw8QYnwMZluAhu2iMRm7TjdQvcG+nyR+/tPFczgpxgEax6jbfAh
q/CxhGRgh+AjSc5NL/yJmnFTDnWqFEBgiVMlBOSo/EMJ3pdj1GCyBK2MDsC3yoIj
7l7+3z20g+vWwuiVcaE9mbZRL5V0RHqe50lOhCiUnV7eQd/7U/oHQDi2GonYJmah
MFlM1keDTYPZHXmpJ3ClbcGbyPri3z9j2C9SDlIv6oF8ebP91t4/bEcJIJPhsaN9
7WZqJP5LbihpC5hNuJxg/7BewSHE1aQK2+8De4nD3xDtVj9b5xXIVAkRkQEAg6ie
qQ7dM0Iq7eQo0Op45IFZVWPUbIBV5QUz+hUTU/fZeNJnuLlhCoA/IhqQJXt5efPu
GPA4423R5QjjRrKpaxG8/OZe4MTK0KmEBfAiAdVdjQq/QLDWCNAd56NSKUGYun6d
xGSBegZiwbcAuHBxstciMJQibc7hOCurAii+qP8IgihUggY41rhPN6xBHXgPYaOT
Vxw/Gmodf6j6IIMFgWUdLI8NOX69Ir3WHSUZ031PdmmOc3AkzetuQgN5/Iq7U5fJ
IwpE/UPM3ztwVi/G4TA93Vxn8cpM1IHyzjJNrpQVpkQX/IzcAwHlWP2SbOLHadmy
P4Kdk6QKSgjPl8oYHQTO1C/kCYP9hgE/blzdYtqpy68AFTlWMBKV7WluFZaD64UF
tV4CDW8IwO7xbU3x0alOXJgfjcFBUU+98Z2gT45iyGDW8LmS0vj8ljsnC7Cvny94
V+3bD0waNCMYAcM1/EVwQY8E3mOBnAdpO6NyCN0qAS/ouzcArkHKINreQ3Jd3jts
QwbtSLnAHfZ9+19yEAiHl930pFJpXdhZI5xFDFkhCp3YkbFVBkTXBlSzceXB+XTm
Prw5VKUDnodvYvi+qnli+vAijZ+6kV+0NZ7h476W3bFGwXse5Dun9OGlBWGEEFim
ncdbkI6L/fgai7lh4eawOEhE0QUgxjTM7R8s7rwHgzUQJB2xKDDykdmTYtNtaWlk
P8QP/WdLGyRfUpB1k+HcPNPH0LxbyjTfsl9Ftm12OGJhJJd7vqJicWTlzf7lHS/H
t/kD9WWaDGjL0wrGiJc/OQrz7ztChPjIbzOyy8lNwC8KEhxCKIyQCuiKZ7m4x9ij
13FonR1ea4jZOY48oPbWVOG4NRrYkcSnhl5eddvE1UkLcSrtAVlQBhM1DMmLGBlC
G1Drzn76P/KeOaYj1qlorQyRK2w4C6wb85cw8P4/w+pCv2ESqACTW3R1pFD07CD2
Jidzoy1tB5+7LsIRBGzQki5krKNSemUKmekJfQBs1hRcwYZWMEJvtYaAhspCJBTv
N1LL18K4MXKlPjME3fzpb/tXUuGMugQt8bfus2acJcaaS1+IJHdqd3oAugxqZ7YP
6Uzst5tFjve+CtM6QoV+wNTmfLPWpCmm6C/YAwgBpIjSXHSgrkWNE1UsA/J3Hi/N
XpIrJkHz0P0PkBaCtsTlf/0Yo0eBMQVE/NeVcHFzJszezP7/M+ckur73SvT9EGV5
vjDmauadhcro0/NMW4RX07tluhfsdudDedfmV4yQNWabb1f8oHjP0OV3JgXjXbia
zDlqF49OSxbC2I//BmoWV4vMRRAng18OIPxBmHS0VWTQfWXXYKAxiT73A3PVQSKw
ojQe83xx7q3Q0fYCROQQ76LzohSRiMwZb0RVrAb7DPSlib1IXPAMGsP7SM+dTy5n
z5ywCn9tWL0mMXDeOiIxhavjoe1sMB8uWX0gsQk087RvD2/2mKV+uB+1Rrs2Tm2y
qsh8NRaq9lkxNakiJ3RskCOBq6OD00sDjdS0l8n/yEJJH+F2wj7TtJOOsYbFUKne
mtDLyGUHLyUHiCyMP9X9tvNFkyDazLBcmIHGxmvhs3k1PZNIu6B7/fACh/mqjNJL
3swTm3G2EXhPGI1cgHwe1NMHGlkvNysaQ8IQ340eFtK9mYkW1YZ+hV+mzyKiSr8u
Fd3rmtttlIKehOyGRgFZ7t9DQwGPSzB43weRtfhS7gofThUe7JcyfLpanmjbEHYN
xm5kTOhf+Q7XYbKTHYm8sjlmSTfzbRVsYXJuVMFRFEY+pOj9I3X0OJj/4tFShk5A
l+x1p2LqlyIyCQd0IwGS9M50lnb3sbn5M0DSGCbdc6z16adnfzVULTuu/BYx9mqZ
v0j20VkZRXW4AUaYkJh7M7igCgV0sXHPfOhw8tepLWJzN29tn/HDdaOEjlp0QOBE
Ffq7OtwvCBRpgY0dqQZowcatREtORQ86uzwO2wpayupLjtNbfqnWdgp8xQ9UtSEP
2S0l0mn8sTwD6dT0AOHFpjH/yPJN71rEYg7eQRfOXTXW5F6f2emYbH5JGONQJ3DO
zUN2MQlos+C+vlA2WS+ZnCXBrxKGh0PRJVysMhld5CNJvuh1LJafSshPsWjImeQM
nQLqr/Ae9S1HqBBi+vvIB85RTSVqmDx4SQTJikVxPCKj9LLTHaBq6hYglfPPIsXY
Ks9XfZN7NIM9PPZxySOHvDCtzBFwMEwVDFDVW0FJu5XRyGhecsASeXRpubtQCql1
c6dR0d1zR7dJKd1MW5H+fz2X9g9reRp1BHdnoqLs0htWkopjhFmh7jqicARXrO3v
2aR/9G3q283m7j+ZGr4nv8jcZYTW80UpBL00ozmexemuIU64MjmOU9wLouZXUkmg
H33e0EmGEpOi8GWa2cTSRCnZrLT88WsPw5Tn3lJ310feg9RloTiGdH/ExpgSsRti
fk0O7OPttvPg7teXZcO0qz6RROND0BY2Y/wHU0bNYIQG0Q4aBXXSORsY9FacGEBl
6hyHkBXjlCYiB5oK5hXO1ep0mBlMDMYkEUn6Wb3c9HL6QsdmJTzwRvYRGm+pbMo7
73Lw3bU6NiL/gplJwxO740sDSgZRX7UgY962XWXyg0d5UNnVHCB0p9uQB5/1ch1h
hU6LmrOIsdgcbj9L6xSpoQhogLYCAxB12rn/RN54gkvs4g6IU3lKTf7dqzULUhPN
5fmgQOPSFn3sl9cMgA0a9oMIeHqaO3Q+29zQwaVUvkNAJSQ6BibiAghoAXtz1hBt
Ye324Q0Tq388KHFzxOR6l/QNbEvnOTfF99nyhC+JHAZNSSGoqIKjeSlhNfyD4/gL
PqXvB7VjAYaxT2PS/2xsHVw3y1cy52Vgh/cIlQFOsOvol9LsKSy1Cyee8Os5Hs0p
DlR0tha3nC3ABShzEPlfNIOzkZkSVrQoMFgcuEJkQ1ljDw6lz3XRy72MXo1x7jha
ritPL6vNoAXrkS77ONCQa45w7j3LAhJYk3+UibvnGMWH4I/3SIFPmtnlNf64rMmp
elegO+8jARN4RnJI8k63Kt23Bfpp5AROt5xkKszYa8SJd+mknIhqwvY8p10IeePk
kkIIKgof1NEGBL1fscmph4Ng1N18rO1uqc56QeIxI7E9C7Y/YYZRcHbo3IySFxQX
JiByd7BxHn1po6MrRgcNJZwc9i0/ic8R0iKwjC7E5ar43d7K2vHq0dJpu8L6MZjG
KSuzqr5fr51Jo+VSx4aG7wJcvCf2lWP3HiemDz5VZY0DuU7lBcbGsk2esYBh0Y5o
yZrf+2JU8jCaHD10zpP/ZiT3wZXssdzHD0J07Zhf4DlWmtWZMRpFikY/Q+i9CDWK
1rBJhcID+trrGA10FXxtJuDtUIaTRXu29EweDcjXrxgIFBUrTM5Ok6UJDCXnW7kg
V+YbWwYsUUhaK5YmNoWGVfuLreavqabunmx9PR3eiM/fhLE9GNo3pFpOON/j5zCF
uEKqab5SBJe3tOJL6fkxSnnKAcbnbIMuWw1kB4fnEZgqrNhMPwToRMIntWPL/tZl
k3B0UJP9snE2V8neD3XYVymSum55WWjgHWEmeFxmEGWJzk/2n/ddv3tBW30u+TEk
YUBwCvCidFaq9Kcs/PnS4zKsaKs+t/wmmAeiiZwq/xScMqkWk5PJtB7A6glDQKPO
l+MML9uhEjvCwvXilhTwjBGwQXiFEzxLbrlglGtzLd/XDPN9CYP4MIsRo5AB2Ket
lEuzjO2KfEeBy0CcvfR3/CSDWkHObBZgVkw3l8hgVznGqAUlzygMGR95Nlj1OAWY
2ZK+5T4mKGZCg/bPKlzjp/N2YdNgBAeSkrxM110zTso0r8ccazVuzi21ZHYT1VhK
mUf94Ux5MYwAqQx3x/BiFQktibf77uSIhkR3w9wxeV2e+stvmhcYqzCTFRkhXyQ0
lF20IpMWBKRLDBkJt03ZT99V5SsPSBHRukC73OcTYl8dFST6au9Pt4rKXxVQaLig
3fOyFt+//k1dOz48ssdkhMoSJ6ipuLE3cL0+2onlTPCvBgMa+IT+KXLvnX0sBDLd
teBOh+lTbVdGD9hpvnqo9qjgK8APu5tewTUNc2KJFFK6UEQAMqB/Ro4/FDudoxBC
e7G6iUqCMYNAPuAnD73eFvOWpt+5mztaxp2/kGEl1/QdPmKfcttAxAwHzYdxrjn9
0IpK7qKa/Aifrlgaiiw3sptogJseIQ1syv6o4XXY7gjfKwQwG60PrMHr6d3FMpY1
by2zkb9cH3cp3+evEtQR4N/IB1mOnst4/PVhWojF+ssDe45QcG8Ri/4cff7ffy2p
5b2T+CNOrGiTH4AyyG3NbYPkvzvmshtZq1nfgGPnnQAMD/xo3bvJZB98czNu02h7
Ct4XVZlDqfqfYJKTBhitz2Dn1586Ti67VNBwbkT9L9e9ltLY+7JikTEEcGhO7WwS
p8JYm6+Fu350AngIWcykkYKmYM9jfon8nZUaNEdiiY3mT5X3y+e4+s5u1Z/fLJH9
vKtaepagZqWh/Jd9ryxxBL83lEuJVA7O3lDZgAPOzGZFZqEA+v8fc6EePwxZC2Rt
MUEdzK/Y/RJOuQfkcDerdOWFbf1Q0ht7gj5uYh1as8v/no+BDz2SK5S1tiV208/k
RcfTamh/0NkNERRLoK0kZC+wwe5YEZLX2uTcQiOYsTsw+QDYLkRWXY6M7gIg6U1c
dbA/h8UlY9rkjX73OKyb5aiGU8vyejax8cXYfMXTJyM1IFfoafenpGRZjlHv2tZv
EGqtkffTszpRFGFnQ82A8zwWksmf8dsOSwX2hg03whwgBQaBOST7imyRKJoBS+av
lx1C0leZoZ1po8xEX6HxhjpWapcDiPAD4DN2f8FY4A5B0ImRwV6r5aHga5PcE4Kb
q47IFBoiKGMBY7jWo4oADL9OCcEJz8cahTErl9l2PN9lacljajZbJk1LMYPekGSE
yn3RXLCruk29Oxv5fpp83U5BA0Bb6EeuP6hxsyA1HJM6fiXlZ/zeDRX9Q8XU6PeQ
CYUAjggqeCaOzDIgfgMR7R3ZoXWKAjjcU2Vmj+3l37+hYBVmQ9Ny+MsoZ5zEhHnV
dmbH8vwZ0iFarc19t/oaNjIEvvIp9io01zsJYrLarlO909CZwMIOM+8eNQU7sWAi
iVEgbJ7iZsIS0gcAy3Vm+/C+y7T6c0EV4lMufjDBjzOp64thZ6bSwlXQzfFAUQdB
1AwGtOJUgxovukrZWVK78E+EEsd7pce9XBT4uQmclutqtq1PhtfT5JnNLnOcIS1q
AuaHn6QiY4QiWGzqliAUrsne4HKvF7PuK7LWKnbr7IT1XX673YQDq6ZHGenQUeFZ
LFsLKeWkT6xvDaLKAagz20NY6WOBXVNnq/lZj7f5IzH5wci3bFeuoolSym/Nw23C
tZvUn1qt0y8+TMKtHL2m0GXvqGgrCAWMMTZxpgGyqD/e0obBcJG1X6YmJth6N9z0
uVcr3zYP4Zx3ApazI4UPB6e103tXSmhC+BwP9E35KJfG/z3CPs87deYUgs4T0vAt
TOFSmrnoFjTYwWd3ikDq7yczw3HudjRFfTRvyYtl/AQLGzH7BNLXx7aj8evOb5XU
qTmIxCLEO2jvTnY30JD9lKfaxL29bKQU1iiSqNRJMl0ABlj7xxK81hfwTYXF43xY
3uEOrS+g9j29RMB/Tfe0XjSn7p70CtpWdA32VoBxHqX074uPMmOlofPCxQX3rRVc
3ASKeduB5Vh6QUL5duAPQuXkMbRWJMga1Q/idOTjHhN3dL4gvU9wEjwkEe1MuKnU
ueGtVXxvGLUPr8lc4eUaCbuB/9KgWAtE76cB/jWt8rwdm4ISqfiSgTJRH/E6Fycf
6VdkYDiWEmk8ruLpY1fG/GuHqwfMcm2CJgJH/DfsYT34LcXauylbSWJFjU490CS/
GuXXElg3OOLwbzbD+IiQ7f+gR9fVesC58j3vmUJIZww0TGtUqu8WPgD6ap7NlhTu
wmbZIlCrOAyDxmAJsvzIPvKKu6sM2dJEpR/RXYD30TmI9vUslFz/zoWIxmiwJCzW
yqAjMbrqj2KLpi6xgl5k2XJnhn/AxJXZ2oGS6dqcZhKFqN4KApOzDxl0DK+oVKth
eYN2FB+QZtJ44/GPsOE+lI/ARzmZ1/zmfYG8cQudbpdP9gyKPTjUfMwWjDGWwEEx
ezPaVCP2UVIOuoU9l1f7VGwS6dSCaqzPNbDEmT/LSve5gmmAI3ew2jKAcmj7Z093
qNejqKksDj8MHaDpRn8uHtsDwppA8jOWPWM5iblOmdvZ8WaBY8adU5oZ1AhcE6TT
Pr181NMl61xfyl0I2VX3EoSQdxFsGhI96DXPuARo+mIdRXXQNabgUv0Km1HxZaMC
JEAy18jzjmgC8RwGO0zeylRQFbDoxw7TikOFxzm2b/KZRCJKdzCnZIMmQ8b8eYom
1IOlaAY4GiWW+PcUqoDiMGf3xyxHo46DdeP8jsdxmeV/EYeEZZNjOYjL0PK9nsjI
Qxp5q5ApQEIOHInz3xGzCNVJ9IbvdJVL9qEhQtznuWQBxGUxIz9Knz7CHQwJA5s+
Wxc1Adp61B3bXOVvhpuQyMG0vxMQp79cr8wReNmzv3rBaJbDm24cc2V7ZC8LKr6g
VgLn31LtrtsN+sVcl6qDRbsOsJZMCQvaFz2s5Wd9QYZ7tlFDScRiVttWlZjTBkaw
aEl/+obf0dOF0ZiqRs/XRkYTCvEZjzipb4RRrWOWSjv1xkA6CeaOUCxYS3i/ADcZ
uje2QKj/Bjp0O3U11T+eOoK31TLYiGeX2rzczJluJX+noV+8C2A8Dpjpq0pwHwfM
M6nc2CIXSSrQ1QdsYn7wgYOZ3pLjRlCJKar2BkdCfGZfWoQ/Db9WJVohDjLMW2SR
HPRjmvvFY70aiI92fOsYLhG6tSNlWuTe1oVW7wTUlr1Gb7Cxpwidh9dmufmswKX4
pFOe+tAFVqZCBcfCgYJ6x48WLx4U6UdX+1xEC0TFfkJpWeaNlOCLCsr7GRBB5GA1
Hlinrfk3xDc57CK5OuWYnuF+IUKGH1+vN2cmNFA+h0YnBEoLSN6Thzb9VMWp0+o8
A7mHExGrLqCC/15zb1yUDz5cPQIqGSrDHNhcwgbliM92jM7ZTujmr4xl3RxdGjj5
+JInKf4+ZT4Oh2lNr0GrLaJ9dJ+0zhMIfq/maojLFP7ovWl7wHBQDhNdpKvMb/vQ
vbwifJygiwADwKq7TsSM2fvr+z/Qm8W18vGsjJCZit093F70iaIecj+gYCFZ48eG
xFRM+abVVfxJtWFEKqwZB2gvr5tM6oFJrqGoKddspJ14RHFQ5hOso/TmPjv+WUDn
omuIorec1OuLDB9XsZb0fEdkh0mfJPVolPq1LcUoS6C9Hou9K+h6Efi6/Yvl5whQ
dUd+4oxzemU5Y66fTAZr7LgoFfqCgmyeATxeFX+Fjx3LI2RR3wmkvPZPrENSiYnJ
v9GQK2Lr+BAuX50L2VyVUX1WgnxukkcB6TEJREnfH2qlpPI5/iJ/NopGOS+RjgmB
WVYmQe2iQLSViOhxDvNwoop8DRbDh1h7hN9jpV6z+u7d3krsCFK8ZB1yejRXi8Hb
xXrqkwMWj6p2uizi+1bO1IHyaXafWdtqnyuB/SK9aIscxhe4XLT5++Opd0HzWOoI
JGyuXGjr1qyYisQmUJVxJaTH2u+pODnoeCLWwPPGg3fgxylLX7D6zSL+NTTHVZUS
9QmCblrCw+wuPs28pU79pqIiMZnfhB75o0ucUtBgaLkVuuIAQr1DgfyFePAG+xHu
VKCod74+YdwYDzmYIR6d8NBQwbBSwJU/g9PpnF5HeUlAzmD4UdKy8fn7iLqpoyuP
v5omW9Wi6j2JuucmtBl6c4Pik8bAWlR8QddTkhfkw3magyxL6mSNI00AZqYxUxsb
/h97SoY06EiUnLyTN8XJBi3GJY65O+Iax1y4aDvwBhOJ48vz/nwQJJNFWDeDBgeM
Si49A4Rh8U3PWxOHQlt/fbFLlDtpK6rx+1B04zpnL9c4ZyOWNdY6prw1/ci2Y9pM
m9rBt8ktnKPLetyvYG0YA5Qvr7hjn7sEGPANo1zEaAaU1Zu64qM3mxDOXrTinpbP
F2ZqdR1fZ0EX/W55PVqAFku3nh92I3EItr7X8ZQQG5PR3Ik/qR79MEyIu1hFmXtX
fuBK01rDf3lsX5rPmmMGbZ9wQ6kLCcC4BkDK86D/o28oanJ255a3zUv61wdBVs2h
bchVv4RmoP4b86HfIL81hBelHQxbGvnBb1nNB/mzE+oPX6pONXGSMqopLdebuhRE
O46RaNoXhOuGh2XLCnfovqO7GS6AM3PQasqHu98xg23o9TT1TjudypS8eLMIlJP8
uLWU6ViSyfrTL63OuWgay5gEXFaWXjw+feH0p4fDw5bedrkL8z855lHMvfKHJ/ls
gsTMo2hGZW3GRw6I3vsF+wmksYCLdyBEsM/sh0TKJZ7ZqtwdNqCC4xa45HZ1iIcj
3N1BnwOBCJwey/G3Z3jb5d0118aDQVq+VOYO+vVM+46S5bA8eHNX2WhGGHG7Re5Q
pYx7NffMHfVL3QO1hEiK5SRzDMDFyMPPFrFINmXusBp4G1SdT7O1eyl+bYG60lTy
y4+G8pEQJLWL8nuo5WeHltTcKEEaJhI/zcHU2SMRfYjGqzgjjrSaV5L8JuFQ3mZp
fdM/8oxm+3MnEwINZWFjxCU/qGtIalK4DwGT7muxPzPqKrOzrF7BQzpa3wdh0yOH
FDkPfxcMRRB18gFMS8qUQwofulnwCzkKBORa8bCZc5VLAurikidnVJLY2WS9XjUN
gFUxCkWEy0kzDYIPS1jloyLEGLVVO6OwJCA+I+AY564eBtYfQpvQ4b2We3UAeHvQ
hdDD3+zP7RjDfbAfu3NdvVL/Ymly9vAPE4ms6oQanIDltKf1//+I79e3z58LeKuA
qSdzHbwIWLWn6n8127G0L54AmvrL6/ZppMztRbuLEuEFnGwnm6HLvDNiYE9MJqvy
xb+z7HvTzsssBEbNDlWnokIEzvoeQBZHdlUCSM8pLjRnho1Rzq5XpgM6C8RZTTgH
Tk+ZhEL/2b1hsv4Qq4/5ZUU5U1hGRmO7mTn24/zW/5UlmPc9tx6AfqYU/i3BFv/W
Ve3pdnh5kdQ3kensZinrqVeKNZHg5km2k5ipLTFAm6G5bMqGLoSKw9Z1ucMErt+C
FyYYz9GwbMqHaP13k6GKlhjlfkuJiyMd504DFbgXBgxBEU+4Tx6VAYKdvVzwnUNo
57mYWSGa9YADC2XH6Pdjqg9uO0erNJVRliDMeS26sZD67QO4nBrL/A7Lz6ZvLlnY
LOWuGweHDjQW+w5eCVpexrwJrPFYT2f3f1xZqArJsPJL6kh/M/uYZPFl1S9iPU/9
kGByEtyDd93X5kEudKiZpnNwZsQtOBuTtIuotck6oFRdYJnjW5/kC8r02GTuaTDO
8nZ1vOyKMzs/muxHAU+1omda+XgZOgpz+PEEJ3uzrYHacWB8Qs6a3upSp3v7OA+i
mneNRn5ztCsO9P9uoTKa9VnLghOyP4pklCfClMlJ5uFepKN2vQq9++OJ9n5xCyZT
7fj6q44TwVEQ1IYr6IdilyaynFWsMZhRg8mSxo7Vmv0xBDix9ST+6s3vGwXZwfLB
uvEI6VFE7L+K4Su6kjBTWAOdB4/depXAbV1XiXpXZVeZ3G2U3mjPE3Hv5UHQA3ra
lHq6pW+6pbXqNdwC/LgIiyryAitxjKppMZa9/Y0UnQo6AjB1F8vrXX2YMZ4MwHLY
zXvqkaHtOG9MobbUwSy9cvEbNEW8ocTHwqy6ECitOBwJ2FiKNR6ZB+ST4CHsmTl8
9eKuh7REDIVytG6FsoeE8rS8kG26RYI1DFQixR2MahmZxkyiDFa9fQVhF7pu259U
liw4sJQRaPbF2izTHYshHkqHO7zLRFbKzaXAKEvIngQwIroJmQplCevZLNcOitMH
w6YbLaUxXXdrEKcILpSkXaSSvfA2G9tfawz+Ec1oy9ycDw1wn2wVJDJD5crwayMG
gN+yaPfeCw0A0QkZ8+vReYO5RbmKZkFoQs17Jh9WqhSZe6e+DKccdI7LaWclE7K6
HQP82vURsqqYODfF8zz4mrFTNyLMzVxVTgOuH6lVBz8gvA0RehpH0jUPZP0BSFMs
MZSH5k/p5aKHJVHC1m1i1rxzAzPQ5s09HeiWsB23aWI7doYEIg+qpdf/CoB7ORV+
boFIEYwFpLqGaBmuAcvMngAPV36fgaPs7cg1yYgyHInNBxzREr3uAeXUsyKUmZNZ
n+nuwxyM44mAUmAScDfYuTjHRdgBD5ebNTKnC4sh/yiV89mLjb2xEynrWyT2U51O
S/Rgfa13qNe/61g8Hq2692isFVdtniyUkz9Thsmn0nqLox+tNRmifU4dbfKVS1Tt
oQFcQqwhVx2EJMl/sT/qpfD3UcUlU3q6mbAanSkphF0VDZDro68mYtap7wXqiHEG
Jw7utXMjW1RozZmuEQkv6ciMfdG5oLeyUI6kOSxnNWbaBGlnmWQG86smYzql4Xer
jNbF1ZY6Am8p48etQm4ueh+A8Xb8UPAB8cBkfJ9x7/UXUdVtfhv3YdI9Q+Xez9i5
HGekB9SxJ5NNxLFphiUmElgWOSoA/38SVLCBYIFDsdq/1wjJo2TX2Coulj331rRX
pQoM2zgMj9To6YAPgdIIhoYBQAf9PYrVbLfn662oLiNoYfleFx8Uz6wLdzrGbhMK
6rTWo0cwTwilk9Oijjua81zxoonfZS1XdeO09RhU6kPUIe71ikR8m6EfZnezBJz0
4eYU+TPfrtWAQ6VbmWvkXJhSm7IUReR6ByZFd5aSKPoYg+aH3eQW5MjnqrOQ/Tlj
0Gt5n2uFpMG4vasV+TT3lkSjow2uiw+7BCnVsLTaGBgzwFnKCgzapqNvQfgnwRZ2
ck/c7TfJFLOhZOa/QmiNZ2vQl40IGX0ggK9vt2T0yqRL0Y3dFhuVsGArvLZuOR+j
2lcwS/Z+m6SGODpYiuU3nOHGPHESB6gOhtE+p3vqfzIqdbDTvLyJ7tkv/ZGsV5Hr
s+plDXhuAtWLLuR/bkRHUqkGdmzrMP1/NHlpOHpQJ3ssD5ON0WH5zF9XOfsH2CZC
0lxusYYTnbdzIFQw3PKDcG26pCdwfwJ9+7xfeyU/vixWfgjpjxxfAj1+tWxAAhEU
/taeI9NVyKnxIbajngIHRokXAd5uptGDbHT7KG1WAnk3F9x8ifYm/xabQD5KEURb
YaY972Xa6i4qo2L5OfkWUCR/RB0Ay2qAAQBiXbM6lU9d8sautcGw4+iS825uP+2s
bmdOye981/AiMVeAMsug8314Dy9tWz+tTAl4lwyWopkK0O/ATplmZshWNZcXkuq8
bvgGfMCWG65h1sA16AX2wOO0lMCFlEZUvNOFRYQnm84JvJvt8KGeZzOpc4mu2h1T
x3k0uqzEOJJD2QV6EHnwvXNQtSMyDbuKt+MdrXtJ5ly5sJKV9E7lc7s4kgjBaXa/
3xnGxD8694EBY4Joc4gvNiTXENMOeDUVajRlhNt1GOz0ks7ut3hyn7QxlVz16NVC
zRD+O6Y3hRojljU7644AEPOKAgKSf0E9uSgbdKOn0UINRA79THHxZPRWY5bArghO
0LBnMvj78tlObx615BzJUI9IxDmduXJ4FzparMUCPeohtUxLWtYIcQ4gUONWg4CU
pN7J9YvANyfoZqGCk0D88B11pTHN7hNv1GyPH0ugOY8XAc9WSuBKyANIRqwN7pip
WsJT7V6BYjotx38NDqyjsYJByU1cqd/vHkD1KrsCvwRCyv5EOgSfaC0XhMSSnHFH
JRyisXhnSPk1/AToQug9HTX0gzSXflLMvDIs+5IJHuH8plMstH61azbpn9IaO64E
0oSLMY7RrWHamE8cP4du34B2JvL7q5ear4MlMjnBPQwHvn87nB9nw2zvzxteZtxZ
SSCNCgsBGq3NHkpiOWqqtXS04RrZ2FtLBKwtx530W+TBubMEKhRRLm8tOkqvVrv6
cjYeX+9QmDQMoUDOD8pC0HjAn+flp0zoVJ1ECDSlk3MRKxVyLSr7tEea7HrZnfM+
Lq+qHSE0GqW1WvI2qUL2fFf8uZaT2d4tVNw3NdPY5oX1JiILg1jxPpB8JqVe8vDK
4Pa91ODH9x6lSdWU41qdQirV0GuGiZkQodUhvQHfRrkBJJAsEksN29kFrPpcFPJi
c450UHoeNk6+W+bAsxWnRQ2Uu1wlW+WzsmWjyn5dv97TaQATZb0c0j/ryNwV70i+
5KP6r9FO34PHnwkJR9YT2PNv+066wO27ON1DfVFcAW5s7VXO7vdA3daMoNnBgQQc
XTy/h87+IlIfHiLn4Wqe21pMrShGgTG/k1umLyOaAd+jPr317mgES34ST9t1WG9T
ZNOkEHoCakEK93mTIn1uovJgXtmP+VAW8gMFg9LhJREZKo5j+0TCB8f/SnwD3bxy
+fe5wfT3Rrc/MJV+WoQQm7I+gFeyjz5vgN7Doq5ZBkg2uycgQBE0njPIOPw79Hhy
LQfzr6jNAKKOjtO7A7eEgLnYxWX71gjQTZ+8upTXQRPC++U/sy1z0cWhN8IiPR1g
g3LZ+DHZHZ6TQNp8c6iZS9Kn4Qmth/WpXjxxsJIXOUTghfQZblAnjA5ZJ3yn9HeW
qISyndmF+Y1Mc0I41gKxGkIzEprlpky2AB4pn83xt+fozq7KQUChyKZcD7tvlusz
W9tNWTWWzFSWkvlzIqfJqsVhm5fTBF2s1HxYrLSmE/Vul0n0wwtVDRqnk3hl/ilC
SqdyA1ymaXH4F13GTg+J9WkTlHzzAsWh8QT4I8Cbwj7J4h/4rjo8uo+3m6NqkA6Y
Jn4kOE8lMJdX6W10lbQXBdOnCo094V4NTm2IQOJcW8AZzl8N55a/YXEUUhdDGhye
FMJHEEbJ2dAdphkuOtQigu14krTNgvv2V+34UpyTswaoMorqvIFdzyND15H7uTG4
ef3CePWdJ1UWMIH/MMZ/wdz375m8eZ07kkXEJRd8WJRVecfA/P0oKePh10DZ0BOt
LT3kwEvtgZ8ga7vx1GbtGRrvZiqfox0+k/cd7TxuK0LxNStY+8iP6ulvi07ClbSK
yEuWLDJG2O6c1ULA+bZ6s2hgSyCNjeCoAgqDDpryXmaDXDnx+5qNibhUDXhCVSZB
RseQZ2JAyFmiwYe9AhGfpU2Vq/t4xVxOZD1iiRqLwvMA2NbgmZxZqwQSdC1b/VtI
l2SsMp8QFIusRBS04LAcNkIx42v1EoWs/7ecPRB71u/rsRZFeFIF9svAD7chmkFK
xVltqtmmrJ1hV2B0y4yW0vBwze8Q0bmhZhNxEc3fPL5p0BgevoXDDdry5WMjwxUi
czRBih5lVROSUOKKrK2hreUBIzQ8pdJLggN9YyNUWBms9Jge0lBOEs84x/UZpnlH
7RKnUzvk52UN3yC9BIaP7RD5uNQYV2noZ37hSC8WRzcrPhucMT3PBzfZUdVaPg4K
IJ/HBTT6Q5IZk7Ga3wtovilUlTawgoErO9QEaw7Blm5E/R4L9/h+BjaqG2DlieAn
hcvMaH+VIuybip+z7bdKVUJwATnwr71LLrzsedAn+4SR6REYUeWVKTOx1M4lffnN
PHrVyHKnn9RDR1w8hnH67X/do5zNK6zfy5QArrgV0rK0McprKY3k/QtaBiiQtVi6
hJsiEVUsPFuKnMgg7ywkRAhmtpR77regaZGFojwC16xf5EQfCgsajAxtwAH8Obpv
6C88mPu5Bc9H2WStlXCDo3PqZw5iGvxComwK8OdMF5xO1z5NKVRF5XkP5hdMePCS
SR/ZuvkTyw6/cftqWGuvLc40vopxNFrO0J6vOSlqo/G+2xdahoGYvX8RH37bY+lW
DNjAjhkK/ZcoUixcN0dtc6Xi/IIBa3NmSB+QeUERADnvubNNvncVMIMxMtnUM62m
7Gd2UGc/XDERZ+k7cM/I8MD75WEmwNTZFztiTFCHjaE7SL852KDSOyh95xlWnJaq
zebitMA3aWm7N5jzjgTyIgiWLN6W26yHGsyq1fmr5j3OVsecOHQQNjfNkNuzWz6s
apstwVRsqKGY5QmkepCquB7jopqE2Rc8RfVd4tJqzUGVXeqziYZmirb1vHD7ow2h
FY2KO2mXYjK9KqBDBgk3xfRztY3yOAEttcTeqwn56H34ZRNIsFs8jxp3dBODepui
bHMbJC8zcUVhmT+DaVF+HghRunztFdUF53ZRkiKbcZaSUYbk7S8gGl2erw2hr/Y9
VE+h5RYgwAZy0nX04DmThFJI9q+erpm0eDdmo9r1+iR0OclqIFdi4r8+RiiEzN/c
ieu1WHWv+e1LD+N+64Dc288IeBhEew0PQZvQ0Sni2L4Zv2DEBxTRvXcYsPJsJiJj
gfghZYd5qo+/KePInWkp4SWH5CsTLgMRtpmbk1vjzOr6z0YK4YGWgmCLCGbQRHtb
VxmOXts1wWt4uA3bxswR3QVCp2zM7RlKL2fErBgri6RmGexbG9NMIk77psOM9XAJ
7eSZrsNOHWZEVJ8gBwjzGrmRwBrT9ZqPBrCbpCoAc4POXBK0hd1Tzo4Zl99zyp7I
og0roCQtKOlQujOtcZmptygFW1+fIh6ROZ+jVWpFfAzOrIHivn43pdw6+mCWTO1i
HmZ6Kwr6Qi2JKm3Uel5G0zmYPWP4cZjB71A43bak8wcPIfVamxDnSvKi1XtXJHe9
XTIpD82pfhpO5U9AiPOaXHqNO1PM1L4ToujLRRb1Qz4b20DEdbd4cv4L2pbOy916
4TM4Kb1SKmDqQUpTxSFyvMaD9R92hhfoJi3Dipr8sbaJQDHUFZmcFG5j89XGqowR
hzRoMfmYCfgcqjhCsnG6EV55OjF2ADjsHz3ca+ClPnU8uQOpREkq/9gOEOScmwO8
brOxbZjYbEUUhTse85yergRCAraqiAFYyfK6+EznQOkoB4Ugavwvs3pMzyFcsm6y
74vjewBOC6sTJ9crrGec65IXvH2aKmAN4vcQhPaW2sdeB8ZGuZ65Slhwr+NSCSDu
dgUlMmK1TEIuJON5OQYvJEouJDzDg1y6hsoH2vpr8tza2Z3qkS3Z8a+j9MjZRywt
eop5zqLv8m/vkcecfsYs8n6t8TrLSmnLnT+tyNXOlUhHImN/Q9dBOzFhHFPRtecf
KQKEQAtqnggmz1PU1s29ef0XPazGpnngPIZ7zFNWjWY0Xfvb5F9ZHTh17GZkftG/
iKpa0RO/dftq+IhxLo1YQBrrkHqCkn6eqtarHWsM7VLEy4jaEK2hxO9rJpS6/QvP
G3YHG1Ihf7Wbfrjo8gFQO0XvhKCiVXhBsgHNiW6GMcV1veGCMkbbojHacnvTmj8/
x/ZEYeih1ANTuEah9Slrj1d/27Fil9i211kTpLPe2zK19dpmopvw2JGCTfqA9CNA
TY/LrKBBed7+7g3L1smhrit08NuwcU0Pwn7l43kwXCrs5d7N140eHbZI1Pw6cuQ6
eOQXD3D8c5qSCX5Dc+my+TC0e2hbo4HuNt54Jf/v0sI/wZX+dDIgLbwRhW9jnW4i
Ewb7cEDDSiTMDko1TsPsDAASsH3Fl9bWyDyLK1gvjba4PSf2t1WPpS+YhQErXafy
yKww4/5hgjnkjYEGg3yoKY/xLwr5AikF6T9hz8CMN5mbejaXlRwKhmgteRaSRZPa
oPMJVWa5kGwxJAVgFX51CcO0Chf7+vTJyuiXmCACICj8/mQuyrqzdwxRVvSLdU85
/DuLUlAAtZph/e6/bJ8mpvotYxZPpVVzXxyuLkLo2AovEyn0Nzs3VtogbdNC3Nu/
P0Vg9lgKLcDrsjf5pMS8WKvFzAaCUTjGVZ1vNQVJXqMPWNbNCGrtcm1RxteQhHUF
LtPbhf5ATSSg/y+NzTj2VpqmwHtVqXF7R5gQv9qWxg0tDLjZ8uJko+15b+22Ep8N
vo6FkY4j87NA8irxpy8anvt47I0RmfjG0aHsYlIzWHXIHzpyL3b/lf4WZLg2IVLH
01LI/azCaqS7eJ38fNbmgMv7LD9aVGMRLB5xs/qnyZiY+J2EIIXZ2QLKnNkqcd3N
Gez03Mia8BQMHwpn8w8KmhBVHxUQetHLBVu/NgRUEUcymfhgtUqIlTqRX//ql4D0
TCJh7Pj597lPjmH4J9vEh7r4PwaFoKSQ9rEWRPHlxo0mAbErSy96/F6DGAs7UwW4
ae9diY9tN6kkS8KjeR+lThJsB4ICa43cpGb/+WLctX8zWkGqV0jZ/Oj1Ma4BJ+4M
E+IOYdsVyjOWDS05qOLCz0XVClTJ/TjLdl8ZwYzPPHQkvroTfCfzEoonANeiAVXT
0k+AB9yGKBMRslgno41diLQhMgwient94i/Q9Apw1mMZhbTeQXV73X7wRDnRH9Nw
5lv5Hm8P4IKzL5yPTWaAFpfsFXv4fxQlLttAZ6nalqUUgLGEkdlijK+IOfL4IRIN
UNp3ksOmGfMvnb1kpp2lYBuX2fSQZ2Xt8oNCuZzHqxr83b9Zo+H543p7arR58eRx
JHdGr2zNOLGjjHDim4KpXiu8s1WStWrT21j/WfrpKaAFvBdbLitxx9qtg/hIDtF3
xCDtdMBjX/MjT6imlc8VUKHwRa5bnc2Bm/FjSrhKw97lAUyVQHp07K94y0Fl0m3P
cJXhJKgToqNwcBEZvQxQsaax1c5o6ZRxNj7MfumeDAu07lvWgL1rxJQgzwQcbEjd
`pragma protect end_protected

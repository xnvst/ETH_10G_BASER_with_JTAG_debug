// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
JWw2TrLtI0Oqj2PEASyHZ50C5ucm3ydqO5F9ChIVL2YHPvR63lCTho0+fW1sw1Pw1bbHDIDxyHDJ
xBWm8wBPZPpCp+wixmepgqH3yzzqgs8JmiQzlb3OTEZL+u2/eBB9VCMF1Q5iWhBcfKpaTOMQyfwT
Zbm+8L57LxayiO6AQ2lRmXEFjUrQJ1MkD1sIrIdi+6n2Bu51fDbbIcNu9PJNUFvzd5WMXxOc8Vli
35Vti360rEwFFxwYfnl8sBvfrGITgTW4UlJ16GjP8LtHBQbjnBn+0QxbP0/AZSR8+aBVailcu2b9
h0Arfm7jjilQHNOaWjazenScmBE0xbB5PvduvA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
wUnQQK4cDm0AB4+Ssn51+ddCj3iMu+VoCyCw4jS1r+fbUCOtn0eIUZ8Mcx7+QuE25kzHfxd+ftHI
EhFkX6jiTXfFiPBu151EeWKV+8b+AmKBE4wkQ3FRvuL93HTlRoIgmh5tsInzYAAT0fIQRrYspQ1u
Qk1SEPSRmGo7BfbKfLosEKSD8by+4TNK/jS0BB98DJebqfzUTZ+x42EFVuIzv6qkeiNxA98I/MOO
MHfe5e4XjCLzGW4Ml38yo5/ZuvVq9E8FgKirN/C/t1GbRS4/egEejVzJEXA4rP8eBWS5sZIo5L5o
Ii7LLjzmVcPy+v2n9EzOA/RmpMqFvwNY5HgfzX++9QW+TZb9uTCnmPnSAaPHCXGOijj9fE36kh5w
+hNl2T4g2s7rO8fs9SJDVkO+oBWNQ3r9FNsOR6vnBxaqylLpaMD3Rc5YJksWdQXf4Velz5Jlp0aA
kxgCxt9ywxenhgfwJ/GYsDKLGAhBkqMQX2JL18A63F0mIxYCaNQC9h4tOSI1raiXypt7H8WJFJ1w
Jb/WPkcLpXi3HOeXBljCQsSrMa24Dgvrb+WccnfXrSBw0JBigkkszp7BI4mbCFpmBCqperVrE61r
qKep762OZbP9b5IACAd8LIbvqNMdmp+PuFwhMNey99KbX2yspp9ik2FB97xG8glmXXS1WAPxjgHP
qxnMHvNO2IUl9oC7B/yNSREl6E2PYdM1noLNJnit0hUbmRoWUo37lis64DqeGlhPLDIWR4A1oLRj
YUwYQFE2m9yHD9DSas12ZYsYjI1vORfcjGqzKheNdt74By9fK7Y660To8N7l+9uociKDsOKvlubp
m9L7DSClHd9YCPYbXQkX5UxUuvfkFxxFkFxCGRzh1Dr+NUHIm96ce1sKS8IF2g7THFHQqmjTiNwK
v3jQkamebxdfpOLtc31uLFhJdiBGhGTgqjUpSOSOQhiDbkVl6n5U4jIpnZtZ92VAtwAWPG/YX0Ya
IL/A8eabrR31ADhaX8p+PEiVk/6xfw2TxBKy/ONOPLCgtaJYEf7tT9VVfhA54bs5254wmFDvpJrU
5FLuNjx2/yj5PQQDuuBiLWXWi4xr9X1UgWZehlIPGDhTyu9VEi8AfjEG9O4NKAR+g62Lpw9sBtey
djCjGiMKedHLg72GuFsG5dynMfY1+EX4eHGcqbPcmY6AyLPoVMMgJUeCtRhgmHdZLPN+rbwvjEzM
hj50KTAGM7Fb3aZtKW4VNziGGObgKKw7JoQKXWA7ryJPw+8mZEdxXcS0R3OaaJ63TQ34lN54+2qk
jpV532Ql5HE6PWR3xk3OBNbZhvw0LOUKR6mW6Al/UjC0dfFUfnf3pidiAtxdIJLqxv5quj190a6z
yAy44HNR4PZL7nF19negR6isJz9CguXEqm0RHELNnVXmvzB7NeXonkOpssNPzwbT4ZSLRcyCYAXi
JVxGL/IAlrdz2U/SnpwJG/99MrzUe+jG7OUbNn6xPA13g1btgeRYUVzrsO8tTw1WyzaKVz7N9ll/
O8YrQxFeb1l+XrFdrHKogAwKndxT/zerAIlpLH4OmkocZgVo4jXYHW4pwmAMXJEvUoxPzOuHGRbg
i0U6lBJN+qOaEqAUn6oAn2Atvw16fHjwGNkC1zFvgLyesGK780NXIUwEWy0ZaUSc4F8V9tWDQqlW
tLq4ReW+ECQJESL41luEl7oP9NCqeOHQIUhMVIbir/kS0358v5zIIvWmuLmx8LkDO1zhh3eY822e
93EZjGjtsszgtxw+1HTUbtBSDi64SiAbTr7Ld1dL9iIz7wti7iSidWxC88ybxThw5WB3oX+TAVag
GQOZV0SIH1yM75RQ0Jyo2EMnDOCNyRAm3ZA415HOsIDhVU9rTuutd1lsaqtzDt7jS+KIRBjIcSf9
+YLWQ9KVrD7lYRIjMQmByy1ZTZA18U8JvBlXtsYyULkebh5AQjQPYlP8PLxA5FACzDyTvEI5jpVJ
nJ9SdIJ3pRCgxHNyKerll6g0gghkGXy3zg9LrMpKGixQ+uvRVhY5GVC81Azz4jU8HNfxjdHc0Ju0
/u07VWcQZoVLUlN5tm2giQrXYKX4I+LUJ1TwhktpWox+cs4C1a7wO6d97zJwoz/gLlVjWfS5pxta
eChL0hmCiiffOYUnGEuJTs4W3KRNejrBFVkx/OkrZLhR0ioV6gsE/Zz9VRbffLbg8XFFj6nj2oCL
keza5XDL7HFwv8CW8Iz2ZQcXr655c81CsNVevDuMB464fTyGZ4yPzrunsZQhubdFlrVH5kH2TbQ+
vBnuUCdQ9w509RiZwaVl9+1VhEZ1KyQef2KJrYKz7Z7K/GL+GfbW+tkngTIA7op/kiN+H/QjckCU
jwuLmZ9ewRY0Id0DHPlsFf1+k0hOzo9PMx81vuSiDqvwYtVYC/rGuarmzax1yF9xokiTkKnVKrIb
zWhViWYLytYn5FiuzIBj4GCyVgOMnmFUnsNi28YEYNw1XG+u8Bo5Be4nJwcz0arT8aoh2ngDy4Jb
KfMNV2lq24A2jNZIGlc1Oi6Zq9Ec+jmaQy7jKHHjayRba+ZlcxRkfqJaK3tMS5e5DPqjFU4hC66C
kP+TY0vR0B8yXH0jjU92/eZT+N7CUdW3szdZmXkqM7RbLrUUc4SXq26e1UUG2HKQmA/G8q7cPV4p
/W33yZZAxt/7eQNNnY8hTyHPycnNTrARNNYvVizqGhbSFk3izXnRO5/SdAh0YFi95D7SLnIfW1re
0jpSYatGSSDm6YlDEZORq24SP40qm7LXiTiS4abTUbVwXI7Z1LbS4woVeYknh53mwH79cBkZ2B1k
EGnizUkBzPwtByvzHvqqAw4HcZToIVI9H/X2J0SvQCGA/A8mu66nd50j96vGPLxPnT6eeMSP8KPv
vRt8dAo68blJJhDh2yBFSwMhXLC2vOHmnyg7T+tbTa4KYnMX5dCdQAqyeLuvPkq9O53HpKlPFJjQ
jSyPcOn0xcrbb60YfVS8Lee1udDDC6GmHMIF9WBPo2LrKJ3baHlXXmzYxwkCq+7KGi6sFd+nluRY
/5zMVuZ6ttqfGuvb/MqcMGXFApJK2R9DxyGO0dn+hZ/sX3PAslAtlZbxPyPNNyktQFYMHindRHdf
DvFUES5vQAhLL4mOxlnxHf/CMyZJH1NFtYNfF1yKIWTcpylycCevUPb8QnzLX14kZuIdYVqMOR6e
SUCYhy4hH9zaXUsIp9hGserKj7O9Fkq4DLPxRfPu8C/Ka1nBfB7MlAPjSose/9RywBqiHHoWs7RK
Op7ksswSXWZZZfWPlfzM6Z4meBBkke/3swJZcmiuQ3HMB213mOh+VMcpoM2ciUT5mQRiz76zQR4u
tajL8dpEY6hznSS3JUBEPFTIUfV61E+40NEGJcnXU3/2Euj8TOZ5r8PjjswFRX+ONNDgPUiFm4ag
M14f59USKWLCXf9BQeQ+h63qirBETuz/hLym9oryhKi2djrpqpyxsAO+c23oavGSlcI9sZN9M06B
JnNbQy5QhzoneQMOWXiPQUnogQ3vsxUIP2U+OBj9E3JU7JglaGPVXgYn0wZfVGfd8K8V4JtMH+Wt
dNjlG5wk4ge1p9ELiUZ3lBdfW3U2eO7Q4tfeFEdOUNoehdWNSknjEQIBLHB9wP5N71Nsex3OgUe/
TCyUE0A5DkhZGiyWXfAI2BFZ++ukHg+Y0aCL3LKUUG13MPwJM3aS4ei+qp19a2iC6IA0Fbia/ts6
2jtp0c8ZJwEmyLG0PsH909Mcb8+iiyBEHGhAzUgdkSJpA9BBBRhWDsJAbEMjWljxIad2LhpT3IFi
rAGRll31mVW0TXQ6DRfZrFRudNN4Ucy9btBwIVwlByWak6D7/+FmH+b5uLiqAKYPzXaee0wwU3Bh
S2ZtVSBCiHGKmUgVqhFiUFeD3pf8sPNNzbPGWAchh40424crfEMbch3p9tv+J+eUyYFdIQOOkBiX
hvHOMJFdCYV3VSQ//Tb/K76OTf/u9gdIgA6ZkKGL6ByUI/R6x1EfN5lLmEbl8/fAdZlzFkAs8nSs
CLLtetaT5qnLUwltlsD6g26CTv/FR5TpI7oMzUt1vihQjAvZRiB2gClX1J71hWZGdF1FqglyHiXB
GIaqP9elMHINauPs+a3auxfpeeGBGVOvfHC/qgCZYFfvA2bcYhQ47yyE7vg9BzBq31Aj6kWFXDj5
YNmoetbbUKbvSx4TpzkODtTlz/qWRYF88ySS3rB3dh+qEOs9uq69e7VlT+CpKIHhoWHFTsivAXpw
SM+vEZqqnL6lqhpVL/eKO67ER2aR8v/TElRaz6a4l9HmdCMgHW00KC6YvXaafh92bFnKEEQgmf0e
7AqNvd0SrkykDD7Mly+xAU515nSerxiGOHiOEOf7dMUkW8Jei4wCqJ7UBWsR9KaOe2mZ8Jj0NR9g
yNdFHoaad/5M9NIJ/xLdhcpBLl9QACETOBOERsS/h/pPArorGQEkMVSit0zvDLV7JcX9MuRa5WtY
fMW2j/BI05ol92as9VNMJQpfTC9uJz/x7DM+dqZ+XJrYpK02hzZV/61w/kcDyLpUjdo5vOHKnoSl
FvqzODLcfop8yl7gwaKXmZmk6maFxOVfXlDIc1JG+HX58XnbHGCRpEwRNqAJYYNS09HESB8k+Txb
G7tE+9+Dm8IcWN8FpOfAB1XhxqYBykeLVUzXoYMAY6PD1ao19uq0/z1JWvwmkleqeuXMmgsUL++p
GqubD87MQsiU6XI1pq4bk+UCIKNWWs9cxomh+fgCa8Ih0jzvTbWlQzs3cVP6segb5bXtGYGNYqFx
hnv1DKSqwdhE4WHmFNhLDzm+bcevxj+ck8ybt8jcJMlH6jw4R0MYvjO3Q/eAgfrjtgK+CNX8nY7a
+odxBLbk1MbgIK4RSIRY1khoKl1Wu4kLJAZoTdc9ePCLo7lmkgGeRr9JJwSDPC+8P7184Zertx6+
m6ood+9LMR1jtzagYGAhFogcu5SNuaLtba+EVX0FyeIvQKsusNBOHGaAcmQzDRZjCG5wkOuFoaWk
YJODDg5G24iUzwXWXutYHNXYNb5isNM927JoSRHnvHWOO6LWQBAn+O0lSO7Wsw46BzcEd5apRvRT
O+JZn0Teh/N+vCxBieW0qFpjfCmSSqDd7rzRB2za/PnDNOLnVgW3LmjqybJ5OtLwwij3Qh3xGkSn
skDWXFSxFmbUowJXivd7MYisxJq8JLn5Je9WJUExMLYHdeOxJuTMkYsAAiBZx7r3BcYeJUmumx2V
mFfJ5iVQT7kcyqTOnCnWQwf73zOtKF8N+068/uFZSPQI0GuePEGKAFyM+CNSpF+IEoA/IvBPazwt
ACZbWDPr6m8F4I37Fco/Lar+4A879sHE1ha+fzLEIOzZYL72HDKHrBTVSRHHtyX9VD+FE9oCSNvJ
lqOI9uKstBNuheFi+9KPYHHjW8yJ2xT+LCWEbsMe7AGUPVL21+XYDKV8bCejE4PKtLJxazpIVYup
t2VwukFi9lFQS5anjUTMq/lkTnOuN9/9nqA4Hx/baynjotXfEwq5bEuGFqrRsc02+n9FlgGNdpXe
iwdXAXiKmaJMug0vLS7z4gXeHBrIFIXa22+lM1cUHdoyKmAvBl33wPZ7KsB8ZJ6G567JiZ38bC1y
FDSjJ38WzSP6AFNIsWAckJqaGkhoGUWXohx6MYpaMFwaCg2Yz77CwCUmiWUwBEZ5ZJ6tL0OLoy50
g2SxzLqN/Bzq3oS8i6kmLCL3Hg1gzj592iloxtK6QuRLKqh5S+oKxCr1Q3OtIgQivci+yN+Ygzwx
8vkd9Ho3JosjwaUp/lvM9oNuFQ1C4y27KxFHZckEU6nbyEjzNLW/Gto/AB5KgPleo5HiTl1vQ1iK
CDX4ttYLuux3KEYuQAJQGyjZIcEIZZTQolYZFr/MEkApxrYn24Xt6zNXVSdspkoOVHLyNwQNnhuK
MtuINNmeAh0gnBBTWQF88hVA8kIT+ppom2SpVPIYsy2Vr8Ae3+/USgoRTR5h4nEjPPHkAZIVo1Yk
SiCk8jlB4nCxoq9kQ2Z0jQfO37xt+/dSD4XMawJp9PJFYoYS09rUQtLsx73/qTc5Et8M3ctS/Uev
R3GsDXMXjY+cjTfzlW8QQMTxOUrCChRKHNUU88yWZBJefNd6YRiJTIG8EGTUwXoZ7+b7bcGkQ776
X6i6RWBSkXfKdQ3DWELBQUPC21IUTomj+mCKYFKDf+qfouV+HMzMDG1mVmLX5HZmKJcxUUdtOMLL
wodcH5Lw8d1DzPnYQ9IzqpnYmzCFJkP0G9e7xP3rKhObucuPzgYzlT2vQKpWwlJGrg4bxvfJzzda
2g/SWjaJLvgmz/OPud0Lyk7npAba7yU1osCr9R4P3qqfBECUZ4x2WDgLfR1zyTfJH7QSWVI9UWoE
yUNfak0AA90fV90wFlTC1YmjPtJ8sLDT0SROaBSdtPNeaQHEr6+PeqE+X0KYE2IVko5UCrSObdZB
2ZAM6MZi2uai6CBa9MzbuwxQEIht5uxskW2g5FxsxRnRPqGoX1X5nPKh86vlhFZ9jTCxrh3WYJ/e
YlBor6cmAGaeApOj10dE/NxP5Z/mMS3f2hw1r5D+EKp9nR+aP2u7QKNHq35Y8ye1ENf0KPT+DWTa
mFykqPiGIcvBWMhSKlqh6r8W1kwyz6b5jYXP65DlPcCGeACTZq3on3fLyvna02YN4THQCK/hET/y
uhGuVeAEXaaarDz0lL+JzLWQdrFSYpBS8/0nNNuiYdBXWpOgYHpjP3bqnz6rnend9zBu4TvDOsa6
al6wi10XXkXAPU0OIdR3XdlhhJOjRp7+dOfA9VHc8fwMZsHv6ulpE/ZnotMzp1kPcBu82eeCGaV7
nuQDVKtpLKvbm3CkJD6dvmhdUGqOj4dkneQslnK0c8JYyB2w1YbzlUDnFX9rgBojn3CpOPRja2n1
tdxj6BG+E+7jeAXwcnWbZG6zdK9zSDPuuF/w62jbmVrMBzOmznFLerjdi0DTWOYUEhTm5K8IQ1mg
XFxmwipSLBcuDWI+EnCXMZDq+6//BB45qMQaX6KuO8tGsABYeMa8sV4qBZ15NKoS69bAdY5zdRdJ
pb5PcXYQXMLRGc4U+uwtupiNi1bqTQKgFHfjbA8/Cm6GWBGTnOaV4E1JYPvmpfFtf/Db0d8ZEQjv
/UvOfu+7CUkWGX95INw63tFAf22u3D1hh4lF09Mg8w5n22iP2+pAUR4QvKe2YXBxdHbEW8eaj4N2
H208zTZp2D3c3QLWnUfT/SW+cJzkcnFtGIXBK4lqQEaouqMVqKFtVvuNd4NPxuQbYertJFR6Ri9W
McXxHanItg8rhjiWKZeYPzFuziiCbi4L5Yjb26iiylm3CJSiq5x9fRoeS9ouEPDF5sf9S8Gs9S/A
Ce9ESqy3C0Ov15nm9SvvYKB5WHRRgbrRJpv6CXVWlmDVVM5k81rygwyPLF8QFiyBUM0cZM4u0kca
rE6Hxtdu9KhLHTO+0S6Ob1iVarHcGVjHFIw2LGePbCOI2eM5Y+bYsFLTiE3wfuEaJaM6XgUfexoe
29cCl2kSyIbO26aa2Q7xjGAhh3hJJba5j3JgIp2aOIvilFT9hLBhfnOM5oOI+bVFsVqHQGTsL/JO
gCC5LjyEYp77ETv7kcIZG9C/FUdE6O21ayWGFTF/CKC7+5jlOR7hLx1BX7QryXClTcMWRj3lyahF
z/oeF4PLZUvS1DHGKX65Kap88wgXlHlpHj/34GmAJuWg4VY7y1IMx6A3ViknhlzuxNEki/CHwBNI
qfmQ1i5YyDvQUeeNmgByi9U5vDabU3AinXzsI9gwpoIRrex24yDP3wgGn7nK547C0F5CwyYWFcbL
Gt4g7Lby3d2NNC+rbA3DkY18ZNB3++NXe0Ytw9vuj0AT3BILcceKAR96M6kowj1wJWJBoehM5U0w
5zmQoXATbOgYkb9b08vd7KxAZiD1wqZuCfKWXN48XLC4Yfazyrf3BuXarL7GtgGp5C95vMOkReNN
4zI9bxcrM8D3f0iOoAqC7XOuO5bNws0MXpU09Cp1tA1ZrJT7GMpD0JpxFYDHFx1B0k37HrAipXan
EWHbaSHO1MtrCx/J63bxFbVe+71hks/WfjWSN2nNdVI5lfXNnjlxkkr1/2C9206ScpR7DNHrEPHy
fnCwO9nbgVRUYy2GUEtv8uKr6mGcJD3LnGMs1yUGYUet+CiR7NaBI9NeYwUdPBgCpVPVwuqftR93
5ihW/InMXoolsYBnAVNjLwseHJ2FiDW1qUjEsPdiz+wwevLosflx01rglw4iAZwL323/mjVHLHBR
/vLgeqQvXLrhkxTPXsERIlm6PoXTGC/u7MzOHZ3ciBT3Kb9FQlMnMi1Ld42N93cMJ/o+MK/ybPRt
KJEV+1aLwHOXJ9vCnoWAXQ2FYbeNeNacb6zbPkeoEMYhWN6CAGH2182OPkKtSA7IuD2pGG3ISXaB
HbpkqMDTltd6N2FxJJ/PHzKSk2ycq9IUecdwm2A8HRfqj51F77pzSaTMa1tksS7zIREnDBOqeu1I
ouWvfFENVe/Ad8svUZZye2bX6ehnOTbihqBpAx7FxOXyZDpzckN3v7KpR2w6YxM3tru7/lGJGt30
UHWmvx9I4b/IeMiVE22E1jYqhbxAVhXEPF8qE3MAxGJmQgM/2PmfId1R74J7ZSI1VPN5Gny6d8VR
Gf+c6mKVXbm2XTboe4YLIChvFH/2D1G4PdgkptNYUDsNZNn87ePl3rDoknrgDjjvNnRGoXADMRFZ
12zigVb2TlorhwCDZ5P6RiKxcxTRJM++ASIVrfQZsiuv+WKSAmJKUA/FCztkuWQL1zxup376x/r9
CYXHoWfYLVHHz71Pg7o3/gckvNAj0yxJrXLmZDTzDazVpEqpSDTG1MNSLHfMgRHWmo/JUHokdwl8
oktYkKgi8sf7vV9j++dqAPy4YytJVlYed7ZkKUW7iLL6qyhU75GOeo8654BdnMi77vzU1Rhfydms
5m4klvEpWBx2gy8eyoWRYhgrJjKQEw2c98B2QsGGH3YIzFbvrLOcwjJMuZ8wXK2MmyRZR334NSLm
QGIvokb7oDqpGZQ3bAEnl/NzM8v2K/uW2n9zF//ovYJePfUQyYwOEtePDBQqb1f1Jha/dtBvQf/s
VSS4Wsq2P6Cryz0882Hzd6K8UU8+6LfLEUE7GLrA6dxCRHiGV1jEE5dagv/mD0GNLQQTx8sF3B1B
31euTVa420HCySlcx/u+YSUiK3t0HLKx/riiDHpQHPC+hTb47V0wx3h/cElRmANLdtuo8NO2Mm5U
NmhfBHDQPeL/9z8AG33YF7VefZ3VVG1tU6QS45Y5s5eP1uUpZ91JqGIGyjbijdChJd6+rM0XxNA5
olA6KFVpNLu0F2HF4uWsnpjySMr8Ws2XqaUb/siBZkivzdRsIwxxXWnaqsUSvRnn+SH+uRn9wy12
AIkxstn0WMC7KJMuZcitWEuzLLlfvP/OyCZL3iVN+pOrASHCfYhWrGCobSh3zyz/ONHG4HuMphNL
nZswX7yGzrDuYIg/MxcXFu8V86hkpDQDcAU0lLV7S5i+/260IRlK8K2hq+hkAtaC0MvMrZkutqqe
+4+rNzMC3VCxRkfBteSkinKI9MZcePoMH5gJrXFQYBXKb44o6Is2GkuhrJlgtEFjq0wF1VgvyU0i
H2Mpd++hNhX+VJKATaWE0salJuzKTyWrYMQM3YzKpvuatcQoqBzoQv14Kc3xSh1CDkjep6sVjIbv
46mrPwWiKzXHEvSbdIt5W84lc9B7VS6NHkBx4fLkJjsB8tlPRTqYtwXC7Dt/ElQO0QmlWmBUQcVj
PNsmB3nJhLDXJQM/crcrujlo/3avaamY0f7z3NZnzuuZb0Fa0+XyIWYufojhQMw3vPLUrX4PB3RA
6xrE79k4kAycWcKk8gE2cpmFufzW9rRvgpE/BZgRnJtOKOV14nV2+8/9MuKIScYy+O6udnC3n60c
qClD3xr2bfKMS7jp7b63Ik3n8Kzjdh18a7qC+tyG/P+sgw9C/2d9n6la8mTTzQ9Jxz4MmxLKP/Xm
4znGRSFa0dGpIL+ZXJLZGZKrRngZAjIGaMDwWC0vGcIgZ/1HmKcHqDbcvWI2jDZQFjvx5No5tWzv
h14KJKdgwPOD+WZi67AnwYKdLjxd5DnKNYrr6nqarr2XutBQCjjc1oRrvLiVzKT9BEQ5BAivE8C/
b5G/AmI5Z7I8qN7iuJ+hPFxS0ez6bBXf5+CQQL7FHPsVivk2fWm3z4kDnkjEUekXgoopkQ6bLOwT
XsxWwU+YqW8mbyoW8pLllxNi0l/HemOX+6TM0Cc+2JnWuxeHXCMX7ywXaSDCsGLHzk2twT5mwx00
lur1kY926i7hM3p+fNvuHp9P35/y5ajdfy8UhbwqDmBO327/GRFy7UbPP7WCKx+7+rKoZoInhYK1
3/BVlbeGladMVF0v/mDl4REBcYi5qwvckNleR9uwnwdo0KHLcP2FVDfVGqFyapejCSuAbrszWaJs
WS2+YdAQxNCwV1b1tyNEpAl0oLfWW7QY5SQLURk6/AJ5OFqKdHqYFA/HHGK0JOqBoSOMZIMHthWv
xEmSSTAy5twQsL9i2brTiVVP7qYTvePXMKy/E5LzB5pqwVBau/jvsk/XL5KGWWQpun5o0Vg1Fsso
ao3DKfALnOJRsJXE1Zly+Ysd1QaBeJ83T5DejlK675eHIflIXTDyU7JrfBEpeUdWuYRhWq6HvlsK
Sge3tQzCK2gj7XWDsaVCQ3Nm56YDzKW5T3EFybn+7amjWhoedO0vpApHAw6jmnQEz2fdoFL3TSfm
Olxpkanc1s10IXzCZwWKPe5HRhwGVhMhROIjmJqT0ismZiY5PI05Ynn8LTZSyQk/gFn1pt7KUkCv
WYFZiSMlzjFt4V3FQzyBUZx0wdhFVBf0XwbNm2hJ5wjHIyiNXj7M6dDs4mkrIJoHP5HxUh1VLPr7
0LPrfPdLAGd9v/hVU5GClc7fHZZ3HwLEq+PNjlGRS0QxKdQ8qebF1ty+y7Uhm2SGvHAWrtFUcyNd
jdN92PbIqFcAQNw4xPl//ZZqkShZshndAFstxcHTO3XTF8TxGZUK3bAFsTftro6Nnmdu3X2+0GSM
dfCXl1uv2Aa6U2FTzWOhIcDMoU4PkZkkl2Ty27lu2EAnGRavR5DPihWc8n+La/mAZTgjb16XPOTu
clI1emPHsa/Nce3gkIxq49+xlmy3T4+sa5n/Mwuqdop4WxnNdn4Dfi+sXpTCYcCwJwy4A51ilDTB
pWvnAzFA/8X8zVRsX3VCozMFN5NgG/+AcwyO82WHYj972JjzevyW5/9gezwGxBcgyEenTgpRwjhT
d/6baUNk1kB4o1KE1B0tKv/tugZokL9AgZ+tfLjgFPAAI66nUi/dKxBKvinuxqLNZIQwyhkXsa9r
i+le7bFqZqXXcooLUitA/5CclNtKqOoDKg5nCpy8z5tntwn5PySzZQAqFW4F0F2C8Bn5cvoiNvuP
nsLRbhLOFlWQfipg8P0bfgY7Zew1rsGWn8KIR6ho7+fBjnp3hHdDlXZQreePjJwT2RH2Dxxd/o2q
b64AuPzX6fC/PR4nJSI5DsT2FR5bHNRERB9gg4WcOWuJPca737JYBxKgVEYt4tcZIGewkpa9LBQp
WkyUiGreycVaZMDqpRB0VrKIvVAQ/cVRT8KVH9rh9LBHGvrV6t3n4p0Mn5ZPwzAc0oJJ6K5vTXWt
XYi2MTf5c+lFenbu0AFjr+IYwHX9WUaw91WhPsnD3uOFWbpNqeTMArXKZtwvj7YJnd3+Efs0ekyS
WwFTZI8XaVM2M8/vDAKrjvrPx0vFdvrrL+3r2RWazt8We5XGIZB5o1qgvTxsAPrDUTuhTz3Pq78j
070vFSmcQDQn9LH342Vv0MJPATjgy71JpMjowMknc8SuTW6bxpTlmGCh+6Hz1Hj8o6+aOKxMRZwI
t2M48/OJd/5X+mzBIGpVl5Ey65wDT8mtEC5VM/cl7J7SB9UFi2PIMpgWki7X8qUxxb7VnYVoICZL
hpSy+pmbw9/scpxIZDVbnq70Zut3PanP5vt19DrjyCaPvAPDuYItEZgH+AdOZYkfmDsQHIbHvPKB
B6y5HVoPcEq4lVVV3Ucn8mWVFgltRiT9O9nYSMPtziJ3QnJFqajqAwAZigHhGqwxD6efClh0KCsR
gyaCN0aOW9fB8XafD7qIbUEM8ztGTgkHGMQl8oFuTE8SXnzDFlWxyMWabVZXA4GEfNzT9v6IPSXZ
EI125NQm8B3Be4P+IrIZ2DIont0ZCJJe6/0TPyiyo6pP9t1WBtWkN5avaVmsURnioTmaJMXQ4xT6
D4itJZRUrzdiY6XWafxevsiM7MU7xdwki/HdCHtZJLkjxyoDokFhQAAsoig+FUl5ZBv0V2uK9dbB
yPINqkqZLsNGxy3oSOAbfmZChMzh6rUCIqBE/vzIncFrI7EfvB6ktB8GEK6VeBnWIPfFw+T+Lwyo
Rs99tbzJo+q87G4ES9jzBlo6xe7IV7p+llAB4UwrIoyTX3yEf/opVn0ErkDGSiHwr4ZJakU+CeIf
+937nKSe06FW05OWg+yBugjwcCm2aBKX2woi+X67u2IOfIKw8rwyQycVFlOhYOOG6KQoMA+jcXuJ
UfGEM2WexX0mIttS+TC0obQp4oGiHj2tioJY9SKJNc5KYBTfdMQoCQoHljM+igVt3gKSf0afITAf
yEWaeCtsY5xDg9UCFyO7AFG1UNqSoWwLE46uW/pVjMvvuWZndbJwUijin+0i+RrOjK2Vcwm/g+Mm
RRt0U92BDhsoBTnUz6WMppiWjLI7bUuhiSgOHADjnpHt8x2r7CaDbOI9aEbjRdZATAjsXrkbz/0a
cVLkNQL7AbGrAb3bcinXQk6ccIbl4L/0GDj7EkOUr1bT/sDaeLlUrJgdNysW6H+GPGM437ve3DwR
PsaL0JiZ7AOGAbVw43NLHRSu3o7RSrN0JNqoDP4ibYsrByuFuiraIFt4uHO49dbAPgSzOUrBdx0Y
rG1Rj+Pu6xvsRE135wHNw86/BabFRGNec86/hYTdduYS9WlAK8SgjYZpY6MZ7k8Hq8hfbEwSRftl
f1ng6/VDa9BYGPCT2VPrWxa/5VKR18EISPRhF09n+e9PXotQQbEHgVBIfAZJg9K3G9fcfvU9T4JI
7EnxYnxJi/FM6bNHuniTykhDF6Tl1kqXX2m44mKk+Bl+6/YKs9S7OgJzag8eL6OtbXx2pZzdxfZD
PX3w7PnkCNvpS/TsfpdK6XRGIx4CpHQzUcqPXfQA/cSS2YDliMLEzRVesvneVXWWlGDSqfIrlOId
DLyX3gLLYijSk4VSXPW7SoUVAh7YV3qDzeaWt8GeykNQCi1Ung8cSkjEpsZkr5BHeivZQL1k8iHZ
MpeiJAWyhcuI2PH4+jL0QAPgjMSg6aAHEl5iF127+jk4DrIZ6iiUmFzXIoh4devFYlJRCKZ7LSRg
GE7NlucS7lxZT3C0dGIW/G1m450pyr0PcoA1MCFdTDG/T/f3RRsB5uWldQocLQfuEKlH17iO+nyO
CBSYNSLThoVV+vvo9DcevIjGiblEVmtx7wRtGZg2TfagRL1UiF1XsIuWesf+IN1O/3Nn+t3wYdKI
bSZdQy8BAaJiCKMwZDAjOXS3ako9HMfRdK4qraLW5ax6cc0cFfEZSGEMKui0+DqymmpPApa+1XfT
08mM9L07b3ECXHRXHso6NlDKfAHwd4h+LI4554GTCqoxuRs4oIE4Ve/56MRD4KT6X+9bX5l/UUGE
QUUGoR8CPA7z+S2A7rn/YeyhIhhMB2fAUJ63zsl/3xs88X3LOIK6r+PYlX6BCBSZy+4OniWPcHGX
5FDrDPpAX8eJS/8Kz5vsEB/+4ZlU4WQzw+b1E1D02IiGTSAYQvwTMOcpPWjtSAgXg+hO5aXbB8qe
HsQSO5PPO9aktkDBrzEiralDwTvPE9SSueToad+tdwdFfcdBDPP30D/Ql4Y30EVbabdn0URP8W1c
7KDFehMadZQyti+Hc8LCzVE3adDrd7BZ4y4C2cHychU4nBW4r+pU2r0NLH+AsPEtnClQ+VoI1VNy
cvcP305NvZ2Ti5QbsV8akCGQ4mpA6ydRVwgWleVHmmuvxuJI7wY0ZgYLZc5bYQXEAT7HzItwWel9
mOMBRrWpqBiz+459zFDu2BR2UYHjVAlzFHQDlqrDiX2Fk/R279pAHxtlbb9pgEGlAdAO731684aA
yGzawohZPj6fiCds3v76GJEkbvRjN7jVF5UkNirHzfzyFSUQyNlofeOBihjm4DaSlhChPgf+9C3T
cvSggj03co0rdWCEj+bTzhRCB6SK7KPNz+g5YkfFW8WBgceXc1NnbWQsVeqnZN+0DnVvGQbX3kgp
sI/gsMWMit+dL4ylGyLPOzEbrTwQR2uGO3sd8tcMwssW5CNTxk0Q3ApfMrAnpqY8441CTkVPaOML
N8gZ4p05PkwQ8v5TgY1uQ2siAXI0R9MyQOFatbcfQpho1HsLQsRbVQlWcCigrez5q02u9JcBmTBS
mx9MqS/MgYTcCXZ49vMMogY0wBRt1zxhToel1FQgtLGwes0q3H16CsmQRifOzvFWQZBaroq2jNPM
nE6IyPUfTTvUwjJbJz3pmX2n5ke3j3osvGoFn+l8lEcUW6cFGBRiMbcPTj6Vzm/ZjisB4xpLhWHj
TgYBFNSa6Jcq84uoTcbbqj5Ga5CeyxqvfrSR31kB9kXeagMQhd7nMcFg8Xbh1dqvB6BRc7Ou8grK
fQ+z28mS5vc+8ATd+jzQ40y/xCDARto+Wut0/LsczeFJuHFvBs57IqiGKbIN9GJd1J/3sf/eyXTH
O8D9WGS0fSscPbLHME7G5qybZYzhTh9W9S8twk4Yq3xGoRFOC6Nb8EdzJrUS9HwwD5kfxjRWirGh
Y3tYpd8tn1HSu8ATJFOW4Wrs39idS6rYfzTkaFrd0CJddBCSdw4WLDcK+SN2VsXpm3xQGA+EvvF4
oX1ArNCx+mjG10DenBPIdAs4nYBZiNqoKGm7PtOUtnkxV5pQ5tRHdGj8BWvSyC/BntP4MffQpxAa
N+00ClH5DZNbHwm7mlIoZQ245iomasVBTcZO9jwP1q8U4nnjNzIHhkS1WBWhTVUOb0TZvWiGy358
y7nPpE2/ZItN1L/8lWgRvveYj610E5/aR3fDJNtJIFyA0PIc7d9+GlK43OngiAcTJzR6zvff9lKI
EWMYcVUjpnXmbiB9JcZCCkUV2ZwjtMAgEkn1eA/a2VRcHnWvAZoBXHzxHKinye4woJsH0tzWYxCP
lNgNFJt+pMzIU1vQVKBWZvJCeIF9vYoArrzkxtgOBu+Mojhp2Jc7Bvm59ivuC7rDKImTNpbJswXp
eJJJ400t1ZH3F+VNWoddiutUZbU7LCwlSf+E8qsarepEICD8qHAkrnXn3CB3erF+TP/OCwG8uyh8
N57Mb4deLNXNDG0Xs7LCeQIgO2Oe+70N+9sh9r4UnwX9z8Wq66rZWqSqwDGoVibV7N/D4b9wgP79
5r6fzd/E1Bq2F4VyDISkFiLGWYqdFkEiCi55aMMWlDmxkDJruEkhSUFwaCvR3LtaA3Lc5q5sQDu+
S9X1dHM6ksl+yt/n9PVI+CM+gcPUmwyXrW8PNcPnOhy9pNC3TgOTUZOVS2N2osbtsdKymBna9PVV
pPgKfyjkXnAX4VrTqfJv/SLutlGFQ92O28Zx+ikjZHhLkTVxCOnlqghy3utoZY5VcISBBDo8/kih
6jCWH21gClrAFBGZBTyuVc4s0dVDD1Dq/D9j8EAfRiKCysGcEYub7/qohYpqvmQyZJ3XtnRrkOUZ
zG8WKNggncLjwoEpKhsKOqtCdEzAc8/PGs26Z66Ijf1Xk/n38NkxhOR92lz4HpptTb8e55oiyBG6
caGA6hIUXU/LzvZ8o1EYxRL9TCkoX4l2qbX23R6KncC1EDsZFFXdRBPjCYejZbrZ6K0jfdH2kZZZ
v+sPiYhmnZqjK9RWatr5Zv1lSeAJ93KiVeau99zV48Be/OWxiNX4cEHcMOJe5HWVSWjHQGlNAyQX
qWQ7qtDo9RUmGgNNoBKS/f2lOBvTqLWlMizdhN2xKQs1P4JxnzQ30V+VOPx8UiTN+3vAwqEhCOYS
aL2xIYlLdR6f61rVO3GYefOlSCwMxBoRjbWxXgD8L16rAAQmfqickO4fcj0J1vk0SH7QPSl+MFX2
UG4T/Sn6L3t6Hc4XWg8iJV4DYE4iNK7eGKpQwqZ9h1LVgqe+GJFvrwxlAEB9ef0CZao31YAu69+o
Hl8yDh3DzrOPM0ZXtShUKUOVsVpRPteZfCChtYQRzWaBhPywvJL6V3AbgPaeh7f66nQildAwW5v7
XbkEunqLCQRqF2UIsEux8wpqhPAUNNdChgiomIcZl7J+hqrCGcQDElKT79nPMEu9s9BcsdhyGf9K
MT/G6A4HJLb2EmEWCpusoQLR0uAX63FFBn/Mz4Ls+AjRVUuvXDpgSJL+YsQx92CHhbbolcSDZgIU
2HfVmUvoQVsxaNLyPd2xUEISCG5TjOSIFtoWl9yMTKLL95chPm6Wi/T3MeIVoxFvD2yPMt6el+Ab
cumzBqm1BkaoCOPWCOBB2lu7MUW9jZkVVr0cgphNP692zYf855bPiUErlcoxBP9HgSbzeUmx3Vp+
EM7xsb+p9CzcgCcGMOWTwC37wEUVYv8Zmzw782XRpqduptvpzIeo8iBWTScQ5RrorK2QpakxRFBT
qvT9XJ6zyAzLigmqEbuFU0VVwWFCo7mUCuKhft3ji9CRGVHpv5iXjDlt1Lf/b3+47uATHJUCxr4w
yK2TlbRhm06aTlalBQcsUF7M9BakSGvuwa6jFYdUVKxe3Sy5ZRmyFMAfIAnxwt5DfklL/37t9AuZ
4YCKGip5brus7A47XukYxZOndDfUDFtEUHPMxXSkv7c1beYY4JsKvD178ka8CvL2DsDnqVUvA2RX
D7TEfxRDeXjnbEbKhqoqrJiQqBqmRTOjomuB8I9f2JXpnt9psD3faQC+SvcqhgWZrowT1yrbeBl1
uY5btO2QK99Am8WauT9u+dv8uoHJNnBKOHCsdJxNndOYwjuaSLOjNn4ZxCU/KcNo+P8zMLG4iip/
x2JqeO4DP7opOrU7b3UTix0pwxaNwaTQy1zVO2KxgsQhPiygsJ7krdxR9klatWGfFjcB4BY20EE+
PoA5ydBONTO8Uq+EYRiXovaCxImMMCOGllJkcpRYyocg6cnV7i8azzuNk446MbJImcOnUHclsOHy
hDYOeC6tGXaMrOObwzFlhqel6BvCLsUJUlvrN8CUNXI9vvioO0LXPXNzl9E+wHuvZF1w8AcOZl1v
knZaefrXEDZzB113aKFAMMYiWG1bPK3wqyfcOPlzD/70ujxT1KE2+ELMnwDOZgzB7eQG0Maxz7J0
aD0MyYlwnYwHs0tS5o6Pkx0aG27qJoJy+HXQzF5Mkw1Lgn+9D+iiDft35s59cfoASH1yxRjj2hNI
pkkvfxtnRFfkYRzJ98oGckP+a7v2AZCO9baFN+wySQCIRYcasyt36hIZwWev04aUZGE6rzEzK9lD
ZdOgR8AJbY7mlStCIJOCyQdCPadxmI/oUOT51HBdw0hAf3yeRWhd4lhxxhTjqKdvnPi69l0nPN18
hPzAlP75KyGvNyRkw3XkH5dEDtFwTtFuS649P2m6DOD2sIsQv4EYGnDy+4pJbG5lFLN0IcFfOObK
Q4UQW5NdJqKmeZ3iGVYseK+TUyFhDnZyfQwS/OPYPtb2sUgx4xrWKroFli39Sy7R9yOwZ8JwqGYY
1o/E2FXvwoSjpaFz5rL6ESdXOJS2akNlOxT21IGMjYZgvYOYMcDu/zPMDiP0krGQnljHf99y2iWO
l0fYE9sXK15zPIVHWSR7GbjiEg6qnRgiBNp2P57R7nu9UtkKKfsUp1GSOCVxYcJLUUz0X/U36m9r
xr+Dl8fyOA9wOrT26vQmQhxKO/o4u5FAjJKjZxBMYOLAb+FVYk9sFC5/mlMM0bsr6WyW1XKxhqsc
UMjlrkI0lhWli+wV4pEcFqr7uj3HY5WJehU27EbnWtBVNpJfYxyDc36EwxMq5Sf8k/vfpJtT8YRC
ac+eCqswHHFsP9ODB9swa9JWzpEnCUHcxa/lLH+epEbFcCV+4qEKOqHTdTxT/5khv3y/duyuGCVY
cz9x7m/zkILfq02RgRs47ur+Qj8yyegXOcEa0oIH1HFQEe9lPFR0EBJlHGzX+LwsX6g7whbAJCWW
DJyRz1+bnq3SDF0WK0U4SJiUJ9oO5jVNWdJUw6ksRHv65XTU6av7GMCspbNCnQiSW9Z08tOe/Fzc
xIRsQqZ1jWvMr90YTWKuE8d7Ka42IpXsk9NhadYirlA+jmKiU6/0J/0ORtq5bSMrGAgbxl8yV7Tq
dKJ4M3UxCHEYTDoH0UZfbLQXMjfdYcB8oE4R+VF7ri5CItF6saWcbAQF60VKyn2PR8xbr70fvVta
MKQVpgEGmFUVAiFu0o4NlkVWfpUIcjm8PkkPuIYd84YwELgnZkx/yO6iKUWI7ey9biSxQsGFgKCV
SlXTAT7akZDBN1JFciN83Ok6R4RDHNW6xMkXYKzE0anEMD3kwgytdTdHibtjpdz2bCYaqAWL5CYQ
eGjcr9h2owjG5kO4AZTXuSrw/wMOLMWk3B7ORX0wZk39WXh/n2HbMMnvsl+J2qnuvDI0UKGkqCEh
hL9i9l870VZho0KSX6cN4X+VVdcN3kupBLbPvGWjxk8Hfh4XPbioI320xTy5CQDuUcZulDqCIdHj
oTNq96XBknM9KSLIYxam81/pdj/ySodXc6yojVhjPjNQWvNA7SIHy1iKD2WOXTCkV+slXEjDaf9D
xBrpDOQQKZBUXHEhzpeiKYW5Tdvmqg+l4qfb7nsubziRRjqyWVbkLfeScNH03fxY1fpXj/e2JPLJ
681I+ZfmuDDeTTJdv3TTYusJqAGKNuY1yeSLjnis8JXUQxC370F9VPt6ORxIm3/Sfuy1NmDld6Lo
56L9vU788x9KdkTQFWvIcK318dOrwDRnYXg9MLHkdxt36pWJ51A1Ho4iZT4aoHqOTcZHODn3Dpsz
OmXqz+DhstvFE4yfcuVL/NXCd9Jo4VzvzrLUbSLJtAsabZKX6mMG+jLIYgPPeGRmh+DyWvipDf+S
P3BQ+EyzEJYqhTQFIDzjR3Zd9Gl75fiaYdTJL08yk5fK3dSXEZtswFkfEu6AQHgXFsex3vZjhhZp
4j9Id3Rp3aG5epI54gRzyw1VNWVfAHPaNtip7DWLk2fOY+6peSQcUfYbqrN1yfm8LWTBFktzjDW1
LZpw+hwhXuRDiI25tYfWnCpgQ+HCiKFrWEQr16UxFjuun3WrcjRGJFFYD3LL9VUZCYX3iqqvSUGS
ALZ5VbabII6CEkWn3hK+6oIGWoYfvfhdwAsUE9Zoqen+TGP6GZVxaSCPLGEf5GZqQgsfYuFn7Wfj
FVtxlcfSvsN/578NplxJscxF0K4oHNL5PDha6WQwt+hoPtsb0eUrfFEr/+ObrMv0C2s8NJPEI4Ok
kVXCL2+T4iOh4bMswVDACIT9D8hRMzb37/uwNzaBhvjr+wOeagW3dNJgpdLq/aQuBc3kL5BzGL9m
08jH+sNyt7q405pVcCaAEp8EyTLpdUW6aBImDoCnyWIiTgmCOHf0QjvLj3zUVDBnhE0uAfZAkUGp
GuatqaIUe6fm3NgjZTbY83nRMGV+RoiIefV1zHrBOhl8pKUKAkf1OkUIcO8cyaX07cipv4q0t8e1
l6ZgbcOTAYeg/s7FXpvlIfS8JvggHBChZA5oqRrrb2iEK9Vv56qm+YLcHmbaP4TiI2taUKbbMsb+
9R25vmM87mFopnVjKhQqvP5AedWMZWtk+UlLZZtbpaapPwbfUeMmxJYMnMFzN3NApbJEfj56EThf
EUCAeYK57xmpZuUp4PXVPVLFMeGbulFp6By135j9CA43bg+YT1x+UEcAPq4YdbSul3RF/TgJ3Yvf
nXZPDrgeDo3VrBC2cdUCAuW/2Se6v8GILLmXi8gRH5HxvMODX9rP9XF7YZmlVHHEWStCs6raVrGO
58XY2op7UPHeH26qq0QS4zn8ni2PbDUbD8k6BjbkVL51ttSkWDMC8Y2QaxNuNZpNp6Mv2A96ekdm
J39u8FtCh2DgljJe5KykMzb6xTYNzBjtKwLO42QwYRcU1g3zo2AiEw+LBRSUu30s5KTtHf8jpTPS
Ybmj+0hzYFLVyqefUq+6Yxs7OyUyn41up/iciL2LIaA4/iMhfQ4lFyQQeQM7IY5D2aBZ0UUGbJVj
xdrHBMynotNPgLVGaivBLcWhiDc0HNcBkhpLsA2dBhN8plnNg86HltGx+KZ2Zqa6nKrEKYQc9Vhu
VSzapNbkin+rZum94Q5o91n/2B0pnccrPQ1AyQ74BihZMA+eKJGT7aTYDWYsDznp19BPyYdETe75
qEDGeeG5rpWdGWm2mKkUeqLtMZzIiWesW5W6njXJhA/l/r8SFXYRqHsU65WmYPHcJd+19Bo3khpB
jicL50nhzRB9kh0VSr3MNebM23bvRXr9vj+8nO0DS22/+3KtxyhXBA0lvm6pr6xtrOtztLYQdV+i
SHj5LQuJFtKYb3gCZDn1fhq/xNBgdAJPiP5v8tlVaBNC3yX002drOqW3OFwpnZb+HMDqIuHyOqqU
Yzdg8zaRR+Vqt6hj+q759aW/cXDVuRFsZjs4EiAQY5W/lTEU0Sm/ISxM1BKvvueQyTBCLl0ULu/Z
eOmviVB5L6Tv3R9GFF2XvhCEUNXCmTNjid+lsTHtth5nGnuc0Hov4QTEkCHEWzPZbiIa3KHOgyDv
GYAMg1YwKKMrbad6rZcf+I0AftDt6DkoLn868hzP4rw6Fy8dwRZeOniKHwu8LPkXgleWbF9WMaBi
Gm7LMcltursGAsIImPFFiWkRCl5IuvISKZbJq6F62K9Xbnnt9uIOCY/rk90XGF/JSFG8Do+Iobdx
VnK641ga7W4y+KY3CMDINt8iPq2LoeNsmQPBoIlPsEiu5fBwqisRHgdFGY0/3k50AfqkQ2KCKtLb
j+krs3AeRLkCclbGmxICYzoEzAOdfIg142BrYuC1p68Co8bnqK8ooOnsY2i3T0M2ZrMcny2lHLfy
8tR/oEw7I2Z2Y23un4jtFfeLFeIv+mzwa3WiyOILVMKpSfsPnlezZtVB0C1Y32JTAwLBzVOZxwWO
8tmFgMhupiJzet5+rHX6menslPDUs9KCk5ApLQaI/atbk390o0Q5Dpacu25tTYz3Z9CpN7PsNaU4
mKfybMLJSdK/q8lBE6o+GzNzpqXpi/x6qMUDOe5KD0kqDIF+OJ4oiY3DzSdzDbHd7p+Sn/AxKQrp
rutBoxE5jm37uE6o12An7QV+2GJ61cVu/G9x+w30/00X1VEAZLFSy3I3eAy3LaZcvWdxsgtZcKCr
sk4vBGeVYVe2spRtq108LiEObB+OodncC0somxgKBm+4YNlVOR3sZBDycI0L6IaY/dr2mhpZDV9s
PSi2AgEr6ObKiV7zFFIG/ZnJRWaTjLr0c6BSpa0N2vyGI6ngyplX/uxMSE30S3bxC4yXOy8w7RCN
hUGpEPQudfCbO9EolRUmBf2O7LP3GBo9X5CPnil0X8BwRf1i/RZYR0dnhbpqof/X4JhEMSfL5Loi
citN6OUs1STtvT4Nb5iU1LPYmrXZdf7nTwLnrr42WQ6Ck/BokATMfpT/A6CvDaoFGCrImVY5rB+U
+iBaoDIH66sm6XkbNRv7wS6RBeh7BSjyd1UF7bZQokCmuWLm1BOqMC/NV1JdKfh0jfeLVdH6CM37
nYYWyISZ0vcde8bJEJjXolwGt5fkOpyzZMcN+AQi0spo/QSJtPgzpAkejyZKQiCtPW3JYx6elSuC
S7xBFvE3y1NSLDZe6PUbiTtMpRIoq5xJQXiWMb4vknWec/ZC8fpaq8kayxXNN4bXnkEgMGBrVXE9
vBOkYoATpst2o8Z3fiphrqTpBx89iIPlDLVJhnYG+h5xTbZSnwMfcWda3uoP/1pQS979nmVneEMr
Ao088shjjzTPvdiZ9BYGOwXM5QDCsBaOxUeDLtjP5kvY0aqDbx0ziL31LIvz/JyYZ1D6HV+FvTtP
qTgIwTDgWRnyItY5S7oZndbwab8CiTR3xC8OoSX1EBUOqN/4pYEuMxDomhqvcb5dfdZ+4jlTMLHc
cnZ+z9qWWivqfns+DGo78qGgCLqMoznSSSf8sCttKJSar1r9jteaw64nll6jiFa3VAEKwcLKQE+z
USt29qJ/7CpEWbaBwSGT/Lu/lRsf1DpX5zpZRg5xAPAeZiH1bi+mrS25fFtVswOhllkFiB+yjIam
w3nd2P2dUJ+PzDcZDzkM4EBCqgQ8hT8uoprhyMkqciWEVyzwMKOglbnrbqoNqL31sHNdFVovSFm3
epp3z7JVBdiIEFnfW1xiCjZwzkJR9QSS6iUZvz8p+5jnkyxpMt4x/xagsuJXeUY5OyGprVC0buot
Zsm+SJRoRWVdrKc6K7eqmbvr58XmzOd7sJourzvERIjN+7ZFXWrfHigsCtTQTMJ7Yhz83DABGuJr
wu+/oet3E2QsgnI31RJc0ctdcp7dK57XMHyA/Ho2UWfedWHaD2yL1Dw7dORXeIy7CJdYhrVSTd8F
Mh7OFBP42Q5bWUR3KjAXMsJ1xkD65mxcFcKgzRCc634Uffw6N+1fMNi8t7ei1oGAwsMf6A2n70lL
2NtbxSYL1+Lo/p3YH/5mG/N9zrT491FAMdJV4IfKZsogkXUkYdBNZ27pTjJYrchvSbxoIfyyROSW
FEVXU59egkt1Ieqb16TiMjWdw/06lbPdMFvp6/OK/q3yvec0fAsz4uoVwN/QUwdXIgX+F+Eda9xB
nSVWIpuvdCcQQ2PcYKSSq7SQRwf5Yhxy6NKstDIlH4s+1PvIFDDdaoiFv3tBxHA/oActkZ4XPoO8
wU5FvUcSnPwPJIyuMYjXBQecAi33MAzS7MJdh38ekkABDTAYwXRrjZaETRVNnib1FYKp+JWV/jJO
QLEjfIgqi4HBVqQeDzV+T4XzIc5w8jxH7gmiZDMzT392kjS3ut3J0ah5PSHMHgp/+QUunNUkX27f
XAmtDlazcTmMLt6CAxhMPQf8kROS+MnrqQSkfTHcNWaoHEmfSxCvtpDIpe14D/Q3jMnyghV4dpXH
wWJ8Mn5tU6S25psSaCdtc/V/HAqAql5LiNbDcRWGWtWxqtfhiV+OBiQGAxIwVUIT/j+Bu90/CMSf
XFAhazbQ8HCPv1MwjObxz4J3nIJfd+Rq0THeROvN1XkPA1gI2NpHLnXOVnlm+c5p7R29igLTDaC4
RtT2Vqd55E0GNVDSuCld9rzvi+J+i1ABh7gP2SVWOGddRmLx1GP3GFdKlIVSSXdWn4iYfj+pT2uF
D0m3Fa/HZXMOQUXI+dfm23rTwPJAcOTe+ckda1uWAHMdjpQ5M1Erz6ZtadySeG8he3IxjAgLKLBd
6iicZWeIY63JHCgNqfC7AMW030F4HnIfIS20UTf3fH7PW0bdaSFsPHVHX4OjSNbbORR80vYEVNxg
lfRus+A561+1UTIGqjiBNCSVhREChV3EYGr6fMHUrrBcXx+emoutOOpyaqKHSaSyoTNJZy7SBDsI
iG+m7ZqkBs9OPqzHDfLaKCt7GiYVmyf9p4ufq6OBrDrzjg/Jwz+9f+YXpLUokS8iVCGLibSL+fCm
Iqsdjf868PUI4p1Vaz2FXpvIw7qKXMQ9K3TB5oUwGWetQ6ANzCWvmXFrapjVAk0hFdrGXGfdYJ2G
EEAVxDCVz6CTFLFgtNJ+0hcNcW5ufYfgArqFl8noS3jy1UI3nXG9UKOkZSQ/pt9UV7GEGFFd46Wq
c9j85OpRqG7D2bH4ViaydtohyLw7Z3JOkIDjp9qp5PxZYN1jrKud9QM5CAnr0bRpMc8nDXeaWw7N
0CEk17rUnhMlnMfttL9K4+82JtL4OxhyeO+jRXctlHfwXaKBIXZPd2hGIW7JzA85n+oaZBs0eZ5A
4G56XyAJ0fHMOOynlITKoOLC/vtbvGHS4qIqHHMdcJfQ55AgDzGJQEvfCRw1WtReKSjAJrpkNi8I
YLpvSfeYHREziO8NtkRjUFLvtQfmEoqZHzSe9FC3D4SopwAhsVSwuIu2puBmtyf5ZVvZvnvsmzlY
4FtmQSq9GWlE/wJ0yp5ilKS2ctstGUQPjuvpaTq5trb973kbEebhD9PNA2/g4VR8pZreTc36msKt
SrFdaPJ3CEl24cloh0+iEr8PmVqFyOmb69wcFD6aK/FR3FFhTVfOIbOeZv+qdOukdAeELyWM72YO
RSPUpSmpbfhS7IVE1raYNdNxe0MxxO8m35b3I2JSc2zhVWBU+7VHWU2RUaD2Duh2iwSSSHKJ17t4
RGPwGNNrPGmJA4S1Csf6QNQPnWRFsSt6sAPBIYALpsZyTfl8kAo4wY/Fv8ju+wkouRmnq4k2Sip2
MU/Oc5llnTEZWhtExdTHiPOdIOXfo7iYPaD1bF+qR4qOgpU/Uzl9FZeXhDQVCIfqS4wR014RPO70
9foIKCiLz3rzML0AIgGdDCDBSPXjBektsHdF4WpRmLGgbjU9MdHtD9mBHU0q6g8vHE5yyTBsdaXj
iNIW4ScI1nM6F5R711m/LpxvCwISKg374MwcUgY3iavavwBNzDL4YYEdm5tRTcBH+dJkbP7kZZNg
yGGG8ePb+y+L3V9m5gmrf6i4TflnaLh05NVYrjmov0/gUSQ/isyMSgwK6M5u6OAopFqpnO2yd4jP
H0b4gNHVTV6zGK/lKk0igEv20e5PzkyaqcQ2/O/CpgXj9UzSh0+w6zTCyBxmAIY/aW2p9ezIwStD
gQSJEMBNk7t9LKk0EH/Slqt8M2FAszqUWXS2bDuR/J3qnM/lmEWZ/jsxnk4jdvW3KXv0iJMIZolo
eHg4XHtYRybkfKNx98N8JpZ/buWK51kRiTNqn53N/IsVMzDxWcwX75II6UdZMlOaxsfW4eqVXYQi
McU7gn00EWapr0kkVv+Gx8XXCrlRu9Vzb6Ci86WQ906ccAeaiuOtRtMS9C3I3Yr4OgC7T2343uuv
FPgyNzqGnz6aqM9TB7V/2IQRjxiv3B9QuWWXMwLTcL3I/Od474hSo+AVg86n8sJDXJaqaXzzGQWw
LvS4MT9TT/7WmZUvwF6XhZ2O3fZg84haL4vBtEjpslG8gD/VYw+iySOk5vycjpZlHHl81EO2gxR7
MRffxHTO5pKcHSa5tRUBy+wS8xPls6Q1xSWedkq9HIgslJRN3+nDMzBsVxctKNItY+rIiVitYW1t
JQpjrXGf07qjI0wltt/M4+UBi8TAiv5U9Vdw/3ETVrU8tn8DibHifl+NLeOFhRh3FaOTbE+ynmdz
4CIwaRvJiuH3RbQQXa51ax1jT4f+n9c/3uTPW1luPha6Jw3S3AWpZ/QljqKUz+44f+jRwRqxzDca
EVHGmIGTeudRV3TZ7Icm2l7ugAbLDQVqn22cU+P+k2CzqT6n2twVIPC0IT3jxau+rSOR3lCwdtNc
fuIrkfoVUolvBUOFVn2XgjYZfFphw5yWGO4LqFUTDnIOsfRn0kDDTSqP7la7bTd5Ktj4/bDNsnww
R97d6QdhILXk2GMFL5csGM7MrUuuyFOLkR5IU0ym9CEbVCOfODLDP5SjJxipYLWYx7feEsD2kW84
wvhENV1KedVOUeQ/zJ80pyx0xZJomAccrpuA3L/A9RDKXCQW/oPVsHPg+xwb2v0rRx6oNcSc3J5F
XwICtKzjhpwm9bvRQqsOWZt8Iv+K/JVKqD40MXZtq2lCOLWoVwYBJvOrCQonjYEwsFX40AoyjdVX
+AvdxfN5d2/ddnbyjlnyZPB/nbkARBufoSq8k6/ae3/U6JMkq7peCXv2U1/EvcgX870ANsnit4kq
tHb5vFRe16cHOIZlPRGRiXC1EAhPg8ogKmCKby5PRBqg594//rZHZmW4ZZJXfgjaaPkck1AY9ofd
tyBxHgpoBV+yngaqIsudgW9DQdgOBlXPN+eOgwZf+nv+jUGwHkvoeTRKMGiTC8Nmt2eOelJ6J/9O
yxGgBQstNCOeAaxF5nzxbHTwtN89XGoao1BxzMlAae32V6lG5hT5NdoFxiCgPwG4SPO0xP2M7TFJ
2yPa2UJPPhJjQEnIobkdTXT7gzSeLI7dneBaJLTZ2PXT3bucjynkxtpLi/h3l4o/ytJpVaHycp5h
mP54FJadf1ofSanzueQ1vXBsLc4jWInM4VKjlkzyczRGmOvXJZcLtS/Ru+JM+1X6fK1YRQS6wKU3
FFhJRkLK60Jd9fvgtM65KoITr+rKgNv81LkCOow8QaohvsdwntTuG9xyxdfTHSINPHqLrStweKrY
yty5lIClX4Nms3v5MZPrtXdBcUeevtMbkHWqVEko7y5bt0opZwgvbBoTH2x9VLRLMPZW/JcMTw9l
ydjIsZk7vBFth7IO21T81MqhUWv9EYE6UPDVTgY8sIgsHwOxkwrpMZiCrwFpDoJYfzH+bHrP4UY7
5CjgEsGBTmyjq4NWs8QdvZHb6/aKw4TommBwbVsvatUt2iVu21JnwQ2XFSbkclz24WYuq47Z4kjG
aSVAz35ZPresE7ugpdKo7ZjLrD4WCdKQCythas19U9c0UOZAuW2F7JPXE/ljEWTbNyuJKk5vXsLH
G2JqwnNLIP+b6frkS/4FjpwSfBRvob20NRM+Tm3MqdCzaYFMsxzcN7AOrYbcTJv5+2vl+8jdpgtt
SHnGg2m5QVAWSux71xF9GzZbgsNDAWx3L5g5l31mcDWT4e6+u0HuBJhT1OzB0BadJNNM7EOnPj4B
9NgzeI5sKXtuUuNGvJ1nzOVf2d0mpYS+B+9+MtAV8lvf0IQa3D2idJncwRFofyuUl4NQMT05h9fF
Vaj0qR4RCQSzDkzYzYxvQNYbfglknqwwLZZBZ5YMZDUWyOZoBwF0py4gPBSc6UPNDw0fS+8LrMP+
HZeK6UQ1lZF4jOYDa9EsXzwhoGz/rRlKyXV0kSpzTJOg1BVtAq2XvJew3iLAzZtvq48f3zqgQHx3
WC7c0PtN4Yt38D76la+CFgjwbMHxcadbfPySbKVNEsEmaxwiWxZnpFAX3YFD0IGluvzL7qgwRnrI
rG4dkE8KuvBTu/YwG7lUOGQuRJblROCLwB+fXKG2wzRY+8vYA/ZTp5ebMDhkMS/ewJLxBBrnhu3P
iJYWJ4SueREh0Lbdiqi4HtRjyInpxapu1TA55uqfTkfeK4fiT0yqWE+yb73ZwYh1AixjZnun5PNK
dtQJx9bMFW3uKjpaPNAMcGV40QDa7LChdvr1P8jFeyMU17+PU/hYq00LT4IiaQAAVcBN+/Z+jj9q
tuQFhEUZYXl37uRgV0mw7HcFsKR4joXNnQCeBgP+2NpVH+NmpspQtZZNtBDRfAw8Sqma64utmp1A
pPy3RYhvaVUIw3Q5k5uAtJKjZ/Cv48zPX4oDCY8R0f3a8FyIz84s9wLzoquqD/QfJFjev9DmAZAe
HqM4G2JMmsze7cOtCgPuJqJrfxE0DnKj4OfKGMMBffmcwm2EfjpVO7yokVrERS+08qr9zxF0zWYT
P2V7wVqp1yDB+Re137oKGWHucphYPm1VEJybHLwVwlzzO0V51sHYwXpmyB4JkKMSoWf27OldylQV
+wWbfyvfcs9OA07r1ihB+H3MXJBjY87tIk3BPgu0VQ84r7SCHChqTdmV3y5xktC4cfopLPWWc2X4
WuqgUKqZHZSI5+iaum9+vwUaQCmeJIcv03e28DYLdJ3K/gd1Ff4d7PbWLbCAG6OpvR7s2jdwCaaW
o+KGdlb+rKzwyjEWGQ+hOgM8LGo+6JddTKSAsVUHOGLxrWq6HHsFcHZjk2kTSakBahLMvCMRCOUM
N/JJ2Z1IDQosErrKNZoRUlpYl8QWwGveQkTKWoHXtBIVvInnXoEE6KMDGf+urn2yOVwBjUrnR5Dy
pX7V0yab+B2ors8bpqpPZ/gSkrKNwUQ2JDx6M2w7MDOzQI7VUZ4JYsrIjzmauS0bUg/SnxcWI1ZP
B0/5QO2DnD+31TBXLTOTvM1Ay7HhoV13MZ5TlfLkWXT2SPuhF0O69cRtxwEZcgu41wLZeV91B7d+
mtcIFVtAqLMdSAVQxS5arh6u6r3IvD53yrwpTu48WDlvUdkp5jtDsOOPEy/CHGQGuV/IzSEF5hm7
WXOz61dKkb5YanPgiysqGeJGN3fq0Jk0TV5cG0+A0PUnBtsZ2TzUmWZdu205f4UsOP7cTU/xgqDS
fvfRwNcqMBfI9XnBjtKoVdQcxDt3j/dnEPz2Xs9hJXi1BipVOMnKny/r4QJPmIFFL/o9QqJNCugf
9nldQwcPbSFZhmqAnY5UfQlRuJsGptHl2TWILR5eGou1dztPMkdh+k1pemMIPEK1m9ItFU737CJe
TMCxl74TqoV7xqJtCeE/353l+qah0KauC6hEGaCSeltdD3Sl36FafU0Z3nBJ8/zzi8H3PcoafL8q
hvig5BPLKpIaoX1TzltiNE9cIaAET05XLuPgGLptgEIAjjcBSq8abEh0KIijh3Ih3Z1dAItIovMw
HoZq5DTpmT+WYp+xJlLn7I5XPYQVD50DW79S3cFbZsebbZ8OBHOnJziLAADnLd4prEQlnLkz6kN7
DoJnWP+PWuabve7N12Nt3wBd8XLvVsmMtmy/LZTAbYQMhQxD+W8x5QbHTkOLkKKH27cD2iAfPe3H
VfowZl8mpho2APhlrOT97KGe2mGtFlYB25e8YY77Yneidp0jYg951jrlIV8jureKeuNmlu3HhFqS
UgeC/kjNNjPCfPYL+EkR4n0L3v8+LnLqYUEFfNdxN0GIHAnvi1BcB3tY1szAwrU89EjnOwdYT3WF
W8zG0Vk2L/a6wSM7ojBzR+jHDb2xsuFKclBeojBWo7nIfMyaHPdRR7Mpbx9iO3wY8MvSsnxVSFfC
QgFWDWcGXXf6i6H2JjTCmUs0iNxH+iNo1kHBFJif82prl963t94QBgT+V94Rkw1wUW0nnPFhredt
8Q0WEdAVo+3Njvt31zRjlirlQfY1xIE9+3r2JXhHc9N1S+ykwy6A8ShGdWmWcRwcTRHREYrkH+1K
3kALqFuN/ZaQ79R5a6llilVReqpu+0cyADfOId8q4+0Rw/iAhDpbwGa00gt+FINSCKA+yqD3SR4u
m1p5kvzA7bg6NvLNfZbqnAZh0MDYHycGDiXFVdxRw628GIgmqaXq9Z9dCujKEJjsQ31rP9K7OJYr
TOwJxuym5tPZ4DaB6xOcOBorn/BXgFR4g+ii5IKrbVugAfFig92E12JeKM8Ba/aHTsg4YyXH68if
QgSGCDe/qkjmYscYmPSZze3jHE/Gpg1cTDmZybXXi3ECsFTxIGgoTEmDxyZADXyxevz6GsxfA3VK
VYtmyi5yLoGK5ZK6clsxP8mCx8x9OnUf5DnVBb1wws+jpznvY20lYPOd8jp2ob+SkcrkLo7XKfYp
64A0kfAYCWdhc4deW1wwH1GCHOAnTvCubDtsuNOEormrvT1qUx6kMDOZxhKY8mrqzBR9BM4eXUdz
hkYDeMDmxALeXbAosA7w0Yz0MiYAbseJplLVG6OKXOmi90CcUtrtsMOQg4NiWvtjGP0Dzy/ZeXfR
Ql2/Tw1GZmaxBW0GfPcxf5inlPnKUk8OZlMAqf9q0wKLNoFHU3vpT7nZ3fFnennzYhg10lh7RS5M
xdBwqC5AwAIn2tZ26kxV1TeSHyFH5HIayMur9cGI3MIUS39M/1pQoFQsmImeosnfX31Nwq8+gEmo
to/74pRdPZ55yXFzLzUqcGtON9RfajyoiME42CGdU1lZmmCWRzRoFMjVuDLGR5Mbx+ABGBA/LGPw
cnUrYmUWCI//YH/Qbyavf+C4t96sZMf32ZlmxVZnz0nuaHxdYGiJUT5ojfbUvatCj+6fx4IQsSPY
s0TWAmngSo92bkYhLD/YfZHj6pIFKdRgDKOQdoN21T4POyiopPyaHfq/ezm17Ta3zaTUdVJKYHtP
JaAR38P1d7pfACG+ooIftoYjcDOsTLF7rqLntRfUBuvZnJON1CDNPAkRFJdysFPElXkoosKuVEZX
fTtLJSvA+qSPTD2BtxvyLFRiPZbc9KKHErGTcCG9d6j3OumCq6HIDhue59C8Vgmz8X1ErKtTwsPG
cR0VTyC/vpO8al+PdGsLp99porBR6AANsk0Ktqb/ShURtLRf3Jnvi+jDED0y0Je2QkWbKcMSh74d
Z7gUBfoTm6laK7ap2bUf6LPy7GMxguahdloYWtWlmaVfXvQ/iFsMePa6is79j2U7Wojzb8fkIoNm
oS7NZHFbKVwDhQ4J+63pB2tkEdWsI5m1BbTjJGqVA70Ypm6gpUBTCURo9DpHBt+hMqYjxHU/VvwW
c85MyHDiT7WVcXlqASpUtV06riF1hGxldoNo4Zx3HRnAvxC1pZyN3RcFJ3Yyf+5Gv886pVAzW9wk
neX1BxtzKj8iKkVxcuyj4Oy+fq6vcU396FQ4GmsVGd7VWxsom350AHCzgljp3p8H5WHNPRESJbVM
WcmmLVRmpN1LZ02oDo0x98y+6d2kcrvTXHiA03ggnpA9ObAaKHOPigQcC8QOjd/0Kd6akyCcY2GD
AHcv6jeBsunHxQN3zjDxqZ9jgRdudNNMBHSs88zMPYvRZfp6hTAPuFsj/v9jvayalU1Inyc+c4nW
ug7UII04rqNN3qangnE48iRqTEqeeLfFKA/BkdPLeuDPQpj4XuKymhEMLIkdNEfjVdD79mdRdrgQ
q/o7eYGOQ0qHKSCLI6YHr8NaJslVITlDH/LjWeSvB0rF0C4pCOhlfRWNIyGC+flBEOmgSkO2Mzo0
j8KZ1E7CTaLiRQfBCJsZKZdiYsp8yTOUu+cvLgOArzbVQfV1WTgOMuvNSHS7kiMqTYrHU8W/v1Bw
Rg9tisMdG7L+KAPKrGg3UFYjQBZg3gyVtrnnkcYNrbWlindCl58I1aHbzefjwppe1ga2DuQTsnPI
nAeLUzD1NqjZ/Y7FAMQJu5DOzFpAjA9NGgHOYp1kNsBjn/m28UWOOtMv68M+JAPSA7raymxdP2+0
6lvuB8SUAKaVjb8U7Osd43OJB6gzhrJVLkVLezsXKNPG26GcqMOYiuTiC46XvswSJ/Cf8EJvxT9O
qd4R9YPw0neuienTAQ/553AxTl6Loby/E/g4WE6hufj3qogkZjtHQgZ6QG+4oTJDfaauq4PQ/aae
LK14iwc6MWjMl4QHTHGYTaYS+lMObGKj66cKqJemo0Jhq5Xn26v8hx6WBKibPeN9C2vsHWsHCatj
l920Y07RK4UFrsVaplgW10JcqOBnFqmVrUJrHJFozWMZ+0CVsHTuh/aM6Twv6Pr/k9F/iNor2XGv
zC2A0bJFzZP1DyVJiCnZ3yDfZu3vFyVpKoVMAnKWO1VJljVRo6pH3DUKgfBbvAkAXgVpL76PmpJl
db+e4ljJBRQO7+AMF4R74OOiaQc36L5AjERPe1/+bU27Yd96/tblN46UJfLm8rPRmuxA1oG9ZYbx
9R+HBThP+io6joGwPFu3sRN0aYDCAif4v6dIB98XGUiZtHP+dYE9jWg1+JBopamNam1BSCYi0N4v
omTy5YPhn1fVr1Yc1Ic+uKBxSUy1Ii+Mo/cKBflDsPzZrAJ+5rhNpXyJ6jDa3URTtYoKx30bFdn6
Z9Tj4TFM9R2YK9PhxV9S938BHmRjBlYwmY7BQ+1VTZ5CMyimEW421SkCoPENOoyVDcR1/oQPxjBT
GliPwbjHD/3ehUI7KfFqbOqOHzirMsN03B3sJ/V5YqzdnqtPW+ZTqHicdBLxsIZpa5d4U86YFiZa
ba3yuRAVfSkkglpxjplYgj8wzAAJsKnAguWd7t2MTqMsQ25OmHLKhoZn+u4212tXtirf2SgsHZ30
bLbaU+8UxrZIjuXH2iLZCdSSdHz0SdmGGv9zfx0qht3ufhG5EPkAkoydyxDtvrF1c+pT/Nc6Lfzn
BmNcmzTjwFvBzk5GdtUB6tKrkonTgnpFM9UnD9ybg4c7D/erBqFEGQr7aNMDdC9dp4qphCRiw7VQ
krPDTafm45MYgdz92jMfHV7MSpJiwDr9V9Blen0CMRD5TVW/+Cveff4rdG6fr+dNX2QEjd9qaiV6
J+lwvyE9HhYmLvPZIsZBh1tgL8Evjj2mNnT7bKpicVMTxPiXXuiK4dgNpeLWh06BTgsMsuL7OpWt
IF9L1mFX6mJr/mSX2+RP7AUNGB8KmwGDvgYWbCfn0AlW/W7gWkph8mjKw1/D2O+tGasmY9nN1Ww=
`pragma protect end_protected

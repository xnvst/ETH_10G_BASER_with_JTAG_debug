// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
omV48M7SOepLCg5Ynd2tjglFZTWRsllETjQg024W+AZyzEKL3EzSGeiUMERbWfO/rxHPqOpOhFQa
KVRmsROoWrAb0N+yyTL3Gk/pKAmeIsvAZ0MEnPYWg/f8l4h9gjuSCtMxbxJsdRLPOtdX3QILyVd8
ezSxnUi9t/lNr9gm7FNwoWAJUkDG0tYeRQ9wf7rtLkVJeuOdBbCpqG4eRN4IxGxnjb0TeZl0rbMS
jzufPogqFs7mCvtUa5jTD1O1/4ekfYj+htZjUZ0AHvABB7Jfky++pbysbe04ruA22eOo/DR/rs49
R2wKni2VzQDUlamT0tV6/zPoWKuapngjWpXT0Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
irb0x4r+4qK+CMyL5LfarXCpOF8pd8Wgjq72JUXaN7v0CEgjRh0W9oEVkV83LkHahxINNQ9L/bDx
4y2ROtjp2hr4OoJqUzkSm2pW3KEEDz/AMUwBrRTHDvGuTCBloxT1kevwV3191TMbYAqCUKCLiRL5
UrDtlSwDCfXoKcddJ4pg5Xdv2wFFz9UwcVEMbNq81r7gnygP11nqRDB8CsQVF1xDq7/++wqk4RnQ
f316F+TgeAUIN36SOC1LpWhEoaqwd/tD+Ad8gBsl+PjK0w2AQ+U6CuQKSnl35bWN3HwFJQWPzQCg
hl2lY1DgynI8yWW8fHJqvQNZYNeB+ytm0mv3ja60QIClvgxMUy6GeI8+3cd2/ofTY7zP/GqoIi6P
bMUJZLPLQOWQSBY+UDr4EWmDfX1Q/EKJX7SAAuwb0DDK8a7n8+s5nBFxNixFdkbUyiK2P/Xv41T6
RnAVcf9kXA3niuJgB4yZAPiz7qf+F0P7DIZXTR+UCVDLTUj1CIuH0fDO4CruoQDoBy8MBXdzvjiz
jgBZVk60bnCgw7OkXg+/sTjh4NVC1kI4RauktIgTEEM8WTJw//kI9AYqZNy0qJC8NAN7caBECIgw
0sSGFy3XoEj4J1RtNEB8TXpDAgRvqFvhwEQmosrWWvmeZLEJLna7VHVNKVc5HHZna7rriEF0DgaK
+48MUNVv9Utfov6I2SZJzIXDiTG3GwIqYdHSqe2GuhLlxMldq+V1KmY19QxCjrz5+0xb5SH8rdN2
75WPQwkb4JdduR3F64zvs98dZ/JOUoylflQG63z6EWazyeLZgKvQcZX2xx+xpGOHTSFpYlM8pOSw
dZrBa5A6yd//kBWcb/8B6Yx4zNnTI457jc4A2nUYaF7m02NDcDqLWAMurC27BECdowN+CIGppEqP
SpoTEGl8qGNP9UAZNEfAM3bpkGI9Fw2gILijfTdMdWAh8nuKD/yheuoyku9e+ROTtO8h0L8CykoW
FDIgmFG14s/kBccRTLxhTYVS0xKsGtz/YF6Y9hIdXKCCn7/XO06kw1tGIBF6vxBD4PLSMMEmCm2J
ebi8rtKw2O5R4BjLSlFDhCmDpmq2lepruH+R9V4qFst2+a0OOG3VoESihJKIskdFcuIFUP+pOcXP
AJakFOQ7/lh6BJD8gmhZT4hU2jE/ID2HUoMCDes07hSmij72ag9L7GCwMKzGSZLJUi+IPSuFq75B
H+wH1kyVU9wRbu4/WkQsg0ip9y18dyRTfefkvMO6WSKhbxyPlpz0Twe8JKRrCnNvEK9Lr/mX/eeh
l2nc5IsZSnxwu/IRISwwix2vgYzSUAhm5a16sHI/vYEnafIFKVbGjF1gDiHPmPhQZTvoBdIVOspW
/9zPqvhW1/XWKtnq+XS/zfqRfqiHwsQv7qnR3MHUUOlWhA/90orMK9JHzR8rV/0ug8QI6yjUsCtN
/s4HZZ1Hmzwx0F3WfUMHcd8n9CHg/c1QIrNH50c/mF2KG2mJa1/vICSaQcA1cNey7NkADHN0udTB
r2Cn75qRgZ0QxyRI484WTQ0c9mkVtEwwTmmQj/E4LGa4Tw5s5ENp15xT9l52noRYMpwHaWDhtddt
0a3OYU6V041KLXWZqhnj/Z7yldI+TIck3uWoNNrIvwf467I6BbHcu8jRPSRTraqL4CnbKMsUL3iP
ug1kLPPsgGd7d4QtoadF5sbHDT1hkuasiV5v4o6+G2yXuPQcgDEq7RoL0vz8HyDZLHTDo7U6TKkh
GnIopd4AsKcwRMbt9fwBHrIeKGTUTBQQSIrElG5VMkK/j4Y9y0nQLx8cF1EdIArOQBcKfg3VoJlN
DCYrMXthzOcc+4iIJsHdU0WduGlEZHfEYkgXl0UbWJx5sXHU3xHJQlza3/Ivdjhay4F7CyX1Bq4q
uroIaHRwFjIsU29NcgR1sYUTWqV9LOz/SoLwdieb1sRD7VVJGlAsSona4tDRKGVF8nkOh+6CxpT+
CxSjejbM0ecLz/04Caj8QGQMpLa2WN6OGlZ8LDquXjiZ3Q0OZ/DOu7YV63vN4k3lYPIs4AQ2a67O
NewyJdm79nSmflnJqncrbbst+nTT/0ff3j3aYutwG6i+7QfdFTV1KWT9IFuO0Zax6j8+XssH8316
kznkJ8rv1496NBOeQ/ZC05z6EqB+W5fxYeLTD+8ZuAnXLRlhvg03ce7Y02q0cL0YgcvMbTSuGc8y
rT42R4Bl/XHdsz2QPWjoQwX8RmlJMxq/81Fb/VolMazLM7Cl0xzEE35dzJ+0hxh98rk7jft3Fqki
bcg3DzCMT/v/Dlp9w0ONczB/PnVmTwZDqO2hzvZo8rnTyLmlzb7x5bFiiKdwIi3c0Fy4cHfaeYqj
EX0xbuqpE+fhPlagWw4Z9yleGlvtAHPU5aA90fXr0jXObClXNFpsgg97Z6+E+LZ1BUixyJ4V1wZ1
OT9U0WHLC0CDcvmsKuQizgdkZgHc9/pK0FAVbCTH4yt3XbW+KEVJbjdMImlsy7SU3q3xNJ3k1ZUn
7KjWxlPIEjntTAJMsckOIUOqn+2osqc5ex+Uup298Z4ALR61+GcjnDQ5FvJplNTnnj1wel70vF02
NLYUcgRocOSpHmWsQhT+HaTkNjAPXTxkLn6fPeDQS4YJnPrXq8rhlZ4DC2cRTL3X6CjZ8eBmJ52i
XnSA2RYtnQCE/xAYVCut3NwZiWt2PRYV2cDAJDIp+5r967/2zWLKFP0/1JzU/34rgSrYaegQA88y
iZ1Z8Zr8mIqQ2Fquy5+U6OKTUtiK+hbtCZ/vqv7Ya4ToD3FYUi4g+HR/Iw3vQ5lxlRAVB1VKMIPk
Iv6mZvqflRS27BL3fKIs/PT+pzMLSmxvv6VZ8m/J8Oh8wEQKraK53Q8LHlnack51y8c8RBYi+FN0
04eUOaeEtUUecFawprxJH0TabQkQhzh4yovoGD4b8S8kBbDZeW+uvnvQRiyf99FXej6QHCQ78Jbz
4cl8vf5iUp90y+fZ2SdDjRIloontizduP8L8LeQpKiEjJqBiGdl4EAoGwD5MYBH9Lp/aXdHlY3/v
9I7xQY/usegbyARzP3DwZ00ZuvMOhVtlXLVsu0k5JTiwocul83HsGXrmPwZgKQ/AqXeGSZVX4FGk
KPLWmWR5/Zm/LggTgJJAu3EKfmCQqTxisWoXgEr6Cf+lO0R65vm+nakv2qtMYMR3e3i+qXUd9uff
ljuBBWELHIAR+wX87DFBK62+62UbQn3gdQ9ja7wZqkg4Ib4D4qHrNCTPGQ7hqtT0TUW+RLVIcnB0
qfx4Np8oB8EC3JhUp80K+oqhi/8RwW8EAKiChM4k1wzJPaFfsoUfCjIikBupJyTJaROwT67FZPof
r6NItlPkkHb8gjhcrsSrsrtC+SW+aKKiDDJHFKLe/XIeMbqxporLvqAo5RWkpNEb1IB1Oe3FI/y1
eQhYz0KGc+l8Nwm1nMoXxtATKu0D8tLyLNo32Gvv2lCxnUGLSf8+QPcq3e6KTYwif2yq2LzZbLXm
Q7DZMHZeCK9K8RMuK/byPLfSWSq8O4mWDcLstDVPXf4A6oNhEsPR/CNdroKLyKtt8c3jzZEacpOV
iGKnircNSpb3e8fq7xcv1Iz/ScS86pJYUToh+c4i4kW0QoXHfNs99NBhRuN5LS7aLp+nSHF6sOBZ
kO1gTMEHV+WsBySY10qCZzNSJw6vG5cwYm084RgFNp4WWsNSk1trRvGDTqsG1nlyukoKXh/JHLUc
5UKdqZ8f0VXP9C4uf5SrdkLQHXzsq3FL5sTmccpzmXRl34dZy+wPS+hnKgJPnZW7KPV1eLrEOmnQ
s2muajNmQ1/Q4/yuHF/4zXY9Mn/RRr4j+2K9bgR9NQry9zrpdwu1TKRt7SDjqQjd/xU2mt/3wCjH
xeM9Y1O4BoWnFQ5ylgwYbryfrFW+AbrjCOYcpDBD3JD8MWa8Bczi2MyJj2d8Sb20kJOiUq71GYu0
ZCQkA9J3nusf8zzPPW2hkcgl41Eo1uEmWM1DMvGEGdyxBN1wmgpsjEbAiumT3YSK1m50P2dmbRce
dPiLIpbIc7ONuufBO/In9gdQ6e9zIoZ6rCq9jSGX3ereU7GTHSNzzZKzvQB6LLp4GldBYeH6mf7m
HBm5LvaTio5Z3BNMrYct1d3HOU6M2DOiD3HopvIRXWkB2bMyYPjhg1sWKnj+aMOfa1XEBfqgD37N
MOpU0/PhC5/RBozh5/Cj6D9HYD/FPhyG0tloMFIarL2rACrdN9SUW+QKenXz7Tmuj91andllI24l
zcfU97nEF+sfmQIry8I+lagtt9a6CmK1LHVSFJtgS4scE/IELjwDVHb20pfX+3eYievHOyZMDWpu
GNLCbCNLggp6EN2Iw9bswJuvZf+3cX+EsJsIUZcdlCw3XwlPLNySWW8dUQvQgb49GfWcb2HsTefA
rCxYC5nAY+9BQYZq7ZE2FLytCM/YG68oSj/Wniu+2Z7zbhKsMMNUYYTEQS7RHrParwNno4d9CFgu
mLpThVs+x/GMuqDKqOVyAnCqSZh4/HFX8W7CePrinMdJ3C8qBzS0iNwn0s83JA22CBRhqvFU7ReR
JtbQTcqLeQvP8FvrZkESCcHeZLIA90VCqyBRSuJvajS1fRZ6J824FFx/0RVHFlJFwXnwtKuBokk1
D8TPncLno1SSx0vgxGOlUMzNjjlJnJexfMLG2S6H/wwICZ1em5zhxTn15biGAtQY/vKULi180R/z
WhDIArIUwQSGObOjGzY097+oMtrKE4r74WUIh1ZZIhqsn3p5Wa8tWNokzyWwE3s7uFMDebH3aZDc
5DfA1+NTXVgcxDa2yxJldHIzujyqRBeSS+e7VglVycMorz51ZtzZVKydPaBwQGB0t+jkIwSD2q8V
qnTASRsHOjIPrzIVAsg96Cav6uPZGLV+goX7ukqsIOgppEY3Rfg5cUjWAIPU4aifuTv6N1+SCJtq
LP0PlF2YZm9mjSgi7Ecjahudt9V5kd3ootNZuNHSp2i/Y5IspivvoDsR19cogYkAc6T0/PX93swU
1n/MOtQUkTYiodWicPO/vqAcLPQXr+VY3pa6ZTGI1/U/9cXrG22FwwJ4s8Y+hdV5Ne41I1K/Y0TX
wERJZMRWhF5Ki/BBmMG8fbxlPman+6F303gopL/SIqn/ThcLeiQUxyvViQZOv3gext9CMazJnBAb
7qrexvRwRWjIaFirtvaV9F4HU9UNchY1iQojNG+Gw37n+w8SNsuHYI0VnA4qXp70r1mqe0UJUeEw
s8Zz31ZTZHxf7aPR2kB7mfWXgOwZaZbUERscxxqVMiZ2jAnZaTK2lnPhYMcKFiPSmNzJwH3zYhAY
HWo/BvRvTAsJBrDMFvJIOfC+ROjUn73pxT5Fou6Hax415q0QgsNi65nPCfedIhbSNr4v71p4EvWr
c5lHwn+70EHb6aOfiwYZbzz11pIYD/XR5qMcabUlyy4GYuAnvmqlqaP0IbWBvqsFZXV24K2SZkfV
YvEk54b7aKRYXDYpVuOIIFRxZj3vGFjomnY4JlspnuylxzHR+WW8cC/yntbovz/ytnwt+NyjiD1N
kol93q/zfiejuJWdU7oy0vNHKKVDMKcvoCfyr69jKjcrV5kF0HSr+9m8wba+vPcfHE+M9v9fgsBX
cDfPwSCcENby97WdPRi4q55Mt4COqglUBvuEpk7trBqToR0OlRmH5P5yOE9SyL0tRdoPLCb0Mrqn
aP21krM1j7GDfT5GUi1h+RQ+fVNzHK2C4Bs9LREOAbJZoI3qpR1J2z2HZuuWeBxy9pb/ekBrwrRm
Ro2RregpaSjhV+EK3Xw0r/y4hxIe+/Rb0tcDNhSHyNcDvV2D7531eitLquaXrEkKp/K3hiV/FTT4
KdM4AauDZBwfUtRt9lhV3BcO3WOL0YDNfPZ0zF0soPdmTp9H6z+QyXmLuyJ2hrdmtnucSIGtNRa0
e2H/0GT1bdvTubYoXB5e+XGvydisBn/xgY49Wa+jCydEzjU9ET8mX+S29GEYWWJLSGsmy6o3AnbD
y6uuENapF/vxcXsezM3xHSKPjseYNm2fxXpM5MTxG2VKsOYj1oxcLrgRjFOYznYPc0RmzWPNw/JJ
Lfpto9fqSoj4fT37zIse8RmbH8gOq8kOHkQOPgvsxNj6E1+MyoVHKcg6NwqyweBqKW9u53JgBhzf
LHnksYeLZ/zy8GdnDC7O1vOF2dT0+Srwc/ov1HaGsgWHRw+CCP5JaF2xsIMEU65Nj/g5RRI9y4rP
7tdZIb90U9DMhCI7OTwDoa0NyvisTx4cGA8iRRlQRJ7oeMS0bskBpNOoGi9ejnez8IasBT4HjcfA
nz0+hqPRAjH8RtZinW+SVMgt5Z70As4d0DeCxLIx+Q2/Z3hgzZejEn8AZx6JOIf3e1C41Mn2va9e
/hSVjMYMyFUNfYUwWyh9S+JMwFDdhgoJCatoVDJzzNcxpi5u70mts9D5xlLs+6bzR8qNVzMs8UqR
doRdo2PaLV+ZsV2DdTpAQ6iUtDCit1xBW7XJXD8QpAQ2dkPm5dx88JkmnhHZdCHCMXG3h92MVs2N
of+Ht3OH77A1tZnM9Oo2fZ3/RwLKa+GvVbfEBaYvIQelh2FCwjl9zMqSwPi6SvsVmh8hi+OtUiFA
+O1uMc7lfmfRWzdZZPr+GWA9WQCxavUiy0pXlrrGBZ/T6eTO+m/p5U3YXNw5/e9S/CesH+GZf8FG
Fg74f3U+bZr+gLynL5T2bbJp/hRw4Kn/LMqFWi3L77QHM19Ms/c/4f5iXOi/St6bfVEBm1xjerm/
zTb4xZ3tegG+3nW8sQ1UFoH/xxchRk1cvQFEu8Xn40Q+1WmYOanpIGIS4ERKNXo6ntlOW2AXvtU4
4ke+GgwfxC5Ph8cT5Q70r8zLWVIl5mOWbJNNsiZYendXxdH68l9zKgAHh7b1OVEG1SaWDa4AfVPg
9njWXii4N/vX7YWEHWPFGpqyysV//qzvKAdka/0d99X3ZOGZPhk8ezBnPjMLYix7KbFGx2BWP6fy
njGVA6tvTkeSAYsrR4GFCGgO/Qz7cwvZVdqxJOh1GA/xMXuGlS7NN3ZSv9WMFVz+g7/DlSi0ioZd
urtoE/5ypUNL0V0+jsoeWULaqQHzFVvj9e2NHrNKdHAyHQRHe9h9n6QWTfhXQeCkzgNk/XA1dm5u
ArobM5qlSf8/Bw6HRh3iBmGc28Ixx4xWJBcP41VvnSleXMnXV1aBJ1Ze2ya+OV4DyFPgzsKTZ/kI
jsT0Mt/mf+2HZvqhSbxuinAN7wCH0VTVDV+mMPZdVHyTMHM4E4ylslUAwZPyaN2KB2lXEPXu4sR+
RNzeYg9W82Hc1se28h2OPxIK65+ChIUs8ujnVJzKOuBGyCIxDOqQMFqXUmaJcubguNtD1ye5aDVt
HE46OhFIS4cyW6b86kWesn2226xOppCP8sc25B1vMOHDhBVuEorfb0Rcsi9gk5aJEZybnQFJrxlk
T3kxR/r3rAX+hLZn3ySBBEF6aE3E9ixbUbHeoccnBsTGKGUqqVdjNzM+4WkhX2mVIFzwGesSeeHs
mbQyBW4soYLEUXgSRGVMGPnLUYsCP1xu59EvnS2t79iYnVmjP1lKJf+7UQEr4hQmrLnUS2FYg+mm
dmXulcW6M4BYaEYj76n9ZFPBCdHcXoAo7UF0juj+Kr03hU22L09kCJtqvdRQZehpoNlXmGeiMDxp
ltltb/BZn9iY/GjK/tpdSIgmzp/LTL5r9vkPK4Y9+8e0A1x19YitvrhmEcxapNcW0+GI4ceJa87n
3XIwSZpfETOJaF62ngzT4mevccUcBtEC1DTyJIYGIRNRDShNVOnZViw8+4rchrfu/9cbGsJ4fjhH
gpB1nAtjImdi0KmxUgq42rqJvuP8O1ix3PcT0elxx5Ks9TJXo+9j0EmucCu1EzHNuboqSTPQJ1V3
aab9Hwi7JDW7ytZQYx/kuyIeexW2GIl0qx3stQtO9NVy+pp/ty1hBT5d0JHTYB2xh3Xw/DiyZhN7
twsqlJEVBAn6TJ5yZ5xkh5Yji9GSc3h5Y/HLE1sLUpFaIVBG6IU3M8RmTVBzr9ealxBsHnlEQWuk
bYK7TGZB6rceYuK2OfFfOA3iWedX6cGyOuOBuoA9x83XmpHpgVqcO71kk6431Sz7aMvMtSckBR2q
Lbw2wZHfQasDpH8dKGbJFdm704/+5PPcbOUZh4KPT5SiXNl0GL1Qu2jTanbmM79AYmPj4/59wxXF
h4s4hBckacB1IexPEiKr7ZNYP26gdHECfZF74mOTf38njeKS/NLmAtoo2rICab7ZDgVpFIvXqvmJ
290WO9jOiDuq5bMsLXh1v0SdRM4dZdlgv2YYKLBtjKx2h2BZmfBbrBcev3V4avoi/y9lYmtVLsiA
248pAPQLB5SXtmTri5nwJZ+tMCiAzOsg/bF1OCI8H2HoiaJ4YlgVBJf7EV3PgzQeuS3plur0zqOz
ATbPhEIfwKx7YN4QLWYrveiVLqXhxb/KVb6CPinyq1jne0NheHV+e8ai2GriBG7woak5xm1cQNKJ
XqSrkOGtygS5ZiGs0aRRT0XvlLX9BB1DZpLWVq5wOeZ2kLxOqxqqdrfSTxQMAKeIaIKCPjhMOU2a
PruilS00041zApr+XqqWxvRDKB90uPpcmnZM9n4dK9IZnpWhuN8l6/MNnn3ol1TJCnxSclRtXkS3
0izcc67k3AF4WPRy9/Uv1xekEf0Zgg2Uu7aH11I8fftZIMyEYYdEPcuGDjtCs2dOgCYDpzvwUTRi
rxPqBL4OQpEk2KiKTmK98nbazSeLbdkDQjvNb+e1IZG3I6WJLvtSp/YvAn4qLZ2AXkc200pMzjo8
nE2f4p7PRwVMVch428hGAHG9um/DNrhiZeJNbR5vbbYBzhwgV2PTUzustJJYFVSuFfsACAvESWcr
TfasjKDQvCzHbj041IH1zoAy9VFO5EAmYGj8Uv2i2S9Cr+FCtjkdra0mpf8DXHU4UVST3pgIJrfe
59ag8DzZlrgwhycNU6l3IChITUNKj+luSu2YAcMBcNgZqjzmz2n4nxcHcpFF8JYVCN1NquSGAvoT
y0empzrclWjbEnZeKLATfp8TPn4DkUatuCnIGS9S0a1FWRNwGNmy3pa9MdN3tmk+pcZKxd2IBofF
dHwoZUPz0E352U1jbB1dLxY6Pks8DPMEbuLfOqD15vO4K4cLYYeOm8g1nKHKPOwhEVzW2faewQOP
zrR5rb1vegY8FgUnWxGxCraDUp8VlzXnluKUFl8U6Xd3P6b6y4hZvtkPXFnOrxC5eJLfc7PfsXnx
hwbz9Rzz6LDLl4dtRZVD5cIrNJmb4sFJx6NqlL8q2P7LI4Q8kEQNH2Zsacz4GsJDthx7b1iuwufA
qZVal+Sou2opjypZacOAceGHdpHnawZ1R6UzQdaoK27p7VhfZO0M1pBeFW0hFh8gAo4yo5CCuLD8
ygTL/I7hgKzGEY7uieG8+rmc+9cH3P8Asppepr+UnDMNGfrEOCJD501ycgoO61Q3+zEVQwWCGgu+
YzSq6NTu7p5HdtgNOMrgxrLXgMSgBCLZk2LpATKg8fUo23w2+28AqaZ0ofO2AJWENyllNw6Eh/70
W3rv2wPw/cvrtmDWPrzA4eUUpP0YwA9IeT6kGyZoSNhSdlVB+VdheVXNuRYfU+vXNRvX5qIlc4Vz
f2M0L+R9WItR9CzoRq/bNvN2JO482PHcYKTFyYpKTuA6+eakVBk7qNd3/AZBZH2CkB6L8eTxP8nY
/4ULnt+Ru53i209SqALvCNQolkp+HOimcpVHVDryjLYGLWwOVHQgKaqcG99hABj81zhtbwJaGxSX
E/gcsqxBxs6GgvBq+8+UdpG1SFxkJJp8oAOCEzEcu7b0TWZT8IYrxxOMu9AKIm4YPgFmgb9bTAKb
0NwZBEPEdNuvR/WB3GDbNiAZuDOlmXoLSIwWMYxYd+hs0eKPJ9vamkU+6YilGemhOXaqE9WvCM/H
fAyID+ZjTN5tooXktN8tj4sgGmutRjNTW+6m5jjyM6puJZhS0ddfZj8oqQputuGlHO185RNN5rLd
L1SuC8Zz9ZDRLHDmGY3E3cobj/Sl0DEsphnZdEjP5lAv1A+ZjWljKRe7xgXw1ai8tD5p2pDk/Kuv
WszOtfoc62wV7KW8n8+t3CdmWihmFSa5XsgkRrm3aC2ncAfb/ZzGV6bVkrrY+SX3Qk6PBLLQ5avJ
xX2O5OPfwEGmNJWSDvG4MY09rC8p/O3m6YdatUZQjLR18PHRqT4AFjf+Mwvcx6jYlTXcpXzV5BYN
obxml6CY9i7MoyMeF/xRoMp3h5Xik+al3fiNXRMhM4QSwW4FIx3wcmn+Hkl3BEU7PC0Hf/iWEZKx
kIdAyRhNebXgEgoBbAQW6fPN2qpRhMsWyf5i9+AVHc00xMWJ81rEXFRTfPkBCZrTqPj/dhA1CtCX
Gc0167Ew533vBj20XOapp+X8rd39Lk+nz7lw8YTP4kMTZXoWn8RpzzjBPX6ye3lT6mRJunOe0sR+
AY5VUVhpm+azkJvuE2cX5OpOYyKwu1e/xeCfRsG/Mw57x7Nt28QXw7YrlO8WsbUb+G9JbhOMtQuA
vSk7AsuVhnxQCt/5T91lZ4JD+3exGlCT9nRD3j4thtSBj8lKogE1LWwT+SkR7pQc11HOQXHGpM2y
qFqM+0sH88vzi+dw8I7E6PAocwby+r3kHwKTsT1V8dqZ+0+/vv9Tr82Lmc1wI5pV/44RCCby/oyT
HqapTDovIUnFYBiEViC14x6WTvsvin+gy9eP31zfBHzTnvmeyu7/Wz3uDWE8z8cx3/e3+WVavVe6
jO0ypRpJVwhvsJLJTN7CH2gd0/BjpyPf+Dz92w80WM9r6IUhhV+vhUW88nE0nFg8RQ8xQV00wak1
3ZZEzKVAtnilpSyLeGbiXTwS9lZ1Btwtm4+qcIjV1OYQMkGIa1Et8lNO3BKB16fwMRmpX7soFoud
Nu5ttdnNCT4uEDFndDtOxQXUdnZvOGn2b3+7AcSDfC2rMojEchBIXHYgyeHArL12klWofKxH1hhr
XXmICV3qVKd20SDfqNRWTOz6To6y7j/NGMV2z8KNvV7uOkzlco8PaBJuDRf/xz1hv7V9bAGwjAvb
XuxKznx9YWgAw69HoMvdr94puegU+hhdhoXYg24b6A0J5zq/1Btf5bkOxqJsMMVpspQQuCQ0Cgww
0qYLV9mupVfQ7wpBWhWUoGEVQqg3o1z2vh1BgNP3NUrzKZEdeqDLcmI9xdsMn2rF6cBTlClDUvGA
l1eIQgZ5zkm3UEOP892G3DZlf4Zzqkh7bQRZVDB4iABOucebm+88Ghc3L6Ibe+XSBfXPodoFYM7M
uvaCyYRe1OzH2EtdDpd//l77+4/64lx6H/Ax5W9rOxUt0h3PgIRWZc5WQVgjSVP1XsirV2nBGQTT
RoganQP69c8UeQvabQTKj5AD/MdYp1ep9RHwVKl3O0+mGVzzeo7/GQExb3e08T4bFnrdK6hIIaIx
0gr6St3nPpnReOw1jTIuOyHIXY+tuWs1kFhzK+JzVG6t2/qhG8Z6UQHtA4uVtTReXE3kfmbexwde
9SLK2WSCeEf00th8nuB7sn6S07rwXfV8P71Pp+XEpQF52XEElXdOLETO05mhZPERVknQNKIvnKKj
Mo4ACV4nV4dAM6MIyx3nfJth12Pg0+NsyF+9WZpmlMX6xbD3fyoTKdWx6TNyWWgcTzlrjo9V7agZ
Z2aNmTRa7CfKQHH96fFNTrcqjfV3H8Qu/FNiqb4kC4EYlgQxyDEI0tgos7pmHTZQ9yZ0YDgHW6i2
8YN1CTZ7UMFKJYt7lBBl/i8qhfcaEjerJuVwgmc65MFCTEMDSBLWqAQ4JeaPHnADI0oRsnJZG547
k/sKXamyBLu8SMcy106+sO5Mbhdo8SBJpBb2OkGjFQrbKC9/ei0stop+9zUWS/q6tNVptC4OoGnT
3oAkIrOhCbtywjlw+tWazEA3eHRVcnxeZv/zmndZMVjO8OqmjOYABPEYTREa4+Zlw5jBhiF7HdIW
lpMHc33gP8ia+MA+zJCoup68KVPMTJgQUUhBRXPFO20t4OIIPBsnpKtSA/NONPB7ogkFus1RIQ1M
M1BRCR8J3gZbfday4qPij6y9BAYxt3g4yhdTOx9oPiG+r3edJCRrx3Kv+oCx4ZwIeJTgra9rtvMd
EggztfOX55mRqAp4GWAZ3m60Q4WwdQ3kg9AnQ+pqZmailb0WEeHbaZxKbPRFrl0M7gnNGSl0cvaJ
H2hdxFSYRm7Zx2qKmmr+jzKJ8lCsBO+XwmRzmKHm6z3nozWDy7pRRzq92vvHvVW3lg9NZNstFAsj
YFVnRtdLezZlyv3gy2VVJiBAmPHantnR9H+W9VTa9uGPKgVFanmuAsg3LxoYdCsznDow6ZZow1WW
z7b+5NnPDxG7w4kQrTt6fANrdJj4vx5i4VPHBi92C7B2AyGILijz4i87fRlJd9RWIjwBEzgS4pSz
8qNuWJroYLdIlFnVAmjkSUncbnISgTKXrZKWeOvo8YDt/74F3vvVVIDPPZXgqVqrzQ49NloP30BH
3HLl5KhhHwEq0mb0TSATVx+OOpU007LmR4mqBW+wkQDXOiL6D7CROMqWX2SUPNN7p5fDUV7MrmyK
NHpy++iH1cZ2c8iA0m8wzd9NjQHDvxsihGbDzyvlGcCpG7wMcnL0l1e5LrKHSfYjpJOs7p/61PIC
U7qSOdjwjnKvHmB6pBxpA/UTZSuf+3NJahOlF/D6+jFk2uKY6g5LEaBJCaOzI7rDySbWNL/P7/Qe
MnITokiQS8rumMyC9RczrmOJg/3JzikLrsSebNxuNJahzIRbKUj7ysRMf4usQOBH5FWwhF/gFjiK
8byH9bqpZeizlDPg5Deojj4LcxBgU7IMr8ma05r5KB7o+Nl0KNyJST1FamvT9nLhldbL8G8V67x6
ygXVc++lc0IDxXUY1roD3wSZHIIi14o0KSQN9Hh9GnTcTfLiaknXRKhL8Z0DCklgxq2D7RqbByRt
cz2+F3E3H0yy7GVoWaaPkcQjFNLzryjDhsPGImw0ugw2vQ0T1GWnt/Ze4KhgxhO4ap921mhDyt2o
uqnL+F2N7/ZfinrOAY+ReIKr+/qbtPArd8A85/3vp7YswR84iAOsMXgFLpfLGV1F3gxdnXjY579o
KZgOfEGDxGUtzFoLLROwpZCQNcCHRHS5AKGqsdmcczKoGsNWx+ojq6bB2H61Pg70bZ12K48j6QEe
wNuo6sbTfzCBJ92BR9kmR/crVOCrdYgC9NX+k9bx7FXY8kpZuH0+E/OFTAzhbjhcmYiVMnzE6pbC
wrWqH+v6NtUXn+F/XIGNbYpa08W1igo7Qk23igcBwr0uL8g58dYlfa0JWwJyu1ttnibYWiGn6vuN
jBXwDnFcgxDTtOmUBt4Jt4XpNYXZcEjXHYWOlWXGlC7pJevwk7DTOqmLiynA86jzfN/8UBA0CXIg
yvf5bOI1NiETdLgO5O2MOD4StCrjWidX+k2HWrfpM/jLZQJhgnoToPJkO7oEukhczhnwaEFv0HA6
joFjRwGWyvD7e/7njQ1vu82lJXQxq6sXmz8qXfn0mGYvSKyiprGHPRHRKKu71TqBLJPfyKTV6WuW
uAQ9cWTn25Uq/B18wE7904qhZjJB4URafrdmFMK2wxP+RN3I4wciEHvyCXJitBu52OMnX/SrxcGq
Abgb5yFc+RO8yKQ2C15/FgJHzyd2jYnnmuZkgdmc6qLIsPPwCQ3gmu2/s4Bk/NwjkDxb9cR2gt/m
4894/+cCGzYcgVO1hgOjdWl1Rq0Zs645EpNiPqZllC4hGAPPsT4NlyRXsllAZjCoNm0T3a90011Y
WAp6P0PbtczS7phehH7WO2cilx/XuUnuvF3wqVy0ImeYHSXcPawYboovRVirTLd0VFtyqq8bjmLk
ekeve8MwFvEZhxe+UoSf4+ZIykR3WUrBqUJIbUwJjTfLVHeDONcw6XHx/cB/JKSPh3fhbW7dN9nZ
ehAdlxWAm29rlz8iw5J1FuDEIe0KB1dbozNB2gn010bSxJaPg9D9ipcOUvBHx2Xl8/a11xU+Jx5m
95M71cQTyyQutDbB/5Iso4b8+tR2nOEGADJoBaxKqSj/jMebsjW/z1y4Jo75lBALhzc3gXKSRV+4
758xpY5tXNolxx1+hCloT89bbFm0UaXbyZnigQGjFBeIWHduttvexIRaunjkajqxzxB/xi6V7fIP
ABeywRWV8wWgIuKQ7OS72rjrTi+XGXCQkMSeJtpZxOXhQQXL9nW/aKRP4jDhTi5Q+AGPr25EnVDO
oCFiVoI7kTpd9VUNhlXGgepfgpPKQIuauLKln/izjk5Wy3su+SKUMApJ5AHLp91YlbVUzBIyyXc2
ZtpX9ACXhjH75ZVQhUvGPlYicG8upjJ0h0rrI3yErPMnQYfzFU3OWREc9sGurWRXRNBu1e3j5Kzk
Cy9za1h0aNk3UbjHvCVKBY18U+UMrkvu8kVy6gx1rzgLkpk7wIY+3JOlbN62G7KYYw/Z9Nk7ln7F
yELjYwRT+GdFlFDXVNBoXzBQZm/w/nrPEG0Qkxtpi13Q8UeyzL2lEryoXsf3jWb5Dz8DksKZyVGk
QjA9+dr/HC3zXWcxPiWW1Kitg9oI8dbThc5uKin2I5P0JHWRi/zMSL38Mr++bDHHltp7aYNyGwKK
BmzpHnwP2CVQ2OoU6wTFprvsBRSwb92fZ7Soq1pBgTYLad4yFWnqs10NyHWcfFlM5wCxPbE1Qwt2
sf7MMNKFG3BqGSr15qplSvMlJfRl9/VgzVtV9J1ShbcY11vrczfe/KyC1xCkQoKw83af3Yz4+KZ8
T+BzhCiSKEgyWhIp6qNPrr2pCXvrV7HQ1Le+/ECV7DW4WcAYXFu97TNheZ5C62LMjtBY1paiopxg
QJD/JQJWp5MhlPmxVkmmRQg7qKsQJtuEORavzF3I/6RCqtzUvRE4hxGbg6VOreafu0qdOhnbVB43
aA4GpRm8ot72o4Sg0U2K++I7LU48Gc1S9gxeM73ly9HzcuC+9oKnRbubs+mYjXiwqyFxWuMnNRiF
gnwzFxF24vySek7by3ZTQCX9Ay6YwybGMDDN33wTYC+DziRjLflfdkdUN3Wo/uPEtMjwitO1Baa3
B9G7mnCuJanjdJ0IAXlmKZJUbDMWTfMcBtRIBVlc43S4sZA292wPxSjSF+kvgBUOdzVM1j2ptMCj
JObVUAlM9C6Yvr34zYkwmT7GPnd0R5DqnJ0Owf2YKIOppxKv7FwsfHW2bBec6jISztO8dLTSWWW9
Hl4ADfYj/ZPz35HxLphlwWln5xZWc97Bnc9Qbh1qfgWs+KLzPJCA1nqPAqt8q8zcxly0/LG1/pR+
ev/Ex+eKQQabUa9FInRZDYFEpDs68iCrwRL82uzKba3c+0GuNXJUd5hSh9ve9aHmssyEa54EUlhd
kMTP9hVZ90sOVEpmEJScVEx43Z+zPLgCaFiCQVDW3a4LxC/KzVs4XkKTlL0gOpJ0ltuYicUKKlU7
+4fIHVuBy8wFICxp6YY5Ml1jf2HrQwhRZZxV9XenhmrRQGqCJF+NSlTDUJJpGTmuI+vuDUTzM9yk
c+Cg1HiuGsp/WAh8SF/a2pTtCasgjSOAQwf4+DdB7zK2EVHV8hEchu2DANbG1xwGmxu7cR+M/4kA
c6sqpGi7ithif0G16+akzzJVYBRSY7KEFWMj5y9WnKx5XM8Scbr2CjSw2G3bXU/HsB1QqQ68KUkd
UxgIP/zaAiu4AOqAiRxZeRxfFi8iBIPkfbbAI6yI2qZ201Fx3mLJaZbSCQmjVJ2IrMw4SeRoHl+b
R5PdMWsSha6v/2t6tlFGSyog3M371EyNPHMo6w6ZF2YBreV4Rf64x/JUaUIOpssMCuLEQ6WMYone
x3Wy593YAzx3MuCCqeELBey0fFGuonI6R5/cV7AWfzOiINpKjRv6aWyRCifbsfZpnJrQmmtGJMnT
lbyEcLbuOuZXLE8BwkkQW993rOtA1azdxbwE8gRyi/9vM0NysKcmC+tJYa54Wxy/8Uu5uMoG/tTN
qA7YQhFUdllmEaUe8EYDNZe5hCbFYCEt/iDikPCox0KPfdFL1yTHBe5bQLOIt/7xDQtcM8eFn5Tl
zHKDg+DqCRn7jVfg++Iebpi8lxFYFucEdfK8QsI7WnDOM12amBnMfG8JOv2LHbDCf1DVI9AOt44K
RwqriKyIhx3/trARF1Tb2Quvr+wmZbfVXI/z3JGrwi7MSdNr9I49XGmps5fK5Eq4ivoBMaCriv79
YEvYRilYwsbmfhchkJYIWHO9znO0idRTAxhv2ZKGoOxbfjnFOa/rJDnbf7FdNvUxU6c3MUIsAe9a
oZMBnps/Fzn7UoSZ2/oAdcnwO+OvueeJlXLav48l8CWaetemGhhMW6Z9jdww+IWhjuR7xaBWeLNj
Ct6Oss0/yjlPC3XSYMQcZsXjlyEWLj42MP2wFKJ6NlhueeBZiRTrm0gBMk3mnXeqHcJ5r9uVejKv
etkR4ww4EqdaQwSkA9Sr7QnD/qW6iHumsNichfh67m8Ev8nYKsYID3tv1hy/DbGec+1mctgPSQ0S
ZezJ/HpqZkBksdXzgmJQ1OEuo3ZgQWHucNxg8trnAflu3b0sW6DxJ1esVeg6w/bHuaV1btrsH3tw
eLLn7biuNU5eMwYOlfYkYzQF+tISsyyTanEQmsK95ozFRoBfkv8JHfwDlOBD7Hs8cNCDTjvQLU6l
P+Ph+DRd6yzRvY7cbxU+o/p0gQHVztBGtm2b83KOVQejKo+v/Vlx+mpaZoIBDwF8Ouif/Sc7I27t
pSPoZaMbZRUkeLStOj4AU5IrWEF37eocpxtiEbnD7+N5uPJM+DPMuKFbw3SxxbblPO9MnIY6S31z
CzRTECMdCsFl8SXtAOoD8lYgJ9uAIAo+RmhRNNU0slUfhj4mVC9fqMJTv5FrBJbidNWMoy0nTFsp
kayktom9Ef3Xsv2nNGmElayvKfLp8dtMGIYWigX2qACVP/vsM1KaZpu2JVQoUYhajendY6T7Vknl
gjnq9VkWnhXkpMxccMA3oc9tJkdE+oEcopR765uZMzWKxOqCsGK84EWtexurIwHt9J/hcmXQRPrp
UeTzy9owCQtNe+U9/NKILfGNZAOHl04XwqSE9ijKBBPHrxcZ+qbL0fiUpXnfq9OqDwHZwOzXsl5M
bXHFL9y3N5bWsVb9i78qU0ROuGjVidQ1AtqjXHShuDzN0lil1UI029VjLgSZhmC/B0shmS8GTb6K
XLyDnFSjZ/3KBLOYyKfp8yWMj9DynnFCrCdZqe7cO7gY6ZiUXxUpHuteQ+RDOx44Jc7RVcDGnoN8
gjXE+2Va0wm5ta5Bsz3fOW5TgMVZIg9RiwhYuHAeZ3v0XUuo6rlnJJcEZmmjA+r3HLqgJUg+75Cw
bs5VuObM+Ot2kYZEIvXkAQ8+q2zv883zSnM88M91PXf+Sw60j8uZ8WBXz7GiVFxui7HetyTQRgb4
AQ0ozU1DSzowksvHcW+tA/wG1DrVDybnfcTDewzbIpxKoD+aCNOikM56xgjIEnuGxIU3WPs3gmBG
oQL3elXxEyR3YuOCpMJqKxKZEUg3eOA8++Uhwu4KIk9ins503CdsFqAZKY5WxQroXVai7kPepAvB
i3Lap7cqf8FlD9+Z23L7O1xitYlIqJ5gXMnDof8yW9BX2qhsx197A5U7P6BLJZFVt+g+GkIKw1no
C6lXDD702KzI5K5dpTHMXgVeqNDUoyXM89huk2BsMCtenNRNia3LMaTe3h0+65TU/4fo/Qa1Pu0g
2DR+J83ABLzqrIbKIm/EgVHNg9zoYuya/WRW76PIAls3SQ1YTMGDRYgdf62ICD9tbyAtmaWj2VzR
OZnwq5/DX3IXSCRzTEb/2So4AnexeHEp6aozRveCu8m0Q96PWqdumnaoksY1uDW2JnqsL6yzZryu
lbKDPQNywd32AT6Pm1kILz4MnTnIxM+Laxmod4e9ClRD05Md2vevPm65zrDTeXIq+pEZqLNz7q7+
3RrdRCmAEo+DKzJHVVA54vM1uKkcEM5XsM+YIHcSQ2KPA+NNhIHldyydBD/yqkEk4hmZ7iLwg0xy
zbZEA+b7SvhXRkA3bSEC3UhRIweElxHCPnfq2pp1SY66YPAfAUCIQqVhd9QzjsATm+1Ba301dLF0
x7DuzqcJnOsCsnSC8ctyIAaIHzMEzUtRGFlWJ8bxVb1XzLA8l0glZRdCQW0PAuLebDhsoG2X15U7
34rK/DmOwuwy3LWX8glIv+Vt5i7+eIzlROJA/i7j/x0r5f1/8/WbEt/0si87bYRV5oCNWVeR+2iw
emRiirSa4paNXLOGbQ67/sPQ3idUH4t+WGxG7n1eUAcnRpm2I27weojysZ1GfJoqljpT8IwlDMpS
QMUTBkOuPefq4R/ZenRxWQhKzHmgd4D+czasSNshCXBJrJ6dp806945lJ4in6Sj9zTrjGDyXI0/F
qqKj0j31/aN5xR70uy3Z5hm2494riOwYvdf//02fH1OZ/23E5XRAMd5Fy1cz8H8qoMjmse7Xw8gX
wfYCVSYZ8533Zn3CXEdiW43CVW/BDhj6q1Gja+1rc/Quc77fHm9tQO20nmHMxMzNl4R9YH7E/nfr
xTJpWWGA4670sdgeTS9bmUBr9abXDh68ygilf4R5cUdqB9ntHQAwE6TPhCblaHxB6AAkFv4pBQRl
YGpyyiiCXyUyZugnV2Ipmj3RjSIqpAdXevngR6Rf/dCUDY9U6cSEeQGRaMv4vUxUwTgDvLTl4f9M
ztFZ511AQuWmTRSVBqHsJPP6cOrDwRtXsWloNPDufGSh4w9cTtmpSubGimHawzs3Lmf1B2cEUO0j
pwWfuKuNGF05OQRxSpbvCLBte1vibo9e7TxHIKbAXWDT/TTWbfUPlHscjRN5I4/WMEBWrvpfAM92
Bo1L8YRQa/2l+iMU0TTfi/3UGgLN/JLFYuFd82CrAJffx3c3xO4124uPyVYdpcGOIkUQrBagLg1v
JgL2Axrf8IyeyQolBRsfcK4P72UlO0GKlAjnDsRer0KlENYD1iHNIaRWPZ71026bdkx6ZLxAYrIQ
nOwKSbji7ynPU+aoOpXihl0zApOYcTbMmnJ8Nri7IxDeT5EZsDY9gvOLQT9eq5Joup24oOQC559O
PImaE/gzUKj/C43JG93O1QVKShVYLkxg5g4/CE4RoAHuEZU5j4IrIoDoejX/pisKnXIRiCPcFksw
nHr6vzXqzLI9gyG8t6xhVyn5bf9Ul8RbNfU3vuohet63X75LnTrmLiDLrSWtvnCFlA6njwXOl3nc
YCWQJPjnAqXUprN0y995ftF0PHPMu+nESPn8DlzA9cCAiMoJqG/IHE5eUwgOp3MBp2OEjkHopf2P
XCKIAciEjyTafOy81HrjovzSTTBa4qTIFmCi36lsbgJzKpBsYeVKcsULEf5i9Kt03wj8tl5DANqO
6ikfuivu0MPXr9PE7gPEpAk5KtxOpY6iQ5rwzkUSITc12s/c3UTw5hlV0MqcXgIv7dkJhlnb2e+v
OsEVubZXylDcETg49loWcMhB21Ed/Js+E3bN/J7hTXB567y9Z7Zd0QUAcKox/xou2c7kUJukL/PR
X/4uWpTVtWfLUKMMadyslhUpELrFSy3519RnTgGpBtFHIcUWdNJZB68nAf49BrlHRdVRBF9CTghA
BAVeoCLWRFobPUAgtYMLWoVPXIDKFKqMQldfRmdhI4sYzHdEfDChYJcY/fsecNe4zUjGkgQamd1U
FFYO0ifewZ/N4re1tHPZ7LIoWtdvgtKRHqLACjmrisJNK6ZdfWhtfO5ajVz6iF/Qf60C4iMX7wnr
Fd8mPJ/VTmFFUjudgUjjHQvvw/2dATN8yxqex1JKlmRRlYslFORHh+f9+2jzjImZ4lQx3kVa3/3v
HIue3VijWjboslYJKh7cYFgY+eqx3R9erPyzSb+0z2q4iqkXLQKMjpnAwidKme9ihTaUxqAbBP+E
s5veSrcN6zj1MW/hUQ6vhpoSVzzmLM2lQTcjMb2HTvGCJY6TbuWeoB/8edHqF31nC7R7lk4sdpCE
+FcU7mm2KIFkFX9/RDA7pShMk8yjF4zLYAZWKRy4+3FskDOFB1OvTN9M9Ha53ObLIJ5ew/F2qzJh
lpxs2yAlDZ+BPhqZInQXkV6Smz9X1t/8UaKS6jYXcgeu71sZat3NXVN7TWvCCZDwa6L79k+FM37d
qQttx/cyL1P2TYeC8rVRVKcLdwz+oSXjvA+cAu+BpXBNFik6/+cAebkbP8dCE/djPBGr/ku3PAVu
prrjEf4FhSRF5fEt4+nD0OImdwGpR5bopHHbQlEUGtrz6iw8gh91JjQ3ftxp69c4wZf/ystLwAjA
TJ5c8e/ZFjtSkqGA/ynOlNqwdGyaN5vBDTUCKvsO8TXnQDW0O/q69DxVqkV/f7hUkiTZDMN6u0wd
f9VV3u4nIYoFvVMIgETwmdRzHkUYGr5ETTZ9AeWQgAWu83mpf0YY4bSxO61trvU7NGErG3Q2OYgg
cNf0TxDng1Q5g5E39RM9vgLMpXSDB17uBdWjPMioVGDVO26XoPUXTH89DEgmcmOcP1TIxP1CnddE
4316AaD/ES6XtchmmCM4rTCJWD48p2qqnU0LwBEqSbJTdNacdiU9Kdzlu+rUpZhLoXNfr6U07Lsd
7pLVvfYsMyXjbjt8iACrzbNWQ3R87DipP7JkOGzPzap8YkPZHEqzUuG3baEEIqnMvfSdiPD6Z1Wt
UMXMcBIIdbDhDBMt0j1ysTUQQj9Jl6XF/QOfYD0447k5N29QPkGlLnBq+/GFWLSSYcVj4ayZeWf0
PtCbsNdv2iExkKHZXXxdXX8Qnw7XfJNgrs1qR51QDdJosRalj+oAcYUfVnbcob5kmQzMY7K7cZM+
tyAZ+/S78TGqoF62BveLL1U7oYUaut8S/MkxT61zvY4U30HYAKlkyfot3YOXiaIAprWYvrcYXXyf
26sehsOy56i8WXJJqGWts9GrjnpMOmQ86ZTuuKxRb79VanVPOqeynuaR/os8G5+Z+UxMl6WU6PIb
UsYJQClR5oT1+bOJSAQ+/ujwGb/dZ+BNcXSCujO33swKIzj7ZcDJ8izajf3SPvGUg0GAITzFmsEz
79cyi1GVyiMUHS0IjhMwllIP0PuRsLoXGXXdtRbwhvdNIICtA8hr8Lc/jgHrkF5i5nz6yBtQIcsX
HU5Zc4MbdfnA3d4zEYWSnnSJO2z8r/hZSknmdAquUnwBE9X0NFCNBUAEc5004pEGAMf8qXS+k/Sm
a/85pz5pxk9FaqIv8FlbMOdyLCqNBCWX+fH544qdJuGf2WDEW7fyI9YvnPNovyiluG6gTSEQhmn2
9WyacQNx2H6YLOaPo6AVUFVmn9m+JEvBgaqT0k5fC+xpdhZl/PIVRKYl+LNSDv+U9j4mczhK21nB
AODZh7tNJbtT2RgFIYSrayT7iBT8lROuONSlUqhPrUpE8Pn30PI6qxl2TjH5Ns4kEe6z7LhC48VH
EeBtxNXCvGu2oB3vLseeeT4vBxdvaxfOq5PBrtN3pLbfNm50yI58cRXu97RSFvlU8mT4ciGHcxEi
6ae7EXRNujxPDeXsW92/wmNUhklPd8Fe53K5f0BN5t1ZMcUTxVqUQ7DGs8Q6IjBd2zqtniTkRXaJ
YOfaccaTa4+BkL1WJbVgdPYCm2RcO1P0YQWyhVHmJVoA27WQzcZyuICrjtIbFLS1qIYE9Gh2Z13D
rO+WyVPaT8XKzC48/IsPtyTT2BxmrshXBTS7KTSUw3KHjEkTIspB9lyCohwAcsinsb+nNIIbvo2+
7Zl2nswoZkj7tgmmeYtqBmH47PKbTyRQjGQYRe8RRiqHjsnAsMvEGnFmpAmva28lwPml20D2cE9q
aZhDJMJJlWVbhwk84JAFAy7yZHKXw/LkPmuKFLmJ82XwfDeXSC4fhyj1O5zi/N/wg0QHcbt3YD3f
RnAJkYkORq5jQqSfVOqSsQ3B4VNDE8iG1iZl9CHkS6c3/ROb8wdc1jAScHv5V+xRgaUXnsSwNRz0
jftNdPYPZO35EJUOQGyP01eIfcgfSHxWbrPY7m7wiQdoiZ3QkVIDJY1y5VM3GUHUT6ER22aB1Nt+
D/9jDhlBIAghoebJ0e0EpDh8eWh0OP6L30l/bp3kAnnBMmfpk/fWewf7x7DG4xwBj6LTUS0BVpCh
cTJs8o0Tf948BDDdB3PC+BSJ/f9LyyRBxHSWq3CFGllaY1fBQZGBY8mcHE2yg2JI/kUM1ez/o0j+
ETk7fhiKDyLjsGQ46r5sBneD/uGrO0MSw/Cd+OhyEZtoDsHbf5R76uxKbJaNNfmSzkSOFVBZvUGD
69OzUofdcIbyHz2YL9Y97KWAySydwO1oEvwOazae/9yzNFhsvzf18/Z5L2EnW5z+WYD4DauKjSpx
htHfkQmq2aEjy5peNd3yvkbZ7MQRN2eJnlBwviYNkPyMYTRNUhMM7OHHxtI2OD/GVJdXCJYj76rP
/+/Kj22cMfVAzQFpAorimV+K/zUa43139+C/SQU9NvYWh7LeKqGgjX6Jv6WSz4pdp+t1fmrsON8J
PW5OgR0PN53R3vOYUi64efHbstRdafHKl1BxU1W13ef5SuyvatRm+rv4Tqxh9BcwaiCFkBeRVucg
AQkTDOgHA6QBVCEZyjDTD+DUPAXmyQQSQsMTvLxtURnng1zi8UfBJQPdQpnq7D/fZ/+ileMUbMyA
b2hERzy268Gta8b+VKFKzhvNrdavFNrdoBVWaEUR9rmXeNt1jqFvGrX9Y7v/Yk2VWbO1P++GHskb
8qs6o0sU+IU/P2skwWHTZIJulXrveY2dyUvAYiGeWNCg9sf0TmMVpV87gnjKiXAFiyj9P2ro9BDY
T7PAeP6RelgVg75NhyqnNl+5J+EWxcVg/Gt5uy0E22RTnn3SHhts8MhhlSDjXNJqWURIWrXahZgm
XoQXmzlru8zLg50jlCkxxSg0ZRCVq+kbEte0tdOJEoSDDuae9GS0TM0tiXhLfkwBlZfs29ROnt+S
CWY6AYrRajglHFYUTvjYcoeRPi72oJlSaumLYG6C3f7dkOZQh5DVo/LiW/dR2fLLHcjR+UukMwAK
CExgs1O43rwpRn/DuIwgNSHcrkltmcDmCbKrylCB5VOTLegdCZaiYz7HTz4koC3iWPxxRyZAkSwz
dyVWQ+1dc1KWm6D1M1g1TPA9qBMCfYnqt75iW/ZZAJjDCnxdzb54Q+8eypSgOo1wI2FSf34zwCXZ
+LKIG1609a+fWpgmEk9/EO7eo0bgV3dEVsHdEqhxo9x5P84NWCp4FleNczPjtndTsgHlOBVFulSC
7o5yTnkBrOUWePlJ/XlEmrsDPtCa0IDbKNhG/Hl/6nxdq7i3yWarp2FivUx+J8qUOpcAVvDcpiWs
HOSNdvD+mYpdBSHZW3RxMcBbAzQWyFOuVlGxKp+5/0trm2L/6tM+oo7KJptHE12SkiQt1BF1UJ8C
qdp2xBI0WZFu81HYt0p1wfSa6d8q4K7HCKrlh8DnUIuMrOznsNAlS+e9jCPD86Tj0gYreMrNMcAU
qvqpw/dGHdaS0NsYPAYrUCgzkRAoF1pUIJcrglZO6tuLrI+6PCscFuTG1rqdYnZhfgoHo6owrpTl
WRdOQNdlo3xNbsZC92qZDK320DataauW4IOHpFfjEUKU1nRgel14TCzhj0nkSgGwBM8EjYaO+h+Z
Zep+KSHY6ss9HN1QVnHyUcknJUvanI6coEKbsRuij18tg6VvdSFT2fCLAWorL8c2d+TrJvRX5lpK
fr2nggS0jYX9y2+I71bvfQ+1XgIxih6PD42xsTeuookJSXphOwIVdw4tnDf2cwKbQexr5HocHqiK
/kHxUmzqQMNvb44iLlIAwVlXFJ1DBvQg3x1NGVS9n5GJFe6O01Ksq4z6QF9tpQvxPgL+kk5m/jfI
w2zrB//rSwPVQutBMKKMsE5C+M/+G+XMxFBevuY2nGO1qxY0pEmLL1noHPOH8jDdz+iLhKKIapua
dfEerlYq4lZRWIfAzIcM99VIxIm6Oq062GiAEHB2JvvIyjlwTs7h1iXCnyyW/kUvGgSBGjubP9VT
UQJ8yEPcgQmkl/dP9WGb7vz0na0sNVHD6/KfMb3tbZgFJMa2CvFWmSp/vuSKiP0sdCvsEBrZzYXZ
qr/Zi1LLsMyDvfV/wX2gE+AxFIrcjFn5bp941zlxbwTQU4HjqZ57AgpykZ+3pWSLPBfLwdnLf2TY
2w+gAdhIQsiMp2UDnS/w5bU4ZNFsVhrTrOhrievQy9G2FvmCFwb1WH7B/YKiFfb/5w45/M+DWXNz
+DftitKWCwefxlCbfxNTvoHsBikkWW4nRWYLcxYSIgnLQg14JbfIdOewJrjpbOtapuuc1P7FXmdM
mhb4N9PwHXMILhS58HjVqDuMZ+9SwoA0NZpUI42+9mHqin5QCvCz6yTU9oxsaU41JYMiClqZZ0Nm
kzVq/bbX+pi8F8M0iUBUnxA0LNObn+/yb2RHeyeU7q8HbDB6yH7h91QtFrbhe0cwklCSfX6umBUG
TTzCibXDk1pNv1640hliyJM9T3F/J4zViDQ1oiBoe1LR968lJnZsqZ2lgUyWhCwU5N04wP99vhrO
AzXOUBvn4hT9vZpKwjb2Wm7F8t9mnB8fG/pUUeWoIydjV+m7HgpdWXOgAVgpKleum2z+jCwXdY7x
khfkXYJR4LtfMcEp8zSSWEwKydpCOjewqkAbTh5DqJ/GN30Tb7UxRMthv3x6sPFMWRdFFSzEt/iP
P0vk1yiZqI0Bm+Pw2676hYaKGlWGIy1gcbWLbRJxPW0ZcJjh94SUzvhFI6iipxAZf5mrWcuOLFE8
Lqc+bF7gV+Rzr/SP8+EZAvtrbAINUH7ZOjr++WqBD1K1trJTn/JQknRin2wD4EOp17WM2fVH/6ZN
Xxu7nXgwaq3OOJqwxU0UeOxRYXYikFRH4tt/4Qd8YK/wdIAPDDLeijV7i8FVbK2Dc5Qc9I0fTaR9
FwsfkAIMrxRYsjHAueoKZhA1eEoJmJ7rOtusEFH5Mj4Vgae2beMrOeqiHtxVe3xI6ZyldetAQbd2
1vGSbgriwNtg+1fyN1kOjILHMk13bChm41l3MJtSl3g6KdJKnA6dlO8Edz0ulr2GzLiJznrB7yN9
juo+6Uxe4w/AZPYr84m31OC+aGNbqtQL6rHSQB2GssN1emOBCP1/4+WmwbIGLSYUUEQAOTMGZBhr
sGR5pZ4O7xq/uaKT1w8t3Q3ob3TQ0hFNRSkehujObXlrQ++j7zTTE50t2x7sjKHQkoYsoU5rvmSq
G6MQLQL782/BS5HKQn3eAS1PansnRBXLmTkj9s0Wr9w/cwkWqXIl17FVPSJcey3nTe7h8R8sutRy
qSCEvWdD57TuoNEs6y5NfegLCiySl75/TL9cu4oALIzmYDQP591LDyh2rsVqBACrTq8jJX6CcRjy
O2AOP38vrZKgP9Pl8shdKEKeoVjx5dzip2G8h4BzGTeP6Yq9mgDDNqeFoZQs3jIXMvvrEvBNHr+P
cir4GBVKGshUJazeEgG8XxgAbLPJrqZh5/uhzOiJEs5s4sodIkRFdbfgnMow1HiVPHXMqWZ3rkn/
fSTsw6xb9ieDPKmTFMZT6nK0g9uUgyCCFo7WnYRPrAiGDCUmDA/eNHd4eXzifHUkT6iUWS8EsHt7
JwO5vmBjFS980jN5iVgrPHEHssdVowmQm14iLF3dRTzcf00W7uTkgWFGiFY2uySYGFbUcOof7XrI
lPRbW5jgVIAgiE+yNaLuxuB0N9lU6xkyargeeDkMDKPfi3bAYUs/SSwZ8RzckSJ3kBGnBeXJ9NT3
OsiwVqqwvHPke9CfZH/VJW0o/Lmsh+A+C5mzK/cl+Q7xIlVqmi3jr4B4a1P7Dss0BqR7am3L1jlM
ce/Q0YRJ0ad64okXKMtkrz+NxmZQ5laww1UFo7YatJlqqowW8ZQV9GtvFSOHQ+HBmsXue9XoIHC2
Jldoh71Kqp+8LOXva4XCeoVynczwFeLTwZVkd2gEaPm2uJwmK9pO+px2gKMcmDWQ3NN85a9iNdOh
Qdju2Pe9BRulwO3r6pexIybC/2RSy7PU62+6N+Vxu6kLEuvOrMWxjGBerwlnfTu2elUPE16lcG4z
xkN85caW5xETJCjA8KYSOYKPcv+Yg16ga/KyDePMYZEQ70O2K+lhypuprmqI4Hxk6buepZo4dnX5
pjUxxcuKzfqRwu1RTKrp7lZWdsTSAqaAdtIpkoTK/3pKDhqG+wnIKgLTOMmgRWUsNfIzz9NBfNDE
+P+LW3GBvZIBP1Q0VbQ5+beO9OTIgZDZyY9GM7W8uaZpSvjXGsogZDpGPmu/WCT7JZo0XQTFRZgO
gxTF6OAk6NgESU9wsMuamJFOFoR3Wh1s9N2rOhKCl4A7+hOfGoCIqRowlj3hVdLJk7gtvSAwQ4EX
TPSna3HBdrj9QrOBrSN3dOUjWUzH3Cc2FgREPlsseXddrw6rUuMU3txODU5XuBeygAXYbi6B7eqZ
2oj6w7sdqhmTrOzJhsgAj+u4l7qruxV9B6gbyD+QuVrvKjU0rrxAR3LJ3vgycXN1d0ln4TuZTRAd
Yd1Yf0kRRoHWT3qQyaLuVwFO6Bepqi8oUheZWixXtSbMy164LsmyKLxcvg53MyP/I/0+1Is9gsG2
fhdmAFrvq1Y0+x9vV7t/QmKZdhRIyDtmSz5RjHP53OohT5b/0X/FiCFwj4QPqAt7hr+SkAZ23/hP
brVw5ebP89IvDldaWKWeRSVBLgWeQC7SeBfBgUfg+sKAaFInMJ5qz5xv157ootfBvsPkDEyAxntA
jtp59UGnkaS4YVmDzjAc7/nbSaF1mhQKIhimjRnWnxE/DUUZwck+nZfpnCxEE55PNYTLkAvVPLVB
BbYW0bIk04P/NCgi+ezFJE4go6vt3xB3aHPlyv41ISzDgstI7U2Pa2DQgSxAY5SEwmz2s7db9GTr
/JcyY2PA2pmfJSsmMc7jnYREDuUv/ZeCzFFWWwmU1PzxTATbM+SCWtSIjLiJ8aqjm/tld1MDL/k6
LtertaRT4jzI+XSkA/5IwkksqCwCJ4OrYpukbet9RwxZPbxWVioG0SpubudoyOqZUBIpVYIc8Q7Y
et6GxmTn5P1KVKqNB+Hoj1lWB4hWumW5bfnY/mktOu1X/TU/zxtetoYEdH2BjIoJrJUOGWyQ6xIW
ZMh1mq1heBUtbTw3dZtmbY1nBq5PKSMmxDdlbzw/TB6nJ6eny4mWlLaZ0LtkGfcvScjM+We9ecuX
62dWQl1jE0mQttGajnM0QkaCu7pZc8p1nt3eyFDtpBqTvGI3BzSHE6wUMVFW2cO1/849Ym0lAWSN
nPzs8FSLxo9wm6PPD3h/fytxf63smEzfn0YAdsclJUekjzV0MMohXgmS4othcHHG3s6OfKoToi7y
kLImgUXvc+Jiq8XrrmsPcI8XaZ22vU8ex/ADoDnWmlnlhwApon6wSLRQ2fZCKeab7EZFmIzrfe5o
nlDVlWPGdh0c8fLd1tLAydw95ZNBEMkRtgkPRnszr4mSyJXKXpDs696fp/E3Wlu79TAYKMVmHU81
l1ebD9v9jZnRNmh/PfrCRXR7EF8OVMD/X128ZOVhdPk1sojwYmY44PkDVu7SgKeCQyyN3sXY1qg7
/6UTgIXHuqCSQJ+es/LgmZ7JOh6i1BY73dSInOdOzMlwasZUSttvj7d/2WIVJDxp+ORI1PjchYfw
f7kKrm8Ais/61hcIwqyvBAk606NEGxWwovvi8PQuABOcKxaU4I29EiRYOwrwq0Voz/Is4eureG+Q
kqlw1UGFYTDfQpJcHyICcrfAsHNlNH1E+5jBxlRWNFxKu+7bQgNy6Pj/8kukZYnMaoM040tRD6G+
G8+Q/mQpqYpIfJge+7e+MHwfakwHJpySxzS9+HULDDv/EYLC0/oyTiBABskJSRtmK8nUSlLez+e3
44CzGY6XqwuL17Qxd4FnYz5hpebNBlipClI+mUiXu0si2F5Osk5YNdaxSYe9yMR8wVPdmvAOzsBn
kyOV08d+2+wTw5wMdKltUQDkgYlGVYSMfLIqQoE5Tf5TuO1cfnlirGgaSDloQxqP2i35eez0v/6O
iT3XcwhJbf1geaLQN0deP4/Utu+2/SnLQW4u/5Q2Z709O6jSt45jtCg49LLEbFm0ILRn9T/hPz4c
61QD8fX5pEWijEnBAjXYVyOBtw6HmndBoQmW0ColcCmZV3Mhc/Od07hKcIhT84qk73QO5Y7P1C/W
p6CNyUG6Gk3PvWiEfCW0C5qFDOhSu5joYBfXriL5gA7SpOoW+LXxB3WsX74BEPtnCWOz7HNgW6tB
Gby8Vu0XQnJIRUdNmnZdlHD/k1m/34ccwtZkIqIt6+mrsWUgMFHQ3BjpChyVW6g6FiVKXOiyvqwh
pwKvzIioWUuens4Hip7m1+WlCILbOQFqRc/9K4qdu6dlCLid8EahmqvCdUFpV9gIoAoOPdZbh3VU
7T6ClG4yfvjHEuxXRAjKopAyJ9MFuEKGcNH7dvkxHagw1NF7nPQOW6wVxsmukYDM9R+GlkzO1QZi
DL2vMqswDz7OujUrHNHT+CAJM2MPpsI9rR/IYaC3Bueu1ZP631oE07XSSbl8g78truBZqHfukPAI
RZX/kCSfyDOEmMNXA+ZqfynSwf0Nj2c1hnU9YwkxOnegUFN8wRNujOg00ZetDoYPP0313v+EEvep
NajRY/D+XLcNzTmessBeQW2xgn8LjAIYwY2O9aaRhr5214fZ+67x/1i7a42VRMNF8V9ZcAxK9J9K
DlnV/3zsGP485SMuXnhDat/FiUgD1J4oGzt3SqWLGi4GF967RmagsM4ePhKRdY58PK79mbHEGK75
3rBVvHAfMnVY0RmxJfmspYWBmyKxdl/zTWBXCrQOJOb92P/Qk4maneKV2BriLIKsz08mxbJwiIKQ
N10vgkPizBCaB4OuIq8J7kw/PyRRvj2B+IoJ7gpgfzMb4T3ygbcpmzZX5rvHvoivOs62IyCJNiUD
SQ6ouj0C2P5cy7KqL5JqlnVMWDCL1264VyMxXDcJJWcQJ4Mmp+sdvKrygSKGiSZ2DYUnFeW9tlUw
U6K6IXqabNEX2AOWWUufa2sugBiqclpCN9DRA2A7ih+095dQHLFrHmbYSOSura98zNF5hiVCWqm+
TbgxruEBEINpXHDPo45mJYOyb7zX3nZMwgnHiGcxp3kDc9oBG7AKkLz3RNnLQDwP02hMw7R+xfik
bwNn9G8f1x0MnivBdGJL+5FfwlWMFSQPm24dHW5meO7a/2hn0+GbAp81vm3KfknSu08/OYb6AYMJ
cTthDMm6qSOru54bLMATJhW24N0S7glpEgnJXCHPl/5RT0eAVuAPNFpvMp3cTsS0vintJnwg7z1K
euR5jeWqviYesk53uzOQcmpKz4EwWygzGAM0jduwCh7JexL0pQT+L/wdSfj3jYcHau30tD+zrvjy
UxzIJVvYaD7L5XhfZLLFs1Y8l1ybIJMmksaM/GYwJIoKFlMw9w1TBVk7i+l3Gk7Py4OtAsgKa14I
zH65lzhxpgQLvrjt8hOkBluEDQlDiCZwBp4M2EDKMyt4vEY9KPOS+bZnJ7bkOKGU5fTz0Bxf+V+z
u51KyL30Pvkpue0SkAL7Tqr+E2PnXSgRB7HUTC4rCOogSvCGfLR2SC+fspTe1Q8Ab8jyLeKZWih1
1vkQxc4w0uaaRKHlXYBv240InzcTPeMZLPLLzI3i+h7yKb1rbX0YJoxnuSomiMW6A1mtIaRINjZP
QWCrOJYbPJL8SrwnJaKDX+tHXyYFr2Be99bIuRMH30q5S2SLb6Jx4ZJWVadAsDf5DOIBI4Tw8hgm
d0AQHFp7H8YB9Ke51OwEwCKoisimEWz1QbUuhATfjoxRV0N4188T0opzn9Q1Okir0vL8OSdcO7xY
6aK1uW2jVLF8sjUy2ZXMkieY/GED3ZTR9l4T1aaibgZ9vUv9Cdg7N5kvAhOF0BRZj/fHg2LkuZ7w
Is8lfnTN2qn2Ng4miR3O2A4zYLVMQx+Ticdk706ql1DjYnaLlkFfRiNINv0k5giTUmbBa7cfjqXj
zn1AF/4cU2tE5tWLW56up1pgwsLJgK2YtDf5P6RfiujZILtgyXGTVDa0P3KO6pHwsUf1pBGbdYs+
B+YnyCYrfLeQT7A3iNhfV1HPXJiQq+3Rl7w4RhOoQ2t8wVXzBbgedxPVV+hxALHz6bEbj1Xjdrel
myh+nWyEZDdQiWEqBuqm4/7bBos7irokkGixYTD1RLzGjIE+dwXJB5jSQR61gD8RN1wW9u3ElKf1
DQmroUM0jgVV7pOd1Vctb8bKYbsl2uH2eZ7bBzU2YiUW/0qjH+gYPXY8tQMlSUhq9zNUc37tjqo0
UGAJQMT1y5QVlvtDxCC8Mnglh2CzIQwCvvbu8ba6nPF5jTcwuXngBaZILLUohZLJzGFKUG2KfuWs
DdvzEGt520hmSPDz+2QUyFJgas9yGaKsIbuDCqh1gsNwL8TojG/uJabN+eNWbZJgA7Mmq4YjNipG
VdHsbpkUfjm3GX17/UGXjJ3pRzfboyIjZraLGzlVKU8kRmWl3ksr1AhjRvGFfAufn3bfSzn26gvv
DV8/cf1vvHbQlM3PFU9Ox1dhs2sKVoW6+CZbOnzcCw7RLuOYZJe13tWa0Ia2ElAGxdoTmrbVcZ6+
7CPckOfNlfqgUnqa5IgKjn4OZpdVGcvNulfekj0IIwLsp5tM0gJy2/g1ZMTownFsH9JMO9KNbp/2
ou2zp4lik57INSBD7Eq2bn6Avp+PM4TvPcw5Yml3jppXSkwNdVBLtpsk28Q/0eA1tvW6D5Mc55MV
b3bzS50ERglhjdYSU9Bqlv6K2JeNCdg8NXXQ1MsDXSRu5ByRXvsygPnlZO57KWQw29ejj9W0yBms
7ecE1Wd53NrPEDZ0e7uaEQRjzUh+zI7TuGJEYp2tOXhsZc9cYcqZt7fFUhxcxVU7aIiQxBIPd+6G
oT/nDmEg3juBL3bg1BZcpQ+RaVRmI1AxKg8ButKsgMYVVTzqtIescYo+1jf4h5TVtuEOWRgcODqr
9ouXcX8WDEuVwlfmWBW/Y3VT1XVoRH1YHdkLjWpWwslY7PMOl85adAUWMnIHIRz+YNEddEDvL0Uu
Fd7An5JUjkCoh/AB9az6XMjl814M+nkCZ+Pm073R9mKgFxcSjROf59OtU753VDf0rRYiwMtS4IL0
OA0DXe/c7jZKeFl7THRhP1hW0aWZ/0BVvTqazdOsozzflG+pIapeOZNl38Mm2LnSRuKadItC5o/P
jb6TQuQRpQQA3Z+Fv8rNlMRv+ubdhcru/FTk56fpO9gv2uk9znXYw1HN8etOZhoQXyWro2hOZPAp
QP8lZHCzu9dOISNskYHql7NSqaTPvY/JH6ic2nX9PkHy0wos9kjAEnQph3yNGVhGCKhxwPXRxc/a
uZ31JsShGV6I5g3fLg5OZZIexRAE36CU9vCtGgvkq8ib7YoxGH+rgFxnMP6LKDvPPd9ohu5KUHok
49mZkpPDw/3o9+g+C2S10Ob9BhXq/rWtRseQ8qKo52S11gGIVR31uU8cjIW/J48E6sZahHTkIC1+
DbT7Bf/xy8cBhPaKgJRmsqhFdUlQNwQ3rjtUv+jQqiGlvrAdb4Oh+qAGENqiIgwfiZxHg1GgkjIz
EhxwjXHh1ac7RuQ6vQhJ9L0wZKm2ecVBYQ8E2u+rq/S2wCtx/SO+i817DJlsT+5gtiLwS/lyEsLb
z5tPG0Cfg1b0z7Dc6jQlNNobb6ALCJrB5ziZ5BfALaAJoZ7Veu6ex5atmX71VJAcZY+RrnxBguvs
Ha5vYpXPT6G5y5iZG4AuIwR1iLSS8vhGIAU1P89pE74pZIs1UuAPYsXZvdxPvwhABE4659qpIalB
1UhpO6HPE6gLCgh0cEvvt1N8D19oA7GgS5gDqISi94tQnn+LWcJapbjm0C8nF4SP+zjh0n5yHT6J
1iW4rtaExzpgNur5LuFMJzVW2oMxZURaUPK/foA88dR1fvGFhmB1DBRLTAIfPDsYXgHmGxNlvU0f
XRO0dxFTcjrIq8RuQr3ia0gXHvSvB8an+oGUhSuA0lNaFASpMKmUWVvcaBMRMNBeJ4PUAUKvrC/x
IhmflGjGM/BnD06wCfLKfahf8sagSMioZWoow98zsbzKCN+LomH6UBkMITkj8jJV0fonTqZKSgXb
MDMjUbCsCB+Egts4rfbPUbM91pr3fj1k/xfoGWQANJWF/DjwppPuOa0yXfVr18JanHqJKe5BDVar
Iwb59JA71j/yGzRF7VULBZGEM8MRtaNNahaRymtrTOl3J5QZr6MpW1mIRpE8cXPcTEnixK/f8bXN
+6dW0NDLEBtKGjEXgzs9oq0mRwXZJFYyvWeKsUT48TT9ZJtDpvY02NXa7KO4oLrpykhb7kXhv9wd
ZIP1HPy1mOrfdKNb4ATrNOaVSKpPht3cRFTlfeUSH3033BmCHndBfB+dnuWvlCiIXjvkYkR+lJag
3fd1pFTacuZPtuUeolaSDku3EESG7xsbuc0Vu7d05a5BOfl2vO2klT2d7Mvdc+UOTjZNFZdEGLdH
E7H/oqZPfin2FMmvvY6iibxImVYrRH3d2eEWHnrZdKXx2CyOIwMWJQFB7cLE9SB3EhlHr6oMzi8n
GLkuC2YTJhdQ1Z2BTc7mmhYN0b4V5ed0m4glhi5W9ydSjUGfQOcdLl7+Gt26ePlYgRNl/3Xyk/SE
g4eM+EWNrtzcLcl/dTiyfHrAh9EYwLnAIK/HKOKgT2AddrSgmPexAHzMtr8k+vBgPA4IBdQ5CMkg
CtaHa/3yau8qROOGpD+dyBLDeLhlrW3iBVoq0wRvWj1CMeAsITP7h0mUpfeKGTjUZU/B/YtKo8/V
nCpcVdFfWfQbSw4bFV9oHbDk03rDCeKlH4HBmsDTuaBlZkmGsGO2ctxcLMNRvfqJ6l+RKJuImIzY
gjNcF0aEnUT5o0nKB2dskas7qtFPfTrL0Fr3iy0xXpNovp4F2JuZEO9qacSneWDXglyPgmlAyMBB
PBemYcxZg0cKRoWHOIafn5EtT3tT153yQUZzEZUN361Yy+GGoNg8o7jRroC85nTE5cF2enroJIfl
0CTyuKBWJBsS5BJrfGgmP/gIpBl2TIFWZIFPz064be5Tyg/20wi/kVg9X3pUNKXleYaOG9frct5v
8vjUok/U1Nq7oqNnbwN3fQsKbG6Ujh8Rkloy8N50Kw48Pe7x6tkyAA6o/hvZvB9h4ICt8gLCkODn
l/0bYcw3VrDPs4G3vQ1sQCjJK9AdymBtaVwtgp1y3BDqno8dqC4o7xfYHtJD1MJQDT/GBPA1pyVa
hLnBXjFw/iD+2pw9wgbQu4GTSOovvvyOJckx62IxF6JT7pOzuN+hvcGfXQfLiNby1iR+DNE7Ge49
DpODW/4HEY8VgwMkGZ9LYEfZc9ZF1QlV22/gYBer0Jzkui4naptiQtsxKFlg4d68ZmjuzFzK6ROR
Lj5Bp6+Z/SvZA4caRHf2ATFIloSWADA2EIh7Tx7BGET3/Gr8iqeoH3ONGeW3iTvW/Zl1eWnq1IZ8
3DlEzt1k+ViqEHQX3iXsiN0ucFJJj+4pMtgsvf7Q9ZkQ9ORKW+uqvzhTPWx75Ibsy4+TZ8wQ4oOE
NPmCLVzYg2PeT5y/vwfv2zR5U4DshRTRmNAyH5HnWO9TJi6ru6FAfUEdXc9zugHJvybqIx7J2DrX
lwiCPx+A+0htB51eF0M/2qg+GOOTovHxQEJmj/tRRs6zpqEy/uMdqtIHe2VDFkl3GAwVDrGlTVIP
6IAi1LyCURxeblYJAkgiXBYJvfnVn08/pq2WAxU7E1l72zCloQMJDq7fc/k2YY6jOzIj08LL8Vmz
YppgHn/k2fexyCap8h2Zqe8GnllFYQnOV2xGWR12pIfbHAsx6+nt0NdS8mEDcglDiz+ltlKwS281
L1chUcJpb9UAdvDa8jG49YiLWRLVPhfTP2/Z9Umc2C249X9hAW04J9iTLKp+zHjzy8PIwBCCrDDB
UAG51zuwSUrbf+RmQZAd5dmKvQ/tEo1dWU4m6mNJiqheLLFM/PZgohqeDGvznm+razzjyE65CEM9
tAQSdjLurhmyRi116sq3DhNryN2WJgeqmAhC11OYWK4PRWa8Q4dNi0FOGsGodbRPXMx0ktf/o4Ua
xF7Y3j7i52qcLqfxwwnIeI+t6TUu8DPwOj1gGqhjcXspoOTVj4eVkt1+GLdt/TDXz+Bb2NUaAh2G
LqUlXDcYXVfgQxskOFClS+00f4pViK5OxIYLm0eKXvQd24XZCY72h/pMBrPM50qntaX5qB2hoo1j
xqdbD1COVSDbhD1qHPXGpREV1RpbtPg2BT3vRHiW9D7yiQbPuOTkTqRCaDu204KFIeWknRI/wv8q
sDe83WAt/bPtshQwbP8arxmU4BJQCdLbGQ7y3nRZcO5ABQ58gVSm8J6pBIjV4fdGlOBkqpt7gZ/5
/enFoM7Y9j3Xux+KlM6BxrhLeECUe2wkTbdnYuon5upHJK5oIxW3tqoG2ysNF7Ph5tLKa8BPSs2+
VMAFszZ1RXetA2HgKw8c/II=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:25 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GRe0CflcFbl/KAtA6LydoBbFCjuB0dZKREjfTzj7ORVK2HgiN8yCNILOX+PmLYKz
aBsb5yxTxyjv1h255IFMg/VyPbiXc9qcwxYrTJ7fmrYE7coZEIGX+Dif1lrMgMxY
JPXFUzNkSkOXX2aoQBtaWwsmpd4gfEHMY5BqmsHyCPY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12704)
t6kJS1rQs7ShjOm5MqlQsCrZRTMkIgxy+4sIJ/lzgrOqj7Vl+gyOl741oF4Os+cY
KG5sh9iHZhULWQw6qZl21DnqwnP5eHt68MPXdbazvmFdadzuOfJ8U5DeEqZg12aT
wtjO+YOzWwZt0FVogdXB/PmL1JTlEqWbuAjadwII3HMwqgVql00AE/lXsoL0iipn
f5hVlimKFTy+JehRHR334kzge6eZOj+yxeus1uLfgYBjbzkcxa2Wn24wEvtx9xFC
yesNs89jkjoZUYE7NwG0G+w2Paj0afSAsuiJUUBl64/bYIMlzmsMeTrCjCguHffE
mMc10pTRDeSXfjPTNyPUaHHdjCCEBCUfZoAWnj4s5pQ0TPMSlAAyzspmBlwdJSK5
8TyMTeefoQNmbCLkJr2htScUl7bxujlaYSONaIYYUdBq7Chnxt5g+lSiOMOR+uwM
4tM9H3kokjEDOxKvnwZh9gmIV2hBQEPTS+9d+Oa53M0DoMOjptD7T7pt977dUpo0
91xfI/jOMaks9ul2RKnw9taAQq8Loe94ZmePpS5Nk9pMaHbWN2+aSxARJdVjE0ZX
fVONFGtOjvItmcgFXOp2qRApun8yH5olGKWlbhaCsJIK9zl/qx5KYqTcnk19FOmn
yFh8hUFPl2di6lTAVcXqqtQSjLrB9jGSQHlHrd7YwDmtQe9ySTx6fx/rbE5qB6e/
XcwsuEfxdtnogM8oRc4NFfAMiH5Q2xcHFwt7swf9tMB+1fBtN8IIsDtxzXqH/dcB
QpVVpV2DO6bGt14sduIYW3jvCr3dpyVfnqx//uPsIokMU52TCIyAJh1EKyebLIv8
z2+ubmoFyyMTUgydImQHXPS9p+lgdPi94LRIcy01idNDM87P1zbUo3deOW++vkmL
Cg3DiPpfBuC+lxQqkGzo/ofA0Uw/Y+tOLBqtzqXvzuUKxXdh0eFxptcmYhT438fM
Lm5KI0lYVt5jTQ750kBOqyIx914h4QikMGJl22Fm+y6Nhw3sMJEwH2/h8MiYLMDs
SiupOC3dQrNeUxJyh00KQWZ+SK3oPqwQgkDBVtJvX48gT7bmPLBgTPdL+k5tlea1
0seHLqJ3aIRmQG/8Nk4I9MtZ5ZqC1ZzzpgJVG1JhSsEYpi0C4JVmktoZAIMSswBV
BTOWu1Bh6OQLnwYzOaMx2DXMwNtcLtlTxa6U/HfwK/sz25w+XmA9EdimxMlyaop/
/cFH5eP/egSc4vglZKok59V6vaQVIAIZhgch8bB2MWMjh70lvXC7eAKDsaNt2dIJ
Y6XAr5B5LVzwoIZQFgaIz5aQwdOAyN5M02QZDjFOtzaIQZEYdoySx+KIckOm9BgA
tG2RLrnZqkDBJ+PuO2xdOqQs+3IM52uwp5nIJIKj0rzwlLv09z05RwVyifmC46EI
mYXHzA8TRBFTUu6tYK02TybgVMq6hNkBtA3Un2qVpG5rt8CXcrIySCZfdEZ4yPki
jKmwL9/WcrnzAR6yr8351kjvAPIYP7rm4EtqUBf8u+PrTUP7vQ/vUlfVZ3BVTcPb
P/yFdR9FNToYlE2RWjM3IrcdxtF0sk/DL/mQ1Qc80FWyBe5D8E1cJNgCyhJIQ/o7
bCrzSUtp8ojjwgr+KysVBpM/eD4ALDZ5KBhZINNpTrHgBNHTMBpTtY8tj0RPtDiG
8wHM+R+CF++cKBOQdB6R9TMwbnzDhatOw99OOsMjILTVz9IDeZkiB2ueUiG1Ng63
UUPepZ/ks+GUO8sNvfKl6T6M/8CRp8PEBKg3my+hBPG9Ic4GLX2DOUvQuMMNEDSA
oX2GUEBcHE+esZcSLllobyTyUpYXqh3o9/VZW4JxXipJOqW2b0XratvAMx+7Bzjm
pJKze4FEpAutVB/wEQfOiwPWa59c9xnT8DGtkPaVlFlJlg4zwFmpnTzNBKsYEgZe
EGRxcESeANQeevAbwZoPWcvqIqcF2gHBGTcrvjX0sSqVhO62IbH/KONxCiJifRsA
/Osn9n8HeRs5dtW6X2Bavpail8HzuX9KZYmLGs3lQF4/uxHa2aaVyePmYoBcA+R0
F8GtGVQS1vJ6foFbOgdkqCUpN+IDgf9l6a/x51kETAIGlvO++0QDDs81k5tkxb41
1uogREeyOup8gSaUBHCTio4hjOOuWacgF2tbJnVOGW6ZeJmaXGCx094aCYV0dEDy
1yqnMRQzC/Obd6n98rAVRqIaslZNGuiU/elu9aylAE1Dv504IBNRo7IZbPrkghyq
abQn6FFsn1CNn/bScgQm5glK0CAGVw5NvnLrVTuqE2Z5qOB96vMCTowEQSQeVgZH
lekLFfhKeQy26NHwBHkE8+aSKjEscl3/NP3rnrgQSirzfPOPD/vp+2mzlJDsDvcB
I5olWFAGfq/5r46FlBXUiQyja9DlXAuHugGcnRslyfp8lA/4BC0BaVmv8jVTPF/v
dJNJo3sR/nh8hGIt4xyVSnoa+5q0PXlS7MjKKDblCSvgqNZ3gStLKKRzxBWLQN+w
FKOcnEttCpjpezeJ0OcoysAVZNJfppCfdJD/q777cbVjv8lLSrwgz205EB9U6nm3
3ai6ricMVM9Sxp5/6exIdjdeayAzxvYpI04h6gHABWk+Dkq+WQTq/muDMlNPNhyv
RMfIo9BlM1Cm8AIctfsv/DLb+61vUsjneQBSLCDS9b9tEmOsCZhtZM2KVQhZ8Qm7
TLmyA9M45nqXHNN8rcX1jTLooianAwxYz4jRi5AWMdpuYp42RmlbIe6AwZiDDgWj
Dv5wVnxa1pqUPfAoGUa5UL7OVHExsUGCyVuc62i8plPvZVkUzCSdbe06x6FOiW8W
/vZzOdni3+cAaCljgEEpXx68SgzWO30TEnQ25bZehw5lZbv1zRIziGe2L3YhWV6d
gzjisZtRRyF2+juasomPOFlLa9TWSxo4VMkjPAmpJ1hKprPcnH6GsTWHroB1L0fF
Bf9rbwVXOIQtSNslaFXir+W7kw+plaigDJTIDOtgDqImEKhqK3LtruALJZI7iwaV
K94+5QoUSS8A/3Gf6fgNp65/Oj37R73BB1dDxQDwx8XvsoADZL/UQ/x62G1//YHb
4SBQgFra7V6mPIYyyxQUzs2FpCWkDl1Dnpy9lRIS4CDPOfFhV9WOdj8ilGtbuubH
hDwumLkjmjWQwRyxq5kQezbfLjX3o0losJRm5Dv0ljM81ewtjJEWZSTPuTMyG6DV
cyjOqtObIo+O79v1Yu4kIHOIQ1u239bfRxaYgZeSWBqpbmow/zY+XtlY6ttWG6dq
DCHfqEyU2Ndkn8nzyHcMu0ppl2X2NWhDXDB8fUpjQrZxygRyV6w2v5cLdrlIsIzL
8h5NIj41P8p5PXSbITIlisSJbc6v101o9MOsxHg2BwLXWxB00QFzAi0kWJ48axdK
LjdAdCN6Ce/L/GY6QtgLOIqqiCa6NizSCWOdWF2wVqJ2O8gkawGYPrtxjMKW603A
hb1qhzTRnX1qghvlf+Xra1Dsmp7fnpPdh95vlMZXGZ4N0zo65fDK1Ksucx5CJEwc
d/6fS1gXi/ZqEo0NilyO8r0QRkjiZLnqJrWoePB5SMxOQz98Bfai2ny+H4itRkwm
tuzyjVymQgKhiEIBictnSKcu95ngaJKB5o/tteVgdCoMURC4VC15K/VZfGutLsxZ
LRq7Y8rrPseajhjKJDhRzNE4vag0bUBDDtoBgaSh0GGA0g9MrgOOr+/YZ+62px48
3iJxB1mIZEj78tl3sGpM8CmhmjEcnnoGYluKegCdVwxjtlhIpNnRG3iB6FAoAeDq
O0NhW0vvITSIQLIQolsfkQNObaS7BeDWhQH+AmbScO5AYksN4aV6VA2R6IeBiOPZ
0as/LWBW6n1CIhVd3ebR3qk2KisogvUscm7AXmW1E2xBZz+oBV2LDUfIb5DMGA7/
uxs8CRDorp3tcABOW3ef1qrduLeVW4sklGrimdi2HnDc0iJ8wa0UGaA/H4UIX6Zg
7bFJOcWWECI81+QmVl0KT99nyDfTP9kAUYKmm6eYztsJKoP4Q4QnvytELaFVv8RE
RzBqlnwRnkLBqBaDpavnyH2bd9Kx0DMOklfxbxOwVVgWZ8oMBFmlGzmAeENf3Yup
Xgvn1ItW/DcrSJ6xwBz2LMdmwgPlIqbL3lertvG0nDZ/eJCX6HwN3gYG1LtpcMSX
LaDfXj2mkbFp+khOGx7gxAGq0w4jsbAJfw7VwARkuHbF7CggcwJqlUT0J21/bGEW
0mCedIsasNE7y18Mjqpm3weOFHG1BisacwBw6n5QFUlZersn/ARNBSpleuLXduCs
kpz8Pf4V4cxJN0wPrBEWsXke56e6z92E1laRvOQqS3i5rWTu7LKFPyWO/oC4OWfS
W5jjnJf5RZZqlFBTvUFU/39jIqEMFJpXdVuY/uoilmG/VVur64xkd1rSXNpAvMni
LP52KOEH6pR11sCXRWdsCVR4krnZrZgCQ5/fBPuaVQfMHiK3T6N7AkPH0e0dy2KA
oVwZGpIgGvwPbkxRYLW/X+VLMVKR1odlXwkoj4YCTvxq55b78zuokrWdWF+Q3TDZ
WqPeGqwem4LdaIze+ASwaMX16LmlS2D0+Env8Cr/A9pmUAz2gz8daUEJ8RxxKXAV
iIxsG5fOdEHRUNDVVw9VMk9xGA37r54DHpg8Kr9mbGFqM/U2+UeCgMblxXX5KYO8
4zArnWdOy/ORPRpyy/aJyWNRpIqKWf23PTwh0dHP+RbR28E2zR4aoiZmZDJ/O6KB
6zYKRQ9j6QLxCLlANC+ILKV/bJWCydTC0XY+2yAUkm2+6Qrzo9pGC5/a4U9z7/W9
18IGmVRUfLADgh6d6g3ZTWv1nSpqBc6IheCScJcqKKlBfymObtux1A3JFrhEQXu+
oHWJ0GS9OBP2F5GwsRzWhvRN4LBJFy1yVsyneF6xa22xUefkd0tibEE2zOd8tyNY
CWD0yKuqtA9KA9okQzrm7dnWfe7iFVmTOPf1AuN0c6/J3LWbkjn53xkG/JgZDM5d
D4bheRUm2ZYXUMOpGJ+NqYNqffUCSECPCLpcgvYOdcwra14sT9Fvilza8m9JxxQK
Lf54RLSK3MSNcTU1M0BOBLwmDinXgdIDyYPKteLtP1Ua9G9KdtS3oewv9FzQDeWR
0H738ZB69W5TANSKQWK24HTdqR8L2torkHrvWWJxLoJccWX5PodOuuYP0fi6SuAt
dKFVReZnivOEwEI7vcUczRj3voknSuV2FotK3znyzs3T6QM4uWca4uostxKrLKri
xtpwL5RXttYcMVl+9wpatBOKxDfr0nFfzM+Tw6/NjczK1Xk8Q/Az0YeFOdxksKPY
w0RwAPAMCZc/qUpJpZ/+eKYJsKOvhZuzGarRHNxhHVOnReL6od6AKkOSX+Bsm8pG
yB6IyzycY0V57LElVnuqoeAqjFuS00EsObVoFrSkXUf20u6MnV7a9yzM3U1h8+Il
b6c0q9HsY4WDoekoeK+YGYnnqDFOx7K2PxCi2cuMO04/nsFGqu3XcDv2AJEFMfvb
/KYHVkehuEVql+WuhUeV7kEAAmIxw/hGeAVcJ2QGvysQ0MWe+YWu5NaLb/HKjpN4
mrmCh0j5u8sZxiYCD/Sl0DYKe9cJ6sigvsAkprXF6BcGmoHfMETud68J1jZYNW90
s5T8Fz4uaOSJIT2trx8iJU+x2YiVw32QnyX0yOjrfLpFZaROJxfKUiwlYlqAl/w7
obSzmFr2IEThIbFfDICg7Mxpl2EXEjVD8aiwrc45bYuFNUkJDXuCn88IWsWrX3wK
gzbE7S3drWUZZhW2daP/WcvKQpUaRYSKyKZwy2aV6fLLkrMmkUwNLzOatfxuid7n
LIo414c5IpZEEAKZRRPhF6bYO8wdt4pfR4ZRFn+iobFTUq8XgtdCzfy8DniOd85t
2kzWIdv+HZAnNcarRlvba3qXanmUTPhYVZCgSRQCEFDn+0Wb1VUAv7jBF55NW6wR
vWA19lwb3uEG9jQvmh2CIhACvyzqp1ldyhlJYM6COJC5+Yiq46shlJM9KEaI9eUa
cRqjs7aMa/oVDmk8m7J6LPXeAwm5BmcKGQC1hsVMhVtR/3WycrGKtoxqldl19tgO
2Dgba1K56Sv50rTVjQQuLXzDrX8MG8/qPicC2GL+dSjSltoA9WbvwW0WwL4b6ahe
zA8h8gAiyBGPnZc2iAs+TFxz0IMuSXkfQgrgGXBotPoLJsgc2AGgvJcKbQ9vnhcT
v84+yygmabbkSRIBtgixMFtA1EPlwkARVq8Wntp8MU3Lx5x0A/sZPoBidbReCnDX
q0x+anqDwpvY1NRhpLkLax2Gbxfsh8gzIEL58uPwggZPG0kLV2WjQdf3Le/6zXDY
Cs5NBgkyv9zIcPU60fxxexWMytXm/pm/GyMLuPRZci8vp2YjYxEH1g0biEUN8Awy
BbhnUdAb9fMsLxugiUViva2N+fn6l6XOSKym9IvkRX0Bs3StCBA/FB10h+PsF8Np
YhKtl2S19iaHwc2UdVkn8myGvoGmUWGhls7PhBUGHqfr8UnIWrAhJw+v/9oC5X7p
XVVSH3Qc/DRpNyYIrjM5optCWL1nORFoBND/qGvIQGeX16SP2cafh+0eU6QxH95D
1qFYuyKLPrAsCWiivhz/JX8/NK04y2d6hlw7D4N6c77e63nsfAiXmDNB4YOxmlNg
cxt5vUQk0krVrookDBznzu/qeHYxIET8nrX3BxN8DUdKEKp/NWX4KIW6aZgBVIld
qaatdof+i7VovmOUZO7nMSzRfO0yvQL22OvWUuv0OZR6fvRKL8WJ0DJl8YLGFtVE
PGXPD/jtwSgkFzsn1c0+mfr28+6IHziY4aAtD71GUIyh8Ui4OQzKgCgcZii0dYVL
JboqOsItwjVX6X21TW3uUDxJciihLL6LS7wiKokCoXxWO4YdeA8tgjCIC+Jz67lc
Nt0LW3BymaVCSfjwNddVzd5jzsaX34Xe4XswQ2uk1slxU+TctliYPv1/pOlRLgNp
Pj1uw+2zLU5bdMqW9zU+k6AKX/GXu15xeykCz22L1NmYk1ZQxma1qBi4dc0pQPEj
EJRikgQrzP7wwUsAZGLmqx83mla5x6jB+/MkyuiWUfSDrCUG5q3KgFoZfcffog4X
dymDNyXUV6PAnnHWpLgPMIKIlSCC5PYJZs5WpcO8k/dawdohiQLo+HVxmAWlkoiy
qy25HAFMa2AAn91WtCjjcpG7AFZZqA6mBI96NE6QsoND893G9+4/TQfCQtPVUmOR
YEpn43L87T+ifVsLuJy5sZST5mo8Ugrc8A2RvewJfYo8fua0BcpDCaPzq6zFjUKw
GjMMtoYRHCzMDZNL8zWHAb6tEu4WH4s0LQ5uWpvqaMCDsCjoTWIlLf9ZNIH05z0x
lJkDCcjRWyf5m06ezLIjvDForDNSupADQXYpv4dMoEe/gKlnZ+49FdoKoYKJH+mA
Qf2m5JmLuwrNnuPR3dJR3Szedrwcxe+Ob6GLLc9PXEGYPoqZkVSxC7A1/SGYrJ19
v6CtEkWDetlTn3zyFUz/Slre+wgCFscbG6gjIUPXxg1tCXGpfdf10w71mVolwEN0
AMxuY3Mw7iDxUNIL6ZR2pNXottViGe7KQ9/B/4Noqrtpw6FkiuYmLPoQUiVd9CPB
1x0R5lh65UZhwNg1ur8IOaIYr8mCVSREzCwqg9Jtq9B4eR60qLUsxCNJ0Ol7tnYn
xn+rp8i703+PsDh9lcD5BjUzE6eBT9bSHaVzsM9HgS5xuHy0zXZpGBKIeGEAr8eP
EZcyLoQNUlNGRqGpZ+50txOl2KvM2OG+lr8G5vvY+hA/zTiaSYpO6OzORDXvhm4b
REZ57mcWoYLygPUhKz/ezZBJzP9+nlHn3FvXXHONP2vbOSwUP2aoGVfsMB4ymy+e
5h3qKqRtsebx4hf2uue7nGzdN4jnDp0zqHr/xdmRw8x0fCNmBhG3y86SrDbh+Li4
TrjSfvyMNIL1EeYTsH9Hk6UjW8dPxBLXUdVPhWngzeIIyMybq6j4uL6TqksVLFNA
XqMY8lnt0aGT5kipfp8rRnAUeui3Ze/qTf3TipWHZB1UJ1bi9VlwMvpJYZIXsSFs
mlFdoysmXR9S76ynh60JKs5muzgFq9ZPS+wN793KSLa+UAm4JRYA1NU9+UnngxNo
N+bJZIvo35wP8mMF6iGOumCxx/ZJaoz3bbrNbnccFwrglFgVM5U4VtJXQITdBG3B
3UnQYMQiu+Z3wii+KKdYA1hNVf8T2az33pOxqdhNr6ycu4GtisqpDrUlrGIx/DwG
fvT48DdknJ2godldokuh5PDxDrrmfo2LXGMjaqYjQNxbYXFPKJAYfZgptTiC/F1U
A32B9KvsBYLBIh6C4G2l48zxESnrEih/GXXG+tDKigCEP0Va8IaZYGR9pXpnoSWm
a3iSuJo+1KVccHYsTUeH1zpsS+T25XKAb8yHVSKsVjEK6B77+iDPnkicu74Bg8px
OkLb/dt7QGPD6KAGipG190Sd2ldgd/yj4Mha3c+fBKVuLYgKVu7fgAnRDc/Fax8Y
5NTnxzO6ceCwgjEXPyI+j6n6j4vwe8gC+oxh97eRZoIV6/75tp5AZwISNO5t+jWq
l6YTCerC5DkinTjAZkXlw8t+nMK4+DXQiSXLPwIcRxS2LU+iYhp+t9qoPm0chNCY
crtFWHwuMFAJflqbsCvLJvoinyOYvMmGCDeAoI961HEQp229hj0IYyQ99WXcEZbF
sKv9xVmVhWpJOcp6eR60fhyDWlEWkS+CmW9Y4LAr4d0K7YvsDehL4LSM/ne3rKWi
955C0xLgiteu7abEopH20bNcBRwWY98/CuXDBKcPEGzZryArNd8X324G4WlfuibX
YnwQug7rhWMuOW8SXwpqRWL8fpgmpdUstOJ3WPLkLRLF+7+MqRphlTw9g0oyOzKX
yrgl1J4xD98XAwQBKBYnr9lpBaFkRErii/bK0BcdF4BPQnlan2MCe4fdCLIKb6si
C4hqTARR+WIV7GdXyO6R2SqFPh0YFNQkNuE4bHwYuF76Ephf3TgHdsljdgCa4Drv
KNJ8qbVg69LSxulurTSeF6xY4cVZ0+t/V76fzz2Og9EYuCMqndJLAHV6X45A1KT6
979FJiBcr0jGVtTKgnbK+varFMLFn+304EYdFfUdk5lUG47vJBV3XEvoMZBXqLSs
J23pWR/DvtKjUNGks818DxYHn9BSrbBo9BlafZOqtw1ScxYDpXx+HjEapkOl6fG3
dLTtTwkjLh0Sy1H4O+vk0a7mMqb5yWiukasRtPXoI1+FvS/pkSZdV5n2YkRIXtlT
R9KRhsclf2est0QR6HXLfSfLcv8a8Bpx8HEFXt3Xl9FuoS35nZ81eDQn/CCbKapv
GEMHYKI2u6y6StDVLcvnNK/NknJDijesetFmtwk+ZvSb8aDUX9GT0xSK2sDacKgP
yNEgQ+D5S93VR/vMWsV5Zga9+Jjw1+Zre4MMVhSL4KstLVXckRJoRzGMCDXSVAnT
xvs7wgnsKz0hMobVwmyT1UO+7wPUealtTu0qfPsOIjmxoCcH+jaEl/gfx0lHqCAB
GIXxvSV5+TlSqc4d7Ls7bgXEYHTiloioT/OsbzlpimnfT24GJ3sYtdxatRulg/ls
BhuLe3hfk7xxZImydaUcldzKgxp383gcSEQ8vKQBaK1LePrl4d8vvc05CjI72Mvx
3qrUUszOiN8ndxnepCzN+x2FzyfyvC/VwmTdrTdyCQZxuEdLgtLjTcWgNc5yvgDV
6ElM74JTf0XX8BubgTaYNkvn+pU4LPW4TMAxzzUdD+KTn2vZWMCZE/jxJq0P3B1z
OD4AzYe+LLspOUdk9Ls+CtLLT10+/2Fm3UZw5OF8FpH0vc+mvv0bzSiudLyHafHC
wJfz8I9hJazJ/FYDm91uFh3WTcC+mCO3Ppt2qFOChQfnsD/SgS0aMSe1ztE+pj4e
ES8UaCTLSQpgzc5bRv/7lmQC/s+cqXDkPwKPEBAio5BFlPlenVFrsFEczKR4kyrA
xhGxb1aMvuN8nEb+LO61CsPzdE4K4XqoPQzJOawW1PMJS337PaUV7xORNgoJaiJL
/xg4T3Rbeobt2pvnubz9wYGZRiYMz/ulXbOiEM2tTdqx0pZ7DZzwcf8SvmKGq+KF
C/1TgQEdpmWnpV6cQMD6+UW50zNv2mb5GY07sv0fGXE0+oxzSvHwZRx1CqwyatVs
ONnCJVT6JnVM+PbNBUe4RKKhviFDD2NWxmF20k3KZbLRgA5ozfzAmnOcLTAPpGyZ
519yVAlfCIw9XcYIBK9TVxUnlpqJx2kDC4kT6ZYvXCyYTUEMlSL7H3/oyZPaGh4B
qomH6ObbCWEhGqslrePIG4lVqoD6Cs34UxkuXmvMLxADbnPMDlupLeBgXZ6Evwbu
kQsnRqo+1GhY8ZLwXmJw3odOwBkaeaeVUTqji/mJkzlish9RlRvaTS+7VjCb84AA
W18RviWce0F19KOMuO31rfE99gR3psCC7fnT4dXK6RZUw29hDIAXr/WaLJIOmDfm
BeyiseAkHb0g36UWUkcfQYn6UfRlsW0on+f1HA1w+gLhypFfE53d35TDLFEVz4dx
yrjlQPmfCjelx11UhUbj2b8ZhFIspLdCWpjoK2mWjQDb6Z15/xYiLjt39U0wxddj
dcy8H+/2ADM/xsmD5Jr5TcYFIJr2YwPdGobPiJ+0C4rvuqUYeN2mY0nboYUpEbsn
Ox8qvgd880ItNWrXcUyeeJsIMFDW+U5dLhncPm5qku8mPi4uX0u10Wydexy5wSU9
Tuj20NOzA2lm+ectwNMCKCs4dHG1e9JRLNVt+ASeF+uXaPbPdEktoenkfuAX0Cy8
syhMcCxsUZhOpeFIcPn3H76JoIuxgmi5OojLwJoKiBLJ1YHPndy03CWSiI9j0NnM
c0CmMKTrXiLl7iAXqqENKOqXkKgAJC8La9ZfMETd6m4tdMzcISmpmas7JJkTZJPy
7l0gqr1Xi1JpeAAkUlTlm6+87Zzfc5Ppzpp6onKm/qupYio85uJZog9Qz4emeGjj
jHdJ5MHSeTVedVUuCuuO+fFFOPCR/PCcLrzqKgZMqpxd/z8q7qBV3RKg0ctqpuJG
+xA8BSXvkUfQGzFtryMjtUjJCdSTVKoGwvmvID8SWfteZQu8PaSEfTcN4IssTvcu
+csYN3rrvwRZF3xmsFbc2JAHmgD2tlGcWJk6fffEloVuGf12j2kM2qoeOoTBpet1
Y1yzf12+QUvqfA6oVtDL+crH9bxuX0mkP0tMlsxvbQN05e1qttuRSi0S62K+nlQ7
TI8Z36OKPVVlHFsUoFNFCSfl+LzUJzQSlI/UmUG5H7BqRHaB5L/2n1zl+jl8ICj6
wli9Ngc9Q90Sy9BN5JFOwzZu6MR8GorzeCPXHKRalYEthiAgXnbQpmxlK4fzhmfu
3g3XrEfWXSt/9eJ0leo7foY+6UCcFRy76UzGnShi24b4i+k+XxasAbm9QaEXWiw5
IIOp67d5zmqDXBfmnAvN9N7kak7FmvhQyFb7IzvUED1zkU7zNmPGeZQqqEwZwskT
0X1Lg3oXWB6PHM1eZSZVb2cf0L4j0Q7DWbJvGGiFf7o9xXLFsXx+ocK81cuY5Zuu
pv6yr/K1luMF/vc+yIM1Y4f8lYviXs3iS7ICc0YScxNZt2sVeI071F5rX3IAFvie
FCi+KCLD/J80RYH4ly1ZBGpNHfmtCYEWWabVjqB+hC31ag69PH02yJFM68PzeAZz
oG2eG4sR8VpOyoSsWJNtLEHb+QsluQNF0VojQYQSY9kV12JAosZ8lq1nJ0RFIW/8
3P3NvZHR2DwZrbJc8t/9O947ryVZCfHjUHl3pScwnhPhmjECbCiYYSfl9muWRIzX
jaz5l7lvoYhDRWVu6q2h8w2j7owH4JQUz+bI7qKhwqhEufAEltFYXLBZIPQmU0oM
A6itwWmehT/oASOk22NuhCKXTUTWLN0hC16SfkQcWF7SXOGd0KhGxLbScYjYwAIN
wf+nnlirTQ69GYdiHu1lh6sZFq09DOgUGu6yTsgovaZKrvRxZ8jDf+XeTlMTApDW
hByuIkoB6KuT2tGSov3VZ+ovz6iL21jfqJ70xighUB4Sb0/LVcb3/x2bTTZ7tV3M
/ZIs3dL0tQO1dLh4gzLoAKAyI0qVdg+kWss/1Wlg5PwSEYAg6/nG2V787kJlaLLa
90X4+1nP50tiiSKKIkFxLBPkP9+gQj5ymHCqQiH+GCDIJA/N/zpBTeb5RQTZm1Rj
PkDWb3bT4hzEw4Go05Jb7stzLb0b0x83JT5vunoRP071qmCbipIQcM0CEulNc0vW
uMWQM9I4mNp3PP5s0attyg4xEsVvwdtzEA0QEPTTXTpkW/+UOGGhw7v0LW4N4if2
CbDPHaDHxy/H7y8/ZMoI7BOd6QWdm7Kr2sDMW+rm7eCPCRDNJUUZzrWewdYWTPo3
80SAYwJqQNobO3ua1lOwjff2kdv77ITPptB5sZObF1hpadFwmbkC18/MWy9FI33I
KWzeXKr9qu9wYtFGjQteh9e2gQY3vGUxqZtw62ychcFtDFtfyMs5WnwQk9aI7Tnm
DeQ9Ruqr933sfEJhwHpIex3kewKbCVupzWBjR9R8lvC9qmaub8wwB4bMEAb5twdr
gpfjKsdzX006QMDfgnGnCpd/EbNKp5/1n24/Ntf1JyQ/6ky7t6/22euA3rth+81t
j56C4ZGa+nq4XVjnwc+BAO2uEanSiyPFZxhi/cbljwpicJ/q4xfl1jFqFxK2/shu
9PeY28IfXym80d2AhXPmuQaL2oqKwrhQq7cFXq8Z01PMMQ47PSOpN5na1e2Co0o+
gnh3K10kbIDtqquspVDDkbzQLLepl/j/UQEPzS7IQlP0GwtIMx4I/Wt+HUgAikZH
QSLTA/U33nEL4c8to/gMpAEzchIh33uQ03O14HVWhfXYAdNL3Zcnr1COegUdCfiy
somnABr1YtArvx0FmhAALtP9e+nZ9o6CC1AODn7rop6DkAHnfUXIiGPsr+wDNkrN
9ES72CDdbrGoGHFZw2F3P5LB0OEfvrITuOpiJ6g/myNeK9gaCLRQqYy4F4ZBWvsL
pEmGAf9guEC2ZAX6+44WD34OR2DQAb+dgWXKKPLg24q+pafYpJ1/4s4ICkcSXvpK
s5Wj8WQSHUWNgwm9KXVB8l5QSophYl5o7OB2e09kKCOImej+bkyTA1tQOUxrWeKW
oOMevENq17IyKXimX7Iwiz/PFy8Mo3izEBYVrfL5HtEP2xgLjUKifFyQ0Nlqs2d1
Rx/GR7dPxsYrPIvc2qbRHXVTaiWfHtXfkrE2PpA2PVIoyRu2KtwegatMRgpPimoF
9qg3hJ+fZ7qiAKGtzQpRmfBuuAc+mZTYAPDDKueCIT1YuFvX5PvlHC267qkgg49m
KZzuEAChGIiwPqhatLiSURwnV6NLRWl17k5MLqtjG6jfM119CUofzgYPwAIZ7knh
Mfrxy2olrbbahO9diNN5LH0A7tLZi86qZ4FCNVkn1HYDFWFXJRTcPGyMXhYlaaqU
ME2N0fq9ZmcPe45Ft+Xzn7Hq8czvBdvIyemsmhEvJ7/bfoFh+HwC7reHEGmfoz2t
Vdsfo3PdXT7kXicyzVm0OFF/Hmrm2h3BhUyGTUfAuyW0KZLL5NwhZX7H0pwalFsT
M/ea+465PXJ0P/d4X24MBg6DA7px80yMIbV9FSLYZHOGcz6okgr0MPMZoEQOnmE1
cXJip9KdX99GuVv7YUnLQibAIW6Sey/kzAMmbYnEjYkSayuFb8z96hiiYTzZItaR
5uwYlC0CwqfVvfScVDItb4mqqAsmVbRStWRfs5ZTVm2ukIUfqswZ5lobXuTTzmvi
SRtJqsJHJZ9jpdBK4blGVTg5/rQOLoof4GqPE9de7FXo5KuDb06ufn4DKugWzfpo
zKqD7zJBJ57ty7Rq4VQNwaRouY10sHmkKyuyq2Sa+YgBzMiSgQKV8ij6eahox609
TLvOPwc1WUMFEQ49NEAPq/nExRWzz+WL7a+GgTy7znty05TYPNbvsExuc3p9JLCd
Up2PHPHAjLNp77kGWRHF5ifr7TVUcnJ7ghSxXeaSUOju1KcRfF1+J4/5iqIPSfHI
q7DEnj4Xtin2Olkr5sDpbMaFD4hZVoct8JjrcrQ49R1qqvF+qHIHf0IIvB7qjwsD
fA6/1DKefBO6eNzyVXK70ajxxgh1D/2WcWINTzGGkqNKPjyP7d73kO6ez6sKM4MR
F1vwHHlcQouafRsW9671OF+lFQqiKQlF2+M7UZ6YDMdc5vCIu7ASS3bNvc3deoYE
JIfR21RZ1nBXcjG6iawqW/7B0PAdc13LZSn+5Vy2qoHj5BYdiIlov1vslpZ4oOm6
g8qc7fHAxRr6YiEwcMxiJ8SGgBntSilM5KrWwogcr6kDYdKP3IchOmnWnmIh1XVt
aBaB3FVAqL4E67tKFDZegXe4OauTEcgdysz2rXs72EZ0ZXPSywFim5y4Atn0qXpF
bF9oFN2zlF4waQXqwskc4tynNzCpLUdR6Rnsx4urbAVjPhOUXr/nbcJ8GqKXK9l2
HojUFrdjqlHIiDERCrDQitB1gc4J0Fw+Oh6UodSM5PHMPlZxDhf9wdDNFtHwbI+X
waOjOnLWQJvRN66c6NmZrn8WVZWanLGs1Eew5ARBaol4o63sVFBtv78R1LInL5wC
gcexZe5UDlhddUJJHq2mHfrIQOJgr7q0moHZMbCbp0WS1vBjOYVb9J2vj8bKxzDP
SgJ8zj7OPF3b15rqzpMZsYLCwhUHTX3+OKREYB4ejX4grWLbwjIVV/9kwW/pVBn/
N/Js+C3e7iUUFHCyRh339Y+49hVGCIDGH263VQl3rae3XQBtnAamMccJ59WSj8Tc
GJWXut6F16bqXQz1MX2JUsxC+Xr9Obi4C8+4t7UQzw1VBZsVFx0iVfy2TreEwojr
eTJHLkGNnE/rxoWqXZICx/VxLtfRbLmq9qLYkSjwJlMGC4Pc+7C8rS/kNGB8pAUe
3WLGiM1vgK5/maC8RrHxWFM1Or9Nn3gMrzfBwN/RVUyKObaNZQ4cnkp7+qGgZqkf
RNuypvkwscHhkbRDorf4+p4YvZ4h/wrSMpTQt3va6DUjjZuqG6v0ytMuFuaVAw/n
D/kBQpLY0IsUouKP2oh18Ygc1s/U+Lq4iOpTfZ1B+Kk8nPox7kKpwkW5/V6zoJmH
wPX22ZXLRfmOsNdNMk+iwcc4TyAJVTe9KQ3weL4/+AJU8ZEzrjeeq2ds0AeMBB4f
cIOiKopeRDwWjizXzIaBtdJEvwYHs83jErVHE7ANBjxwBMLIU6DN8YhhfHM7secW
PK+YV/uFj55gxxLw1JatPSn+Sb0RJIXWwvRaON9FL+I56lIGZk54gqdVfxCc/rsA
SpCrWZ5OB43XHhxhAR3nyrvXb/EExZAQ5/l1m8SECl+TMLqMXgCZkn/RhVr+GO32
dj0f1OkiUewVM3k6zdfMP2hesloe6JRq+Ab9/Vm8LRzPKnqDFZHa8/AHuFrN8Wke
NrCCesn45I8+DNyAAf6W9hJf2Sq5RhI1TZCOA3TmQPfrgIAKVcM+hBp/ZUv+8bbB
SQKX70L+jJSPA7r7MxTwWRbE4n5iW/3e527v1jp5fforIqMAVZF7sHLRySthkIDZ
VrbNy0DYlqwNwehdU1uLd54eQUxGtJcOyAabT6vMCCd6zZf1RSmv9zBfRkDm8Mp1
KvjaXloOy0qvPIqO8Rj9Xy/hcgYDy6htjYfIDo3luXS7uff7oAMq/S+1D8NXAv9Y
a/p6E55kV2Sznx6zqOr4pRKMv/eUWOsUVLN0aZ5/Vs6GdfgzknTRZo/Dk804G81x
ksnBbLW0N4me28gaWhSNrI3L7eoqg37d0CDhH0OvudYc8rExsYuDlSvf3XJXp23v
dDhx2P6FnNjERtVjzeCcR9QZiME/llZU+nm6BpZ1rsQ40lblBZeg4hI/FRY2njcr
FZq5t3YITwpCMElGOUmsVed5os9rDM+6YN4UzRyuRQn5botwMgz1Q2/7r/lF0NY9
RJ93bH6YMMllk9+N1JAksxQV+5JHxeqn+tYfTyPkmG3FSS2auJkH/irQTOJNZCV9
t4azBEffOqzgjA/cJecSIxHBuVKz/FdIg9gDlIABmZKYPLIUGDuxKP55Q/BKRSbx
ei575p8P4RFDwXhIU3fU1l0QrDBA1wt3EWKIb5uszH/2gVG92FamUTV3LvDaidpA
bsLULwxhO/pJMY1s7Vbgyq4AWb+1nLTrQ0tXeiytaUnL0VVMgFpOQTP/lahfcHhi
+KBxWh1QWKgb3QvBYLrdvjZLVqJjHqJP/U7cfYZoD9u9Y6lyXp69XLXaBmeUh6sn
sbODjMQRg8R1mqYHab+EuJX/CbkUdLM9G9Z2irDnu5fx3VtwJF1my1PwKJ43fMHJ
97yJbmEXbjZMSPP5MToWpnq3pbfZrmazF1GiwSAID0c6Ak886YfuV0jdocCyoOE4
QwY1pRPeGHmvI8gZiG5VgYN/gu+vQjT4A4j0Ob3PCO2FQrJp3bdDU/ilnrnRramV
jjSD/BBJUgsvSsU08+GVWenJGfkXv3tCmPDwfpLo5qTshUZcW1JR0aayOYkzPNjh
XmauU6Yx0GG8f3M9FYnnLILxpf8Cod/cYpqJ3BAPilkiQbjsG+6j/o/4dFGBJteY
AEDBd8jYoNRPpBYvcEGbMz08vGI/iMfg2iMTtx3tfCWi2YCaNrjSP8ALVHTJxAcp
MOtAPMo9vo3fzjTqBKVnnm7Qv0shZepCKjYWGGxOgENvuM9l/Xo0lOYshf6biTmF
183yoYE+o6ndDSzRfw6Vwtn2w8tcBACL2arw59TgIfBH51+smyBI/QST0hQyQf3m
T6xTKQ9advkprv5Qcwg81hcm2AN1FC4VAJdVNu8mtg9ybunUyieRoSoHoN27tCdR
D0DR1Zr4gRCjkTwDw0Om8tNYsKpCYboKKQw2arG9aPg=
`pragma protect end_protected

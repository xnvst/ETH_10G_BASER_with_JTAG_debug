// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:43 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iWpmr+/wU7+UAcTBLFmgAronNDkAKv0Wu+yVaTGAsTbqpO2sBZQKgWzEj237OStG
7OZDspa74VA8UC6OwXSOl76bk0jvuHrXYh25UC4af8KFMT9xA/2mFprsnWsoirKH
UD8JLbasT5ORtzbIgO1rnDNfD1IXO9DjO4ObQJt9T+k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2416)
mWNlzGfpgMhLGe5b6+iLTkzMo8sRwvX8eDQ/cV9MlIhj6myjEtKm4w8eF3j8RdE/
fpw7qNMIQWi4JxbcFvGbWAZ9Dt3ZRSTSQ0eOrLM4WUgZirfWZlx+SgLq4spLxIwz
08LXN8TeqWWiykNubUhPqeeTg1Tu/nlTRmzg6QmijpMnemGM+dLQpEuMQt1TvYga
0g+DAI2YA4kO9ZpP0T1Amup+uqIqtze35U4r9UponcKx7fJdc3rnChCKBYasn30Q
IBamLzaV3lqmdy+kFN7AHxGEhRRpG6/OKHrDbARtXsb9khOdKvXZBA+rJKrEgAX7
zAV+euytozuLxxMqRDfrFHrTetXEpCrH4fttnzJm0iZcIEQ3HSeppqaIXw1zMPs8
FdfHYvabE2jmrjDuuC6IKPBKviKUMygRjoHG0di3MPkQuj9j3OuUbi6+gYZ2/EIb
gY3qzHdkPUQIZD8oR+hUfEo7FQ1tsIRhzFsxbcOxt5XwvblJ+kl2hFBGDQA/J8mn
yu1jxE+2rr3Tw4oRIaAPRfrmfCoBJ8GytOZ8astGIyZQjytSFxXvZXRMO3ybjO3G
F4z34So0h/nsnbeURsXInRRCN+t7CVckFPXfjcsAaocINJv6dYQ/EttGaK1iY1st
ycY+HIF8awzq19H+VulKDJzkZd7o1Oxse7K5dIKXOY2nGZfHJ6nyU6BccPaYpEOf
6ORLdlHQvbjEBDoVgvfdfaxmkh4KZ14/zgtsATsLr8Oj20yhBCbStVLhlbSKiQF2
zLOdw1E2YygwRDOhmiwUABHpm2iz8IDgHpX5Byt5UbI+kKGD/r26JqArJS9yOLe6
vM+se3yiigrLdbheWYvy/VFhK8eaLWnfwOigqayPOy2StYn/XkSyrKW5zznOD0B5
4J/U25Rrko6GuOX+5zlrWcuBPBMwIy8DV5SkPd5N5/ZlCPXRIYJ0GCQIxKCMiePg
Vm3gOESLuUzgntNGDOOQvnwv601ZFmxvdacnlIOv1t3s5J+qedqLF0Zl0VIDiicI
sLSfPAAZSUVvywvx3TB4tRMHiqT8Phk6n8mxJ4V8j8UQjW7VLZhjKaScqCX3N6u1
6gCvxLJjd+vtD4LIMkU36/37NTWUXmTxhUnUC+kqRG428+CRMYkVT6SYggFv3dth
PROU+05b5kfFS97q1Q6Jh/86Teuo5OxacS3ZsB8L9jFstHfmgB7oEuNxL8aPnmZO
3Xxh7YZo937Eh0gQ5YhRSrZD/q3v7qds0lp5XRZBHS5oXIOhe8I8gR23y8Jf/e5n
z8HymvypOZerRsjkU8M35vPShmr3fCU5Hdpuaw1dMIWFuOJz48hkiGMQE1CZfFJq
OW0nFlwzUvmM/xXDlsbHXLcoYi7sFtPDQnLf4w2pbDsEnJIYXM0jmR+ayg7JVnbs
jl/4vVSPUTTISFXXqJaLFwpHIRVrp7AigZ5LDKqgwZt7CDxa7gFHzhP6dSmzL3Jz
BFrDmKF+0YjqQ2OwlGw62gzzUftsddLDk8xzRT8XSC/3Eeq+Hw049y6L/4T9lzwq
c02B/SV51mcXDpGOS2ooxJWESwQCgVJR1mT7k+bp3XhFYp1oILuVceYMwnR1MIbK
fnS+JUG2zkfJXopxYLIjQH7yPTl1wVmWwmxUsV13CzKWZDmotH2RkN34d+DL4qOY
qKx5hAm2qg1evnnDUOkRK4EMCemn4UpCXeuLecgMMrikihBOu35AMEdtlzCi3YC8
TRIJLozNjxSIrOGAYgW3cPHox05WD5UIJTFzL1+/JZxG9cFaqAsnu89a97oCCxb4
ZOhoCimqOtqfSoLMZAQsTnvdFtrrtY78TBU0Fw9aScZ5Cv/hl+Y4UNn5E8ckRpZY
98Q82QYY7ysBzCOq89SDlk79aYckyVLPxwbp3q6s7P1RXFflRQhtUHn21UwUPWQU
P98NiECeApcS8uUsdAXFGb1hZ0q6sY/tLLbiV8m87waOGRaBtF5fvJDkP3n6qiNG
dKnz/kl0fPkQaBr8WFz40Rr2BibDO8v8K2dmTFXli0xf+OmTInYHGGUCSSwPFLU/
5akZF9YE4AaVOk4tcoy/ToGogRwrIoxIjkwmu+f9m8zt0/5rvvhOQ8q0QTDoykiY
HzvJyxpZHgJmc079D6embEWGztC1nRkylYzm0+66DCwFI/dX7ev0BWjAsCdXPRvm
/fvbP0zyM7wFJ6tu+r3zFok0J8UOsc3WnA4CrQabkOtPGqFdNtQns4gmTlOpEn+4
IiPUZEy2Dn9UUvGRraYAvqdw8fStAwjMDbYD9UBU0Kn37AHPFlkeLL6G1wc0Ssa+
xZBw1DKCDODkTMown7EA1rIWOcvl6VnCAYe6+39KisgXtYepalpL0i61ir+zUoJK
RFMICWrXkPazGnqTLNCYOnRpJmBlM+JUAsajMT2HAFqzICDMsO0jT2EtWcDpma1v
f6dX6GLsTwJg5QWoSFC73Qd1djonF9QRE6Sc7hfLVue7x7C4ESrELDqySruDpABe
KwEFYaF9v9vosXXDHToXjxvAvCP0buvUfawiTLaWtjp5NYfIEFYhcHE7SsNTzYBY
00ImqfMaApnCF5BuWWuS/4eFOvGsr4hpnGVSk3PNejCWtBbx4/UgemJJN0xxk/WP
IxpwT98bQWvUw8ggypjq0Bty+cLunKZY2FSBdFVykRf6lD5KBoUZNsckyzm6XhIW
aldThVoeVSBedoQsFM33juPalH7kjAWct8UoE8+niGIYN9t3n9N6SCM2tWN3Tp8e
IRO5GS1kvNxeDWTKZwdnj61hHde3tdq57imesyg9NwOEuHwiItC2QeVfuhvXYarq
LlHR47bgWgUl2eFW6pW/ZFIcEmlermSEYwy3vQcPwXByjkvTmngJipPh/b5Jqrs+
EJrD4KdozGSeKHEx4KNNxAHkm4xFbjY+gHUTgbQ/xJZSoUZ4bwoe/PI4u7p38qAl
IhI+uWOUU4B/suPUULHkXzzQkipZVyalYK1GZ9gRkQ5et0Lym2vyXbbD6oyEAXV+
gn9WUqjh7wg/JUKYMko71BIpkp2r26wqz+U11FG+xrvL5MLWkqMvoSq6RpaJjwzs
cqR4HmB6R4b/t3T1LeqaPSmv8s1FlkcnVA+jwmDV4DM5IG5I+VpzNbUvX+TWEVw1
8kqvpGoN+6ycgTwxBLaDXBwBk+yLbBKSCBQstxAP9q9pYLoqePq2ymrNly/xilF6
Z7Jrg51Kgi7f+FbfPoP4kA==
`pragma protect end_protected

// avalon_mon.v

// Generated using ACDS version 14.0 205 at 2014.10.10.08:30:57

`timescale 1 ps / 1 ps
module avalon_mon (
		input  wire        clk_clk,                    //          clk.clk
		input  wire        reset_reset_n,              //        reset.reset_n
		output wire        mm_bridge_s0_waitrequest,   // mm_bridge_s0.waitrequest
		output wire [31:0] mm_bridge_s0_readdata,      //             .readdata
		output wire        mm_bridge_s0_readdatavalid, //             .readdatavalid
		input  wire [0:0]  mm_bridge_s0_burstcount,    //             .burstcount
		input  wire [31:0] mm_bridge_s0_writedata,     //             .writedata
		input  wire [23:0] mm_bridge_s0_address,       //             .address
		input  wire        mm_bridge_s0_write,         //             .write
		input  wire        mm_bridge_s0_read,          //             .read
		input  wire [3:0]  mm_bridge_s0_byteenable,    //             .byteenable
		input  wire        mm_bridge_s0_debugaccess,    //             .debugaccess
		
		input  wire 		mac_rx_status_valid,    
		input  wire 		mac_rx_status_error,        
		input wire [39:0] 	mac_rx_status_data,    
		 
		input wire [63:0] 	avl_st_rx_data,           
		input wire 			avl_st_rx_valid,          
		input wire 			avl_st_rx_sop,            
		input wire 			avl_st_rx_eop,            
		input wire [2:0]  	avl_st_rx_empty,          
		input wire [5:0]  	avl_st_rx_error,          
		output wire   		avl_st_rx_ready,          
		input wire   		stop_mon,
		output wire 		mon_active,
		output wire  		mon_done,
		output wire   		mon_error		
	);

	wire   [0:0] mm_bridge_m0_burstcount;                          // mm_bridge:m0_burstcount -> mm_interconnect_0:mm_bridge_m0_burstcount
	wire         mm_bridge_m0_waitrequest;                         // mm_interconnect_0:mm_bridge_m0_waitrequest -> mm_bridge:m0_waitrequest
	wire  [23:0] mm_bridge_m0_address;                             // mm_bridge:m0_address -> mm_interconnect_0:mm_bridge_m0_address
	wire  [31:0] mm_bridge_m0_writedata;                           // mm_bridge:m0_writedata -> mm_interconnect_0:mm_bridge_m0_writedata
	wire         mm_bridge_m0_write;                               // mm_bridge:m0_write -> mm_interconnect_0:mm_bridge_m0_write
	wire         mm_bridge_m0_read;                                // mm_bridge:m0_read -> mm_interconnect_0:mm_bridge_m0_read
	wire  [31:0] mm_bridge_m0_readdata;                            // mm_interconnect_0:mm_bridge_m0_readdata -> mm_bridge:m0_readdata
	wire         mm_bridge_m0_debugaccess;                         // mm_bridge:m0_debugaccess -> mm_interconnect_0:mm_bridge_m0_debugaccess
	wire   [3:0] mm_bridge_m0_byteenable;                          // mm_bridge:m0_byteenable -> mm_interconnect_0:mm_bridge_m0_byteenable
	wire         mm_bridge_m0_readdatavalid;                       // mm_interconnect_0:mm_bridge_m0_readdatavalid -> mm_bridge:m0_readdatavalid
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect; // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable; // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [mm_bridge:reset, mm_interconnect_0:mm_bridge_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset]
	wire         rst_controller_reset_out_reset_req;               // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (24),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge (
		.clk              (clk_clk),                        //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mm_bridge_s0_waitrequest),       //    s0.waitrequest
		.s0_readdata      (mm_bridge_s0_readdata),          //      .readdata
		.s0_readdatavalid (mm_bridge_s0_readdatavalid),     //      .readdatavalid
		.s0_burstcount    (mm_bridge_s0_burstcount),        //      .burstcount
		.s0_writedata     (mm_bridge_s0_writedata),         //      .writedata
		.s0_address       (mm_bridge_s0_address),           //      .address
		.s0_write         (mm_bridge_s0_write),             //      .write
		.s0_read          (mm_bridge_s0_read),              //      .read
		.s0_byteenable    (mm_bridge_s0_byteenable),        //      .byteenable
		.s0_debugaccess   (mm_bridge_s0_debugaccess),       //      .debugaccess
		.m0_waitrequest   (mm_bridge_m0_waitrequest),       //    m0.waitrequest
		.m0_readdata      (mm_bridge_m0_readdata),          //      .readdata
		.m0_readdatavalid (mm_bridge_m0_readdatavalid),     //      .readdatavalid
		.m0_burstcount    (mm_bridge_m0_burstcount),        //      .burstcount
		.m0_writedata     (mm_bridge_m0_writedata),         //      .writedata
		.m0_address       (mm_bridge_m0_address),           //      .address
		.m0_write         (mm_bridge_m0_write),             //      .write
		.m0_read          (mm_bridge_m0_read),              //      .read
		.m0_byteenable    (mm_bridge_m0_byteenable),        //      .byteenable
		.m0_debugaccess   (mm_bridge_m0_debugaccess)        //      .debugaccess
	);

	avalon_mon_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),                //       .reset_req
		
		.mac_rx_status_valid 		(mac_rx_status_valid),    
		.mac_rx_status_error 		(mac_rx_status_error),      
		.mac_rx_status_data 		(mac_rx_status_data),    	 
		.avalon_st_rx_data 			(avl_st_rx_data),           
		.avalon_st_rx_valid 		(avl_st_rx_valid),          
		.avalon_st_rx_sop 			(avl_st_rx_sop),            
		.avalon_st_rx_eop 			(avl_st_rx_eop),            
		.avalon_st_rx_empty  		(avl_st_rx_empty),          
		.avalon_st_rx_error  		(avl_st_rx_error),          
		.avalon_st_rx_ready   		(avl_st_rx_ready),          
		.stop_mon   				(stop_mon),
		.mon_active 		 		(mon_active),
		.mon_done  					(mon_done),
		.mon_error   				(mon_error)		
	);

	avalon_mon_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                               (clk_clk),                                          //                             clk_0_clk.clk
		.mm_bridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // mm_bridge_reset_reset_bridge_in_reset.reset
		.mm_bridge_m0_address                        (mm_bridge_m0_address),                             //                          mm_bridge_m0.address
		.mm_bridge_m0_waitrequest                    (mm_bridge_m0_waitrequest),                         //                                      .waitrequest
		.mm_bridge_m0_burstcount                     (mm_bridge_m0_burstcount),                          //                                      .burstcount
		.mm_bridge_m0_byteenable                     (mm_bridge_m0_byteenable),                          //                                      .byteenable
		.mm_bridge_m0_read                           (mm_bridge_m0_read),                                //                                      .read
		.mm_bridge_m0_readdata                       (mm_bridge_m0_readdata),                            //                                      .readdata
		.mm_bridge_m0_readdatavalid                  (mm_bridge_m0_readdatavalid),                       //                                      .readdatavalid
		.mm_bridge_m0_write                          (mm_bridge_m0_write),                               //                                      .write
		.mm_bridge_m0_writedata                      (mm_bridge_m0_writedata),                           //                                      .writedata
		.mm_bridge_m0_debugaccess                    (mm_bridge_m0_debugaccess),                         //                                      .debugaccess
		.onchip_memory2_0_s1_address                 (mm_interconnect_0_onchip_memory2_0_s1_address),    //                   onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                   (mm_interconnect_0_onchip_memory2_0_s1_write),      //                                      .write
		.onchip_memory2_0_s1_readdata                (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //                                      .readdata
		.onchip_memory2_0_s1_writedata               (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //                                      .writedata
		.onchip_memory2_0_s1_byteenable              (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //                                      .byteenable
		.onchip_memory2_0_s1_chipselect              (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //                                      .chipselect
		.onchip_memory2_0_s1_clken                   (mm_interconnect_0_onchip_memory2_0_s1_clken)       //                                      .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO���6��6.8Y��5�|-�EV$�q�)�Qj=�(T���ɣ��ϱ�@�͆D/���s��Vun�*D�%��g��ͣ&��Kjb?���n$�hn�!2��XX.`���Z����j�x���5�$�x��8�x0A�N\�9e�<���Q�Y��q����kT�Sn���z]u�n� 
�fgH��
���$�x8^��;�eɇ�2�_��f<� _�n����Ĕl@ˉ�����0#/�;�����吪����ے!q	�c��o�o��:*л6��V����Nqj���^�בgI?�l��B�ICO�[�庐��'����[�\���-�,�	���|�we������a6iM��E���X��vb��EX^�M�i���<�Gx��icFX,GwDR嶙N^R5l7��@�	�����?,,��h�s$}��x�c�I���U��߉�+�"�w��U*s&�DH8�y�Ȍk��;��+K��ddqj�i�ӭ(/]\��Fn�A���W7�|c��U/yDV^K\6�������q!h�cl��T��;�E����*]�T�����" 8u2� ���I<�d�N���{���^��:4�e@S�2����jζ}W\��Ø��o�r�������	��)�#5q����&4��'�:x_GM����N������`X��+� �,���J��F��A.9Bq���S*(p �i{��g֪��+�yLՀnE.�0��fs}�y�ԙu76?|���r�j���D���5��1)����Ӻ�  M����?�TQ���D���34�T�=��lt{�v��M�
�ʰ��77mc��~KL1 �����a��2�3�gBe=�~fP���������fK�����^>¯���࣪�q�db�����KsV�摳�#z�=d�	�'bw غ��~~�W���M���;12J��X�W`<9L'�K�@�R��t����K�\
F��Ψ�=$�==�KL��hT M3����t�"�m*:��u]�,�t��S�r[u!�b$� E�iE
W�5�YL�)����k'�۰i��/����(,2:�M���zܵS5a]�N�ټ��}�75�!HT��4���h���i���� ����c�����%]y��gLe�Ʃ}᦮2�m�uBS��A�j���d�U��A�?��1pԙ�W�X݆�)�{�T[�;<ɗ+�n�Ro���^H�>�ʦ"�cL�@�e�����\Ⱬ,��U^\s�nu5��J�6�O�$�K̥N�����@@�;)k�U�c��N�B'��45�|*�u�)��	A9!Ę�>�)n{�� J�%�	ANǴ��
r��r>�Sb�%�y�=���i�s܊ ���ڷ>�s��je�d�&�s�mNBw/��}��ƫ�����
�7 z�L+8�^��P6vڿ���r*ą����3�&	
=-+4��)0���Pd��v�B�,�ɪ��i2O��gNzG��:5��"�;nnm�fj���vC��{>y��� u@�4��,�L���~��_�L���S�ٽ ��M�"�@��c�Ί��&�<0E���>P��b�7E޴���>�H; s��᦭G�N��L�S�H�}��|*��xWς�NW���:�`Ӿ(�Y�V���(�CFND�6 ����m5C�*��;��쿤#����Ѹ.�z�� �����^��/]�c��.�+�o���
N��YH�v;s�p����d��mG״�M��'ذ�e}1��҇�+��&〥c�,����N���%������.Yf�	@Jxo���Ru�6Դ�?�AH�� 4"갤�� ����V�q�CP��}��hH�K��<"8!��ھ<J�*ݣe����G��pӀ^1Wv�s�����a]�L��J������1��\�L}$��:�
�UEΘw��)pdʨkw�g�.�u1�#���흣��k�Z���eqVE�L��)�T�ƭ���A�V)?.M�'����EF";�-R��͘�S��c")[���	��j4�ޠ}��@L|��B��Ƨi܍����YAP�nm#r]�ʶ��RKa�F{\�V�CK���I8需#R5Ļ�[�('�����RN�K��[x��
�Q�'�NQ��T���{��1�����Q����K��\��eH�����{*�]/���Y�M��)K���������`1
�5B�̇j���	�
ejFd��n�55e#�?T�޶6�a�#��"E,Pӽ���+�?.VqJc�n����"y�K��Kt�6�xi���rA���ki�NyЄ�V�ѿ4� 갮�GԬ9�OÛ)ĩ��������6�c������7y8�N�A��)Q�y!Yht/��*��P
�T��H/KfHZ�������:]�V��6eT�!��������b>8%�q�Z5�z	.��$9�l���qd�gV�<k��^Iz6�נ�^/һ�|����h��"��q���	5�o>2�� t�?�(���5^�=5H�_���^�M���o�͸�q���Ry~[���|ԔT��<֍�Z������@]d�Q) �[׃"�Ψ�&G�z�2�)e�>���
N�!>2D|��O�9ۿ
s����L��x��r �t0����|b��]R�tȓ&$�r����[���b�|����u�����)|�S�tb���,`ESUM9��z��v�9�e$&p��f)��Ϣ&��r4
�S>Zz�}��,�`{�*���lGS�3D����24�
C�D-��Y�� CE�u�����Eū���3�!*�Q�X��[�2يf�|�#��G:��++=�N?��W�_�����9d8����B��Л��H�J�}�$��9�O;�g��C���hu���(���sߔ�P��}5'��T�U��
U�FS�W�{oK�a�E���Z���[)�Xr�5�xRIÕ���X?��ZC5���531E��U β��3�~ӋTx�����'�L� �A�s���X��C��p�p��CT�g�JaG
	��,�#�I�W�l8�c=�S�iwu�u��m����c�C2�	_=BmG-�m�J�)����jnT��Ɖ�4k�:�����f�'���L9&�l{�������AQE@��2�%������ h�u�P���<��lr�/�qt�`�\9���>%u���ur&�S���2��9�[��҆f���u�e��s�g�]�u�A#���y�S�z��+�C,�A��=!��'�����Kt0��2z��A�!�[NEn��!k@Ș�<��D��vq�6/X�m��[�!ȷj���	/��[P�'������٦O&Z�e��?WL��_	�ȍ39͔0�r����z�8���}��i����S�4���c��g�ɻ�J�#<��nn}g8���1���+�r���x7�i����e����L�E1���̇r�!����i��7��r�S�z4MJA�јP��M�dM��P���!k:M�X�ΰ8^6ĩ��_A�!+�����2��;�;X�;�y�`re�Q&ŰʚZ��)�e�0�ɧpN,>p1��m:�֏qQŮ@`I�Ǧ�<�t n�!��<y�?�X>!���_��A�P8W̎��*����D�`P�c��9�(������k��za����v ��_ُ>i[ǎ�DH�J�������cYo���"��_���2�`�=��mɎ!]�.��d��.ȑUZ�&�����>Ij��F�w� �g��+{ES2%��v����|�0@��*��P����#�sm`���ǿI�����8�U�QNJ+qAn�$��d�b;�q�?��|5�3ţ���&���c�{��C�os'���~/���ߌ<��E_+�&a8d�	��8ؘv�z>ҧqݬ�LBՒC�Ns���&I�Mgع+4�����������u�J
X\�c�qB�ϩ��gGXͺ�ԁ��N�s���?Av$��8��!9Ӯ��Dz?x�\��,�����s�y�2��4Y7�+F�-���d �?0>��}�#�Rx�S�$�er*t/xӋ�R)��M���#����l@}�8̚�4j�BM}�Aٯ>WZ��-P-�/���r��zB�vu��q^H^��݊��%��1�8�(ܸ*2��p��kԪlz��A�}.,�L)d����j��/S�"�GJe	c��#�B^�h�
���,�jt�Fy���E�W���>�����-�|�8pn<ˎ
���߽u,��0��C�x5��9�#�RL����[?5��:N|�u~6FS-�{�>�.OMYc�]Q�)c��lY�G��q`%���
�(�X��+��V��Ŏ�+&�Q�"�D��5�Q�g5X�=a���dfN��1_fi|@9�-�(��I�&�A��W�v��wt�lW�]feE"+wy�Zf���4�]��B�Lh	���N�a�,���Dn|��'>3�$���*��&$֚�pȉ�`��Eݩo|+�.uv�Q���/����'�mvϩ$fZ8�����^���I�d+�����~�dѼ}�)AƖ�DcW�Ĥ�^��X�M9ɕ�Ry����t����ڷz���e�T�C��j��}f���L��8e4�V��.s�H���o9-�x�9m��%ER4��PtcUx�9�5��M�f4�t�s��
�����.XȂ�F�do�${�Ĭ�C����c:?_��V7�5�#(���*�|��Xr�-6p5�E+뮐"g�H�%j~e�Z��#��ǆ�arn�0{'��,�*?�&u$��j6�X��}�]d��qc˂Z���xӧ�ح�K�rfVG�'���;�J���=�䗳p(Q|��dGH�Đ���+s���q���A�V�O�OtjȤ}=d�hX@GF�U])���h���=�.���G���` �;@b�5*qՇ��߯��R�3G�Ÿ��2�U0)���I�7+Y����,(�{�,6��מ.�nV,���\���()����[���^�{��! ������k '?�Ғȉ�N�>�����q��m`3��$���5���=!x��[{!cn��Gm!�~�A�D�{�P����o�?�ʍ�2Q��@v�k��e0�< �/ԙ�7���B�T�W�V͐��e�5G8wabe�.2���.�[��u�?�?I"N7�;w��sl|�%:*#i����=]F��q�D?��u�V}J�9����^3:`wF���)���}&y찪7��T�c ��B1�_��qڰ/�#o��n��I-zUy�(8-�u��
����C��7�o�g̍��`�8�Y��Gi��Cn�a���x�q��L=�X�m�Ľ�7u�E񤸞#5��zmV\@dC�\��V�)���?��0�S����U����y���IN����ו�nڭi�º��%���4�W�����J��T�7�x��s��ܛ�΢�!6����.'��7��x�Ѡ	F�Ռ��G5�}ЯX��îW�U®ge��QZ�ŀT�"Us+K��io���;(���z�e�<�X�,�7J���硑P�-�?b����0Gg�B��k0Q��#�'u&O*˺/� �����?����E:�9CMl�5�=#o7!R�I	���M�p;�e�ت�!����X#����� ��<�u�Vq��=(HqԢ�K���C�J��!����<�?KQ��Eı���vW;�jZc����qim'�f7�o�06$�z�����f��vL`�)s���K�I�hi��.���#�tDw턺���Q��O�9+�)��
��#�E�p)*'��<�K���>��n;��TT�EF�?��b)�chGm��vRqpk*����w�7v\��k2F�Qa�o\C+������7�������0��n��!C_����g�Y^fR��+�����8:�g>�ơ��1	O߀4���Z�m]u��Eb����^�&e[�x�tq�c3�x��gn�W�z £kz"�ZzI����,#�:�.�*s�r��Tؤ��ٯ�n
�V���0�)��P��	�}G���=��&��E=r0�D8Ikyc�4�>�l,�A��\>�e�S�P	�M(*�n��he�[r���/B�Lf�1�v�:�)�����L�q+lk�Ơ�@dvtu�`QoNt�hb�&H` .�:��vc��TO2�"#sk5q�H����g�_��x��մ�����"���D���VQo�ȓ�+��6]��.�9�VSb�0C� 'SAX��BX��Ϸ�ԯ��F�s��+vCo:ѻ �rC���TI�^xV�<���� Y�}w�&��c�����]�K7Z��-��.)S�Fd�G�"P^����<si���(��:�=��n��A'�U%�+ۻX���)WP��?b����Eb�6
�,���q�I^[c C��oeO��FW��0�Hc(!��0�j'b��ٺ���?�N�py�J9(U�qV?�;=e�KǳHT�rF�j�8�R�L�4�n�^��&����ж_=�a��y�j�5�C�r�CԾs�S��i��N�F�QB���C`(��欩��켊�JeD�C�mY8;�0��������1�J1)h����+�y�b[W���G'H��)jr����q��2%I��H�!�V�|���f�(�;�s�s͂��d��_o��"��z�ӧ#c;&J���k����I*(������kŋ�h�t��X��{%���-f�%!����Ԗ[�n�pW�Ҽ	�>��i�L���=nP�~S,��#6v�,N�]�to\�7C�ѝ�[�\�XW��F����ן
��<dP̞��WFo��' �]K[�\N�ܝc ��v5��w�ԃHuK�����Kvf�(���P=@�?#(kq��l�)w�!��P&�=�#�VQ����;��}TCq �V�Β[�Q� `�"��X���Y5�08�9>��\��ڎ�xq{�0e2`6��f�ӑ���}}U����ZI�{���Pe��u)���KCX`���K�%���v3\@������.����Tq���*�p��.+��c�Lgi)����zcd�i.�x���K3O�j�-����`���@;.:�ȯ��ԝC��m:�df�,I��������̈���j�O�p�q�=�g��{6��HbM�ςź�Cq�`^u��Q ,Q�x��p=�*��^h���X���}����E����
vo��n�X�(o��$�hM��h6�h�w�'�}ץ�G�_6^{m.l-���А �_�p�F��y
��;��)�r��G=��i*���5̈v�"]!�5�As����Y�Y`h�j;��{B�� ��$��^۸<��H;rZl�X懲�.$�ub���Po��g��yX�T𢣛*7�ek���8��D�uXT�Ō\��M���f&�3��!�����8�Zm`�Y�h?zA�������5Q������=�"�oIEj�lSF�v��.�C��gtAq�VC�����׌�S�KLЯ��R�;������z9�V�͐$��RaPذ����?�Zj�b�Ɓ�¡t�bs�N�;�:{j{R�L�M=>��;�s�' pꉎ�+��;dxʉz�����w���J�A:z�L�H� �!��"b
f�����˴�1}�0���]{9�8'�㊁C�ه)�F�ٵ�}aR�i���D�?|b���+R���<z`�fH$e$�!�\���VA2�����A{c��Օ��Ӂ�{Er�^�gŊq�EQ)�e�*B�R%��a�G���a���2H�Yc�`p�Ϲؒ� ��q1�V^>��`�aN�0�3�N�d8V���X�q���:��lc��1��Mш(!�
vc��������_S�}��wK�W�ף�9��͒���V��y\��]�.���+�*���؇AS����ko��+ʏΧ�ZD��C@9�q�u���ط�0�RQ _M�I��e�X� �ryo��zJM��_6[w�4���B�Lh�'dYQ�_ήʈ�ƨW��/�_>�4��sڌ ׽'{`l��{z_n(��Mu9��C����#�W/���x���[|8w���Es< ,�?�ف���D��:�o`+��= ?�x<��myˉ��l�Sc�˶�D�=�&�g$����x~�?�^��R@����-8�Tʦ��� ���ō��벿������|�Ȱ�h��c���G����m���A�V�0!fJ뺚��~��T�֢���S�\�{�ke)��ʖ��x������p�Q;�T�mc��Ԗ�>Y�s�wyYv4����
�o�e(t��}R�(P
���N�ٗ\�� ��9(�,� �%y��q�h��"����4	Ds��k��G&|j+��b�����Οf�a��>c�F��l�̃sl�:6i��'Ah�ݢ�����ȩ�'=���-�n�:E�Ț{]�ޭ�L���ME�2����;�Iu~����ѷ����Rz���lxz{�y�Ho]']p9�XE��%�>��^�>1��O5�u�c6>"n�|�-Q8,�Zi��^�I�LXcȰ�S�c�b7���瀙+Ǌ�;hG��AK�Gi����	D-�ŝW=�
KN\h�-�4�Vݔ�b#_�OԘ�ؽ�@p�b�%Ͱ2�̃8�ޜ�B��B��bB���KTnW��¦�]��}vPf��-�����5 ��v���us������:WO�Y�Qhd�ђ�X��~�7��,W��;6΁�)B���U���x@�SY�m���t~����O�TP�0DT��N��[eq�	�a�O��c�����P����� s��@���{�!�Fx�T|Cn��;��;3[2s���f�~�@jN���{3|ި8�){e��`'q�+Z4Y�M�c�s�J�Q]t��'~%z���>	��_��
[�4v7�_��]���s��**�)��ĈG�����F79��>���@5�q����{�^2V��9d�}���R<ʉg��
�6^Q�E�C{:#�ޔ�g�	'|�P�,qÙ�~��z�-S�\*{���iV=M�[����i�,��k��l\�������B|mr�Q�>�������
��"�!��E�XS>�"ˬ.M��0e�z�}�����T�A]{`;�EM{������X����/�@��N�Kg�q�&,w��]�n�)"{�N;"���a���>|u�����? o�x���3�|��Y�XtI����G2��!�9Xg�d�~����7Y��`�Է���``D��?^�r��uy�"��F�k�0��l���H7^'X��_�Š p1++״���l^���)�����`y���vs�:�q��s�¢\a�t!���=��R���Xb�f��(E�>�ݟ=w�~�Csb��a���������Π+��Y��BLN=J�3��.K�,��N���̧T�wE��6�ɤ-���(͖�F� �J�l_�������A�pg(�n?���+$��������Ee��?�T�0����H�&<�f73Bʳ}���[�_���@�ާ�ڿ2	�c���K����8�J��:�<lu��F@�a�'���n��b���JO�,t��+�
p0������A���.@��b9��F+^��O���&�
�bX֖�o5��ܸ`�2�=#�z!��V3��k��Ѓ�N���f�<u�ڒ�a�N�.X{Y�O�} �B!�0e�A���z��-�us9W�3���BS�v[��Q����E����Q��R��}�����X�R��f�Þ�PR�I>�5ݰ�[P�t=K��o+�;w��H�$ts9U#`,@c���5�qif��B:h�g����ظth� ��qw�
���l�gm����l}�`��Aj{�B���Fb�R��ݣ[ކca�֛>K:�Vx�-f֊N���Mm���^��y^���L��~O�6��l�ߚa\�f�p�����D��H���{u8����AkPh{�[�0AO�H����y��[��"�B)vf����1�H�M�R6�z���К��n7��yc��.S��J�z��9�X�E\��(G���١w��׀ϼQ�Z��k�&K�ʼP��L [�+��`)��,����!Y�7�M�%]L :`pn<�U�f�!{G�`mO�Y%�}�pr���q��DF:�kYE��˶����[�,�Ro{Z�&56�{;xy�Oy��S�����?�Q�T��B��/L�V� ��^��g�>���aϢ~ဥK��2zI#�/��j����w�`t�'�F����J�Ip���Ă\�C�p�j��2Y�\��)ùۏ�4�V^K�S�)���ͬ�~��dQh`}VN"�C����V+�%/��ւվ���}� 
EH��C-�?��o�#KI����<�X�d�Ӕ�y��`0��8v���r�`Q>����BWJ"z��q��#e-@��*�,�����Z��J����.�N81_�P�Ê{��B���a�#�ߺ�Q�zWluf⛵6I��E�kG��y�A��՜�2�ڳ���`vj�����M�)l3-�ا��0�p�b��k�G��چ}S��v7�y�d�lK✰PS��j �w�.�o�NE
�f}���g�9�M�L�ylơ�t�T��;K���S$1�Ot�a̞�_K?�1�7!��puYNs�b|��R1����(|�n��zH��o��s�Y�vh�������%!��t�k�[��
�f�'��`�C��>�~n�T�Fs#`�[p�)�S3
*k��� ��t}�4�xi�Rś5,w��!��3ؔPTԤ�9	&Ҹ�ũ>��;&�s�v!1�͕�I�^��uU؇Q3A����T6��M�v�'��a�Y[_��t�H$�U��j�y�Xg��D����&]ǔ���c^�[�h�Z�d������jm/�v'6�f{Q��89����G.�`�	�bf����.o�6��`��<$۞�Ɋ�"���e΀�d<@Sȉ�)+Y"�	{����V �[ɯ\�Q;�6ۛ����J-1��?���cs�P�����7�ݵ���{W���?E�ۮ��T��i�یa a�)ǹ�H��]n��7�p��(�EZǛ���"'T�����Ǡ<y��U5�d�R�Md"u��Q��햆�Zuq�=5�$`�+�����}e�x���F�7+�����.eS��BЖF����:1��z:�I2�.C�X/j�+#��������0�ܘݳQ�o�*����O����0)�H�X: -�m��������� ��˸V��gm��fv�G]�~�VAE��uJZ˿�
󇡃�]-Pq�e�|�p:y3,o�߹��`sD�BZ,c����c�E��aqo�]�x����L�[��Ŵ��qco
,_�>LD&�.֏����$]EVG�׼Dgu��.�|����z/��nD{b�X5��Ǽ^dz��6�Q�ҏL������Q�|�i�f��a�c�@���"������r~R��w��߈y�H"�$LMD�ey77��*%�W����d��g\��6z#X,��f�y�����;�?�"�,�Ǜ��$�����(�\ˋ�3���&���L9�N��:��O��$%�r¾�a}a�h,���v=5�t�C����P<�`�z�j�82���Y_���vk��O�?w�̻2	<r��D��x����������5	$pȀ��B:��!�������;v�?�ʶ��Zf�vC$�_8��i���oY�1e%���5�b�٬�I�[&���cy��Xߢ?Z�T��L��zÆ6���۰�)�G/�(Y�^��T>��7~Y���Ռ�^�\I�t/��;�
H>���3�g�q(�0A�3�Qxm�'V�K�%��@=6p	���Za���c�2zyݛ�Ț��I�Ræ1\�_���������A�\4��,���i)3����
�
;�0`�f����P���~�~��?+��	��?�O?��)�#���a* r�Tto��(��|o%�Ym�����Ug�����D�\W˃�,�ɻ-��.��?�"&VdR����c5Q�Y\ ���(J�Y1L���i�����Z B�X�[-$�Z	>5�wY�Ɓ��VQ�f����$Ql��}���#���
[/�"xjS�M��7OԂ�L�Є��>�yU��BW�/�&=  ������><�����})=0���c��'%Z�`���u�0K�;|pv����r*Bēb(���[fc��H���7���#oҒ�O���+�#��՞&��;#M��鋍���kɿ��$9�v����(��.�z�&-z̄��b_��	Z�+�iR��^�oUB������֠&��NbT�N#�c�UfH�}�\���C�҂��:�vEݮn�
�h�<��t�&L$�Tp��@ �ǲ�� ���h���oi��.c��޷h��~ w��D,�.�.�!�A]Mͱy̘0��х� K&������A��Rs~4�5�!��aeǶ�`^��"�~S��@�����+�b���8h�Xlo�v��" ��. -�9�"TOonw�tAadىs�C�����U�ŁX��`׋l["u�-��T�g:K$E�l��҇;��4[O��a���FA��!�|�}�y��8��O�H.$���M��+�����&U��tg3�]���?�{�ڽ�;~p����䁩at����?Z� u)��+�4���j%O���BZ�<z�*��M�b�h���T"|X�����>��S�Oc�=���z	�xC�(�e�_U^f64��J.蟍6�/Ʒ�P�c��3�*v��u7�0M$E��)�ec�z�1�bL��0=kf���V���S3�SE�|����W Ͼ&�D�W$�MHNrW���mZ��(����g��N�mɶt�
|:t�:�_� �⻮9����R_W��`ƅ�UƷf
qNd�D�ɩ�u��`��*�!�B ��cC9��
F%5L:|+�!���Wp�g�A�&Qh0 �-���Qa�YwA�BY�6��5m�g������)��Mm%�'�#�%�z�WjGd)ZPP%(G�Er0��bN�#��I���͇��'��ĵH6E0)�����������ߏ�@:��C��al�Ms��}i�_��&?��6��xDI��/�����P�-KɐeLt�7�	�t�-&y&9 ��'��r���6-s�����r���d���g�-\WY�џV�˽��*F�M-��qS��'����n��?���_%*'�K��8�~�t㬅彵���).���+�%w��[��_�r]'^x�48����J�S���	P�#�#s��G'7<Q��',_כ"�0�hP����	@�����:�����1R�M�1�L���D���L��9�*��%˫t��=�/�x���s��׫뱶;m`�4���D���B�p��c����๧�/ �;����-7d?iwަGfBS�FV��D��87��zGF.�/�/ wE�Į����՛�@]���N����:#�Յ�)��ч��
��P]L�����*ד�K�͑ly���yx> �Z�8��z��{-C�=��,ie4�M���hh�Nl-�!{�ہ�������/���U Ɉs�k ��:Q�|�.Wy��s�A�F��`��|h���M m��Հ�*#�҃S0������[>�|�ņ�I�[�Ȉ�h��P(��b>�f.�oX�V��0p��5�,+驔n�QuM)�ț�:���*��W������b>S/ �x>;cil�՜oV�v��W�Ch3fc�I��_�/��B��S�N���x�Y����F�ʃ0����)��Yo��:b;ț��L9�R���P<���(J�_2:����DdU��}�$3��Ҽؖ�j�B��������s�C*�"'/7 /�ˉ��w�!}��X"�A�V�06�K��A(���7�P�.�B�&�O]x��e�9����%xR��t%5cm*��|
DHj� �r;qǩz���ӀiWrCy5C��6�w��h�$arK/&Ү�"Y�V�"������C+AS�A8R�y.�j��<��o`��,��#ϱ�	���t*0��+��O�O��"!�dz嶾�L�v�9�QU�k�#/��|nE��Q=1�&�:�9d>T��y�V�`����Y�hw�7eZ��f���M�Շ8��]�!�+�&��H>b;ެ��u#�Q�m`+��6Ɏc�B5�.TV3�A��;'0�� qc�3��6���Qx���t����%���o'�2Z_"�c������e9ĩ/R�M>R������G��l��j^�c'��iz-Qt�hω�A��U-�Ş��O���x<<~�Bz����X�u�#(ys���)R�،H�r��_p,[���%9����Z��Hx?f�X����/<��q�_4J��u��V(}�$E�_�����R���B�c�˒���������^$�>.|[�����h�1@@��Iϛ��:��!�\dyA������D��?���ou��)���\�ﾇ����׈*�E��,S�C�Ũ��Ee��Қ,$p������$�d��<��K��X{����oCy{����O�����O3��e�k��-*3��Ԡ�m��ǯ4�Fe�E����hƮxXI�oJ�
�!"��!	���T�p ��+�岦��9��� <Ù�J��+R���G�f���u�T��.EUb$����-�l�p���G
�A=�&����[�ȫ���2�z)�;`ڎ�_ʏI�_��[	ua_�Vyɏ�؄<������T���[=ҍW��$��Ŗ�P����A�m#yʮ�s*�j>�a��'��S����F�7�/,�\�Y�$���'%�)94;��Ӱ�1)|��o�hIn �(�ǣ���3eR�Y����^;�9�:��z1s^�ˁ�C�r���P%<�u�婷f��I7�Źd�cFо�X�:�ē
�o/S�&]��"�{�������:�q�|Qm���Y������@��H��_�/M'�9�;,���0]�S��X�87���#(}>M�ٿ��lڐAH��e~�Yg8�7���IS��zghr�0v��	�V������#-ۜ-�)�P=?�k��6\�4xKy��������v}�� pN�1�v�R"����*ĝ&$�_�֨D�B�Cou��*2�Խ;�Xeh��(����s��ge8L�6�[Y�:BnK ŉgY�N�u�ab�9�'=�0�2��*���NW�MJ�	�	��H�b�pxμ��
�b�$�Ǧ�A�B�(�tUǪҨ���v\���WˉX�^�SM��Pv6�N(�c��j6�/�wS�9�>�zgsF�1�$�(������[�:NA�c�+Ĳ�A�H���qî��Q7��l��C� ��0U浢�LӕW	2Fg�!�*Hp�n�q�Y�\C�v��i�{�Z�S��B��/� ���M��R<Q�bRoרp7���s ݳ�7� M�
xcGN�����p���{-e�4�Zb/��U������^a�!��:�e��l�ԷX��� ����I�@=O�V$ͽ�L=����Hd.��f���U�#�!a@
8�;��n��&� ~*K��Ϛj�rU}�+.�/�չ�'<�G��
RZ8ބԠ�3�7^���7�%���*���@�[��
�֔�2]B\<�r�hs�R\���ӫ�IC�.�b�t�5m��~����d5�)�t����@�!�S�L���1]���J��{57���P���Q����[�АW��k,n��3^!��H傽Ԛ|v6���%c��Bo���s�b�OD$!b�q����E�%<�aB�߅�A
��lFnl��빭�K=(Z���2��A���������9����|�r!rtʃl]���ʎT�2%[�+����Mc����ONjvͳ��-B9`;�9V�����h Y|�󞧎��-�k7k/~�f��i}�pt�S(Y8����/�L��k�ϝ{�48oq�e�
��B	�[~��g��R��~��&_S��h�۵oJ	�Zy �m#8�1m{�0hGX`a=N�N���K�4�9^-*1Xhv��c�x�Z�S4�X@*}��EQ�H1j���a�3�����"���E1�0��:8cΜ &T˫�r���y@$�Z��@n����	wd�w}	ʬ�/Og^$��ݖ�e4��A�Z��ʗ��2��f����P]���D�S��?8���y��Bf��s�o�G��\n��P���	�JA��	G15�5ʣן��̛՗���|D��豙�	�I�'
d�ȝ��B�L����;��D�ፗ�f0�H+m����NW"��%�ڎ��JK��|�[��(08�˟}ԑ$'�	[7����7�2H���"ѩ���(�Ԍ����T4��C�Fuݴ�����2��*�'�9��M�G��D�6��6���rRP؋D-�{ �kj�����79Тdy��2��p��!+��k�<"?f��	;�2F�,פ���ʵ��;�\���,��=�tХi��"��� �hM�|؋s��ȩQ��e�PRa9���U!\ ��FI�˾k΀k.w�[>s/�b���p���Q�,5����J��;it�FGwoqŊ��f�N�6�i�������T��,�AuV�N��%&���ͬ���=�dr�@.g�}��=-�vL�PVd�����n1@,�S"��{�m����R�c�lXL�d`�j�=��\L��$��Fϡ����aB�ȍ����#��J�$qc6����g��O��I�ږ�I�l���u=F�I٣K��R0m;S�A7�goś�`��R���D\�''q7 6r��d�$�)�aS�/��dơ� k���Vs�G�!�g��ΤC�5�y8
f8��t���i_�������. ���Q��6�7�X�zw�4��֛`QP���҅	{�S�>&�˾�>M<�U*%�VapY3I��7�yy"~U���)�X^ܸr�l��9���ɑ�z�@Ǯ�r�D5��<�w,V��6�u�LK��O���!Y@�T;Ȣ�\X.ϿS�2����Y=`l ���e��{"�I�&-_�,O�#�e��f^kw^~�tN�b}>ƀ"�x����ט�M3�~�Ք����J��D��kLN�Y���B�A7)�c�����@_� �ݷϷx��)����I1>���Vu��ʕڻ�L�Z1w�գ�J�n|�tKx��L)Y�_��b�yj�C�Ti�TrGş#W3?�&e��[��pF]ǝ���J].�P j�i��]:�1��j�<�&-�y���߉C��#�4�멱��6-IzJ�g+�V���
����o�\����,�ji#���R����bz �S��_A�=5㉷|����9�8���n�G�
�!�2���#��Gg�U�7�F�{m%sUy�éY�]��u��b4����~������}q��s_����g>~Q�>�Ƌ�m�8i�n�l�G����$Y�]����S�Fgy�'�O��خ�� �&�D����|���?�~���g-�����'���w����6ò2U����җ�qi�}�]��T(U�;4_j�2�|4�h�'�M���LJ�1�ݧMtSI�o�t��g8�����ZQ��K���|��tH�O�v�M���O?�����:?�4�WA'�c+ľ�[�W]d(>��!Sb��D+�u���fp�Qk� 8������0$��!���/��'D�SK{1c���\)��������K�]�ʴ�2":{9�]@N���]r5�!�S���fU������I4�1N�ɪJw�:"s�� �,�w;6<����z�pQ�Y�aOX��%�w�D=p��I�z��#�tsG�A�N$GS:���3|���{�/�/�k1�B"�B)�vG8�����B�,�&M#o�݇��z0Ø�'�mz�;���$Y���[ɂ��3a�aj�Wu�*�u7�I����&��CR���	�rH�\M��V� ����)9�jS�(��*%y�M��L�
��.�B􆨑8����H�ΐ�Möh�1\��0?�dQ��R�BB6�M���d�U2?_��]�C������mI�ׇ��@��CWF�AwBQ��X�:T��a\�P�)��CPQk]?צAM���)�BޒY�a0�C'_+�h�-��	���M0��y�B�P��Z�@���#��%$БF"D�_{[���4zw3�$2k\�fK-(�4��6P�X�z.�N�S���"v�ڛsH�m���:�9�wt�ި����"Q��-X�����5��H�P)S��/�TN�&�!�H8��0����!��9-�ШD ђ�+��ƅ��<~�����?��
�mݍ#�іi�߮~#uq���P9�IQ�YJuF�
+��z.m&���Ѭ���� 8����B�U�9"�xv+�����_�4K�����ȭT��^YR2�$��(˅�J%��o��m~�#������tC	r��.;-m:�� 1�"�C���O��!Z���ɂ�)R@��sfb�)�$a?{1H&��I���_l��p�ZXG�o�BE�#��voD�y˷�7"^~:?
4�%�ٓ�
�O��-Z���Ի�A"�i��6���ؘ�u�o8�ֈ����@n�#���9ξ��y��ɚ
T���(��Z�o&��g�Ǽ�;ߧ���{D��" ,j���we)��U_	ؚ�x�zz��Z*Ne>J���+�HL�u��C��$�D]4�����|T
^�	v�.�&�eu&	)�k���)����GK�X��(�����[E�:w��/���"5ISJ��zP�9B=h���UDץ��^�|�2�P+�H�%�uqy�o��<�B�tl�W���nb��e���`���ȓ�j�t'�>nlU����I���Vzu:�^���Ǖ!���\>~)G��7�/p�X8)�;������RdR�k��U1G���-�?�)��S%c@Q��&b�Ǘe��-��Fm�p���r"���n��F�qX[G6�;���R�����a:6�ZP�8�nU�/z|�d#_��2�W�Yҵ����^��A|C.I@��dA6��~�+�!�)Q���϶T�V<w"}�Q��D6�	U��0�r�����APg^7���J]ts��5��S��k��uHG���,]틬��f��cT�}S��\�,nE�Q)�u�3���.��^`rGk��"e�)����R��o����)k.I��%?^� n��A��w9[�lq��@,A�#�e�ڈY�4r�}z�Ω�D{�m=�'ރwq�2�>w�¶���2
s'�PWo�\�/���ډ�^�^��<`fSs� J��t�D���c��B*
{P'��<T"6���a�	�~���E!]K�����<�hz���KH��'����L_Dqq)z�%�N� u(���V�+Ş�kK��6�m���?��\�z�)�j.kp���UmjfY�]�;�쇰|`D�tk�6�/�Ӯ�������h�e0]�:핑�scJ�PRGm&Ѭ|��NI-|6��d 4?��``���W��8��K�m �=�C)�`�s�xج�/zʜfD�Ŭ�D�oK��*��_��a鴣�?K����D[&�{��&9�k#�i�j0�.��C�̽�w�>�Aо]N%���n��G��|C���S�Ηg���2co�u�QP�Z�;�ʷ<9.C=m�ۃ� �DC��Fi���}�P+�%��M�@J#=����bh��J#���7p��p�*:&�ɦ[��䭃��Ҟ�o�$(c�,/�R�_�"����rS0��R�{`� ��q;��2�9�,*\u��k6��U�{�V Fe�ܼ�e�����j�EY\&�޼Qk/�:�u',�ۂ]6�R�,v�Cj��!��X�=D������ha���0!�*I�i�a[�F�_�0E:H$�7"b�rq�!�9�bT��δm���jd����&r�׬в_BݾYZi�Z�Z����8��vv�g�q}�1�Mύ_����t����|(��9W�V̫ye:�|��tmc�kt���"</���`8�)�!�a�S�8a�0��w+h3)=��o��'��O���b$|�[������䆞'�}3'ᑡ!����_δ3�$�2���K ��lǔ�n�E���8�oJG����_�8�����0�+�F���gw��Ŗ�u�f��8��7#�/>��[��lU��xF�3�Y���o�6h��I����^�Wɠ�%y�|#�?v��WJ������Tr�w~р�m&�җ�����C�O��Ǔ����&��4����ɋ�B�2���7@���!�]{,.�1)��,�[cEaQ5���y�V��ށ;����1]�nǚ�a�Fȸ��e��AC0U�]��B� 7�)�P�|��18�`���&�&����̍X���(�_g� �R���x �� +��1�O�̇V�-�5�~���� �>Yqbq�!� �xJ%����§�q�P2˵F������J�+@��Aܟ�S]2����5�<�5ק�AX�bpd��%�uj��i����`��Ib��w�e�������(��s8�C���tM� h�%j�r���1���8��
G��������H�k�*�wN�gr�5�n9��N[�+��x:L��{�
���F6��d7�����-G��>	�-0##'0����;,W�̯z�7�T�]��qt���^'#��"2����v��c+I��}6%�Ǘ�͎�>�H��[s���q�g�������;}�<�
���O���G�U'A�_i�_�ա��v�@���X�!3�Z�p
������� �;��Y%�w���7ެ*�e����#4��\�k�ć���X���[��ɮ���h�T��rɑ��P�)�{R���:�ȯ�q6�`3�F[�a8�&efO���=m���m�kʢ�OAt�a�b�8���w�"J)��1��b%�w~��h����Z��F1я�-�5q��f��&��c��6n�v��w��R��*���ypqɆd�Ow�
+�j10���J��F�a_�8��_/�l��Oz1%]B1����2��Fg��K觛�J+�
�?g���9�֍@��u�;{?��B�m��C2�����V�Pd�'k�����-�6��j����j� �e8E�Wa���BF'�7��J�3~�G5r�#ʀQ[xr�H�	v��/v�S���QUv�7��|y�����O&?;+�ؓTi�@Z�$���"��달�E�̷� @�v (��ARL��?]��z�$}E%�y΅&��V��/t���F_�-�87��g��(�K0B##l���:K�m�H��k���3TI�O8[^��Z�t4E��;�����F�4��}��+~���㥙�玛��ԩyZ�.�����1db�|gw���{�y��y��L���f�qZ{j�K<�B��)��_�7�F|����PF�tr��=VC�k�V�Nf�g�U�[��𮗲=g���eVF��},�,d����J�Ex��ѥ>�sF�#�E<�(|�p�mV��&�H����WV�rN� t�O�V����Pu��|t�#_+1��}U���d���>���%�|-�Q�t[@%�=����I�x�c���-�Q-0�	AN-_�4t�-�t�hw���X����wzT�^��$r`�exl��4}h�|�B}"5E�ƻP�d8��$r�b�3.mm�c*4��e*�)��B	�G�؄'�qD@QZ��>-��,�V>�i(��3<A>�0��,M�~N�!�����0�Rh�	\.E�&�Ʊ>o/�)�)"�n�K�`|-�z�ҨÖ�qrfvүI�3����~(�Q�v*��.)&cc
���9���4ކ���b��	[��!H�=�x^������$�}�ͩ]��#�R��.?|��ۏ/p'�hϕ�x�m��#�+�!���8���T=�3fKWN44�JzMs��b�����5�P��q���mv������>ݖ�֡��d_�z�&����qs;/�qߌ�8�}�NC��\l4ӭ�F�1�@y��%��1�5c� ��͑Y��2��-H��f���� ��w+ê�{��O�K���� &JL�Os�s�f�H��u=���"���km�I5�c���2S ��C����Ȉxᩨ��R�7P���9:暣��͜,��X��W<b���F@�Dk"���)0
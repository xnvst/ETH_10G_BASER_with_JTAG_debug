��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡j��-��l� �3Wʴ ��ȟs�/�\�Kڰ��n��T%�s�^�Xu>���Ş\tֆ6��¬�⩼m=�[��P���'�x r�Ա�����C&Oʱ}�"�_xsVh��k'�׀�gZ�	HB^g1��M�.�/�#"y��	k�v�/�R�-���(p8LD�މ=�@�tuP���aC�kX)[?3�9�J�Wȍ�n�{j�xU�2��=)e/@nҋ����QMt�� 9����������ͽS�1�
��,L�G�$��>T�4���)=�� I�W�w&G�u-��CMv�R��9�w�!	'�3��غ���v�2�]������Wu*5AT�z�y��	��(Ԥ%�Y}���	؄��
�����2�H� x|bq�~y2haYћ�H�x�q����^24���%)oo�m,�c����T��/��-�a �����Jj�P��}i�?/�&�z�2����#h�O�X��.����a�&�C%Ԟ��#茶�Շ�q����"�#�!hc�#4���]�-�Typ��h�)� \_�a��X1ع4��H7FuՃh
ro�x1�<���""���WV"D����^���y�YP1�Ѣ�šԎ��E���GgX甆e����tz��W�pߌHw"ť���CJ�Ӵ!����Ԕ䔓�0�/��>m�~<l����> �,,�gV�Bm�%�4<�֕��@q��8�l�Tw �1�OV�2ƚ�2�u��i�_{mf�qI식%���q�;�{�4�d����vb�DCC��@�cK3J�O�WD��#����B�apgl�s�N��g�����AsR���p�	���QsuA�i^2��k0Iη�/�4�,e��u��k����>:�8l�-)�.G!r���E�L��M��2�wn�һ,S@"@7�{��j&������o͟j�0D��,´�A�C�1�Ц��f:,G�2r�y�z3ɗ٤d��w�2��-Ɲ�4մ�RT����+�
�����{���	ץ����!,o�a��\*z�R4��g�uz �.�ù�L�7
u�.�P V n?X�ݪ.�\6�$$�:o��8��MV�����drw�3��۲Ɨ��$!� ��!~�<
K��NhjM���mݗ�Θ9{�ŻHQr�gَ��8��˒�-�쌭���	��e�,Y ��[v�1��kgȋ.0;Ekܕ/58�`�`�P�)F�v�(˘ɥ�1�"�(*��v
�^�N~�<�	K�Jk�℗�3ҙ�0��Bf�J3=�{���>����
�B5���K�C���"�@&簊5U2��F�l�e��=�[��I���C��qo�x�t&��pT�G��8f�W�=sTޛd+��y�q���E�چ��H�O��~��D�g����9y�����EQn3\�����y�h���d��ؠKw��CQ�B���Iư�覬��SW#@�g�@�F~���K#�*׵�D	����-��*e��tK�:�(I*�"	�:��A������F6�8ϯ��q���!�u'��9�n�ޟ�}029���I>��b[ U�Il��=k�1�q��FeHǦ�#�(0W�i��B0������}M��VS�(Ԏ���o�-E���F��q O7�����j�D�k����1��!���DO��pū̢ܲ"<�ɼW�>��������Z��`g�A@=�$x��
o58Ü���S�����!uje;F(OSa�F���!���a��-�AF<�H���Իt��!P��*��;����kE��E��WvcWP���b�!*�dF�g2,N�v�����A{�� �l�����W�í��tW-���t�NiN��3k�\@�m�l���˾̊]�l}�%�nd�v��%l��s���������K�.�[��e�*���Rr�k]��q,kv:x�o]5���ޢA�/R�ſ�U]P31�8��nR��.1k���4�?���uo�`�6!��6=�D7���~� ��ݏ�)�P���x?��G|��t�u��3�Z������̮Y�ni�b�r ��F��E�CZ�WCܨwŖjƂ>��S�ǆ��`���iE��"��n�I�&`N�Y\�觜���`>�&���3�}�f�(�Cjm箶u�=��gF�E�O\�(��t�����L��?���L�膇�����l��Z�>p�jWmF@zsV��M�(AT��l�P���ױ��A��O�N<fY�
0"����1|$:4�*AE#jo��]�P�%�2�9��}��2���PW��,]S7!>{�nōY�m?Y\g8a	���JĜwj#3�I�Yi�t��h�b�wx���9�㍸ �/�o��Xj�V�Sy�,k��]���M'�G [��2����p?�"ҨI��z:p�U��9Ka�rܦ]5� �6Î��^JZ��d4���o�����|�]�5�K���h���sƲ~�e?�|���`��L�{���YMs
lٚH�p�i��p:�Z��&-Hg&u����Wד>'������Z���T�S��͟��8���.�q?D�
��u"ug*0~�ҍ�y����K�
ح!țv���L�h�1K�"ĔU��2���Ŏc"h2�J��.��dD,��։o�5�����4���!Iszz�%b���|�|�����؁�&�X�a�l�����&���b�������I߹^���r<D[<����o�0���ͧ�8��g�����5��u���3��I{��}5Dh$t��҆�g#�S�~�"�Q nL���\�qR�m���ZIϷǌ������0�	@����~�4���[��n�O�1��Y��^��b��,q)�����XxL:{��:B�7 |x�<��/��,�B���I���"C�M�	����L*�h{��������S:����P�f�l1�I����D�{���!���(���:^��8�����a��'���5*��r�#��\�.0NF!�Rt"E��g���x3����N&�mj�K�����F�wZ��7FH)� ϶(��G�j3|1�$?�'���ξf WE�-����89�-�f&�)�+��fƈ�B{pB3��;�1�ot��u�ebH/��Q�˨[��Tn\'b-�\���0����1<z�\�z�|��P��ؚ��z!%u��_}�8+<p�:];��\��q�J<�G>�HΧP��Q�\���#9�|���}�E�_����ZU$���M2z�T ok9� q��}(>i@�e˴���$I��m��/�q�!ؤ]L�hJ��5��$"�� �æ���Rt�9�E�3�1��3!�~��d6v9F�|t��	V�.����Y�^Z̖=ʹ��As|6��kPjQ�"#�e!@߭c�vӰd��ࣾL Z�n&���D0/`;�C�nX0�ٝyc�;�ɱ8؋��ܽ<_�Lh��TW��{�6R�p�
:"� �R��2ǔ#� LJ�g/�5G���W�&M�)YЛ���H_�䱿7J;#66w����l	�� O-�0�YVg��&)��؄5��Z+�j�C�����̿V�K�o�ٲy�LO�U�^3���h5���a,���dә��W��J�B껪�\��n��u�lD�ļ)��.[���J
]ɂ�L�ݔ�﷚o�2`�bG�u!���h;�d��*��Y�]�W��.~���6��ѻ�����t9��}U�]m��gN��!�h<h����!,h����G_�����I6��l�h�)��9|q.~�Y?�ܥ{��������*@� �\�5�y�ܩ�à�!�[�ԍ�
��MFkFmH)=�b�+��0pEe͞H][�(�t��Y�b%��7�*CY�E�����H����X ״a�;Z4r:}&Z��r-�*%�We�6�8���dĆ��řc*�햱޼�+��U��y��v����Q�yƃT�h�n���l��[=aP��*�,M
x5�iƨ%����8q-e��#bƸ��]�S,S�n�>)_�q�p����n�
Yye֤,;��C[Ӆ�u���J���$2}�Dt���)s�3���{��@���<g�EYks�^+�_�;������vp���$�,�\�JSt��Z����I��3�Qt�޸��>�O0{H0*�*Xj<W�1���Ĭ�A�l����d�8��B���_�GS�2��+���9�fq�dw�S�}�Ҕ��Z���7���>� ��V��W�[�J޵�V�M#�@`T|��~��F�	@��i}3]O��b�C{� "M[�?F��q0搣��F�KI,"�t�<��a>�.��s���'�����-���S���J�\*��F�ْ���V�X`Y��s�p��3��Ѓr�/��2�h�Y�C�mV������=�����!Q�^�	��f|�^��ۏ���;<�r$L�g?<��ܸ��ԡ/�C�����(�O�Ai���!K��}��uCVI�e���ɞ��-H�9�I.�C�v���􃑬3�$ ������a*�1�3�
?Vڹo���]�%_T(u]�K�#�����J|`g�E��7�V���'��VuQ�=��=��D��,�b�����Vlڬ�#���:��LjO���=�_��Fd�ä�����[DC�W��X���Nw����©h�[��k+���|�X3���Ja�>k�|S��.�����N����{�s/x�k�(I=�@�#��J@�|%���!<����6g��k�)=��K���l�L�� ���\����XZu��iZ�&\9 Y��i����fJr�������d�;�X�e%`�7ːSd�&�h;[�Ry����տo��#��(�t�s��Zn�p�Wb�m����V.]$N�"�ؓ�U$�?�̓6���J��iH
ݱ?���kLp�#!��V��a޶w*̙:��x�������%�eZ5��dB�]�𺵐Ӝ+�.2Y�#�*E���櫮�~{>�#b-oV�����^�Y\1$������W񒓟HC�@.�pm݆��"i�݋� �! �_؍R��I2Ϫ$��O(�����)_�a�vRu͠�,h�w��;Oj�B�_j��	"��gN��I�c���V��`[���Lm%N�(X4����B_�.{=�c�'\Z�Ʀ�HD��(&`:�$rm�8����t����l�Y&z(�������m�*ޱ�;nL;��M��~��,���a��3�*6U�(�w8�F���袢�Y@��6�:d}a3��6�߈�N��e�T.}�Z�gξ\b���H͋ί�__���4e{�nn�:{=�{��ߡH��GS��fp��j���2L�����:;�Vk���i{Z�u��sL%s�(�(4�^n�_!(Mݝ�ص�B�����g�ko�\<D�ՃJ�B�@�W9�=r]V󱥋�@J��	c��~�%$���6�$���\ʎ��b�?ܖ���e���#d�<��Cyv-D��mx�F���fݳ "(g��[�����݅s�
,�Edu�rM:��X�ҥw�Hc����ͻx��i|�?*����=������w� ���s�l��Z���k>�p�9ϭ�!���	Cch��(Wu͂�ze��� z</3� I��"��`��Ae��0$���l�_�s�����g�;R�*v>�^`�:����H�zz��^��k[��q,(�V,��ԏH8��hAg)���)�����J��v3*�gMP�,[���"9u̢�ǈظ���)8����v=�*�q�8�����^Աh����v@ٽ3��&��S�p�	�i���3��b�v�m��HyEN�p�ZKy�<?�d�,0�N�{�3�#1r��w�j�(��%��0���)�ӣ��/l���'��N�������7���?���� ���a�������<��!�����n��c1��� te�0�[��l��f@��W�>�|�[��H�[\�Uz���qo8��~h3�D��^�I��|y�+˲X����A��†���/_6:(5T��J���.�K���IW�x�D̀�T���w>?�4��V1))�j{�[���r���������.�A�::�� �A�Д����@z{'�PѸS��]x:�(��3���1t�˦��{�x!
Vt��2���x?�aI:��M���Ǧ���9w��U�o��y ҵ�d|~8���������a,�?��ab� l0����)�B`H��\B�.��L���y[�.�Ad�	q8}]�S�ym��]\��6�;�Zոmo��ﶴ�0���2A'l����>�{���q\�����+�[S�LB�xQ�h�$tgnɘ��;�S����l�<'^����fAz���n�04�;�sv9�v�+��H۷r����5���Y���~�p����N��̲�Lk�����H���6�CҸtq��nd�>�!b��]��5>��X���=�d���}d���M��8�T&)IY����h���Qۿ�1E� tr@_h̐�rh�%���)��qii����#�ɏ��fד��g%*�N9F?ԛ�d�r��]'*�i��\H'������g�tak��.��#�L޵i�Xo���|]��=����KCc#b�ŝX�6� 1�)��Ή����d���k�b�t��d7����a���%X�D�E�=+Z�Z���xGUH��>O��O���N|s�8ЄÛ+���~nn7 �-^6Z���~sT1A+��#��p��\Daԯ뾶7��!��+]vE7��%�Y�%MU��L�/�):T�$!�Bg���]�v�T��k�`*�a�b^~��"b��dK�7o��8)>"qRH-�ٚ�\��Hqu�P�������=K�t���d��"BT=�UJj�G�u�ne�hCg�qΩd�\�&���=��ɔ��A������90�V�f����L�B]�����?�P�΀0�$��Ŗ��	�Kv`��HD;��3���G�M��X��^�y����e�}�xFW"T$C�PJkk�{�-KD�r!��-�h�G��9 x̸�w����f��D�����ݛ���19��f-	t�����E,����� �<��ΞQ��(�$���;����q��ؾڴ�Uo�jr�v8(_��gE��G��l��H����C�
_���|����S'0ٻ�&�At�WU��� *�ë��M����.[_t��I�:�>��%�9��!�/vI�Z���[�Ȇ.h*��ّ�	���0���ɤ:w�؁�N���r�Y-�;�_H�Z^X��4��mY��9m���,���xf���o������R����f��l#�섹�
�+ ��S{��c��`X+Ff_ؔ���(��c+���|�H}�\�ń��ٜ���3c���;����S-��:|��QIj��v���u�z𯕨G!^8���G-�^d�^�� ���鑨�)jt�c(���f�aQ�xǄ�k�J݁"<�2NF���1!6��K�'�|����!���:LЮj~�&e�����h��������}���l9ޜy�$�(�p��8�'�gO
// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:33 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Uzuy4rLy82H0WBn/aCWZ/CQHjnO7fAhjmB4QtpOaj2Nw9406Uw/yFZIF2dSq3LAs
JLrEg9CQWuO5U6zr8oxUI3Q6aHLfbJsLCFngq8w5Gqvc5b3ySSlXb/n4mNtT1A2a
nnQoqwtgux+r5MvfJw/GhZJMGV8ouK3xf9pC2DzZOqc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13472)
JJxAPZlOFZgn0j6Qless+3F1Xz74P7owkGuJktoe0Zc2ZYWga/Fv0msCmwtMLhVQ
4Vykt7Fa8jHElXGHtXq4kQfxNYGdpywj52qA6L18IaD8xybA8TsSwhRUO5PiCXgj
6iODu/d2gLDaAF5uETPe4E7hGv/DZ5Cd1Pf+vK2XnJOqI1/gpCwARJqmVJb2xSXi
33xlTqy0s5GCwzpwQFgs778+Qzi2uR/wTsPakMKSDep+4QYiOi6/goRjwT3LJvEc
J2wGmmqu/1YpVyeGtBairMcOa+I4DTGeuvN90ksrMPkIvHfARzToMqxPs+Swp6z/
v+urDdcRH6Y0t98KWm61tRdqFYwDkLe3IfIRINlokj0BOm2RVYlOqqneOU2hm7m/
SnhQOF6uLlF8qB7gb+l1sz1x4kzoihKpjq6ZziuPP+J/Ifs4h3VVxVfpOsGF7f/y
bEJr6xt4fexKt8f8c0Tamus8GwT1viQK1WqJ6hnrWh1NijnoqTCHFraX9LF2BJl6
LVT8x2pZw51S9g0KHHjEx6zh8D4rA33NRmpXaQIOJ7jMpCoFu7god36xfqXH1SpD
H3KxbQtLVnrUvxMvChr3Hiscr+BJIqIWyiOLDYhsrvi4fZNvZO6CO0iM9M9L+M5Q
74v0UlCCIC4NS3qmbrPdRRN1tYsGNzi1xsLzpdctKpOsMvp6rJ0hc5UnxWJZnnMs
gpnXKDywSbqEh2SlQ1EZGZexOki+q8pJe+fQOA0ADz5GRT1/cz7FSneEkjaHt89J
SqYLMsZFWQyitb6rDl3hvDOUnJHN0Q7WLMDtSjkvRMFZW+tc9P4kE0v2vU+YRKVq
m4vlJgJvImfNYnUUC+HBwjARuGeJ7YWK9f0m1fkK7d2jeiS4I2Ary3x+0ebzx9Zs
PhH/i4nXXUMwHCHO2QwyVOxTi/d4lYgRq5ArAEIaOSkcYKE9JeK3QFIoeSk3M5QA
9G5Kb4e0w94vjiR2onFQGb0MMenkxlRXyWOCjL91HvzW3w4JDEy01hyJebqLfMeA
3cK7V+1OY8+d+TyQsZB3peOE8x2Vetl8487t85XSwFfTXLflAIr+Mj6Lf6FaXK3a
G3nkibDE4axEV83kN5fRjNGz3iC1K07lag5oTtVB9x042sV7DgAXxKL5s4t+CGVR
G3f5LxC4WeNw6toGaFgApy3J6rzc0HXtcXWdl1Q+0jnPUYyL4JZuFr9CCSXbjzgy
aK6e1hylAzQJM1tZsrL0vzbu0WNhxtQCze+BgYj4dTIMJKCpU9mewUvgF3vus18N
XTLuvkA8MZAJvPx9KuX8aOlVRF533Lh9CWYZB1fyTwNbTa6eZtynx11hrqNl9Rd0
qMnZplsdjxjFyG0yNjmYK4d3+ndo19IBbMfz5GyM3QwbGCTem26mR6+K7st7O8Mw
fDnSmoBEoCUTtcvevzP+oS4DiB6GRzOTZgQ/ao0CEaRjel3wkteUQbS2zzPP3M6E
XFNHlBFNwytV5/d4RQfjzGa3vDy/mDyU1olw9Gh5so4SztWRAmlTbOlZKacFe3vY
Xx2MDTDKKDXo1Yt3adhgISchI9ZeO1YjNA0eRYyTL1beY4omjd0TF2X4Rw5oQYfN
bhMVp8eCS4+M1Bn0PRXKYFc5lpxZi8G1hcKrE9fzWI6q4xFI/CO3RNpncCznVJVH
LcUMVwpYRdk2Bt0qKNeDqdbX+Pdx3O8YWeHBsMXEG2RpATqgY3l4Z8QeYq4ppS3Z
C0m+V2QIuOH9eyIYjYuZNlmWFPFKjt4DKXaBDfpbVRtCbqlJYQ+xi/RsAOgL0crw
VbqWurnNo++Mr1h2cMvMejozyrHKXyvr8aMLJq3e0JshzBRQ8LAz4Bazo8RIXgyd
2wi01p5eykGWWumLJFN3zG/k0OtQAzsFe32XEhHrbncwvrJGOPMGn5IxWbZUg+0j
I5H25rkTMOWuWypQvHtZfqBzUN1jvOrmLpUX5yItfeCqWd0xZGEI8N7w8YonPMKy
CztxSXxNGhjV2sF+dE4IqbqGRLW0q0EmOy/CH9Idh8flTcMWv6dnS5dsYpiMj7So
HLesZVLhVjgg3q58NXQPI8Ec23Do1Ukd4MADfNDUb4y32x67avcKEzg33OkWXgu3
M1BDpB6GmrLsX3J3yA4ILEbSPSuEjkJMmI/VBG1Ae/PwIertPIbX5IA1+tFJrEgg
qyeujVwPZFlP3hWR1eDTW22z2OvRXU6gbtIDQXm4N96Xdc4nrihZRI2pn8DDmGUF
+5ihS8HaKP15swE2i3F3QrN+zWZydwwddEUcO/RZDeG1PbY+nCxp1D+8aYVbMQK/
B438PdIfU/nKzA5lhrk2uiM8WOOEz9E0QuenQ5kdpOtl1yl9F0Ke/BZhDXocEmsy
86MmA3ibJPr6MU464SYxIC8dJHggFqugZOhZBDxS8NgYx2dsUWX9EbXe6MEinkmJ
ZXULr6HI2uz6fdN4SyUDpqajDeFBPmiFWBcp8Q0jNUkvuN6pxGtIeZxlKpIFZQPu
Rad6T6QNWZIwr6AksQi972YclRyL5pF59IXigy/FTbkx/h37gxM0mADhe8y3RZSR
uyvE1whyDBXCVWtgREE2qB5r/YiMTAt1d5WDYv1dhWspihINELFq6tm9U9s8D4ce
zL+bnrqZvxf4OvQCxxwjDlOydtBJaoC6xwUzpdbuuvYcnvf1cIwKUeTnTYbIJTnA
vXWxKqtZcB7bW64SSk8W5Bjo75ZcpVabLedm1fJ3OFAUzAFAXmrDqd7iLzbQIdW7
XrIFrB1EIMi3raChZF8/FrOJ0aV1/Ka/OAFR4GTxMk65t4RkQzwPEXRAuVnExdG5
P7EP1wErrHDIJBOT42hiEBf/Y+GlTOfIr5Y0O9AKV1X3M7h/6NJ7QTi9RLNTMVbI
8De0/EOA2LyFqJJMFizaCVE7ifIaIPa7lcifONXMGTf1WHlbtjZP2BdBHozNhJM8
kNUszKgE1w/+EfzPu1ScvKkCf3cZD2HIy8OecHv5g3bp4z5e44E7ceUQf7zVmRqb
dn4pbfDH+LfrP7ho0OT4sTbNbHDAZL8pb+k3J2qqtlRSC9VWXGltiJaKUAcQ6Ob8
IjSbkODN3/YDQ0YdfcNTXJeKE16ViXtRiqO3aEPgU3IXyrohjt06EDhKaN1RfAVP
NBSGl02EPo5o80Y3BoMcwMpj9KynxFqjhhoyvbT4jOMJZCJy9OrcW2/l0jdvTs9G
Xn9kfI1uUZxH96+1j6brq0Lsx1xZpgdUDiESBkuCX2USCh0PyVNFq5jTvA5dB63q
kzGvC7mExqJBoNczYwcrYo7CdguLzbC+HUSbFwHZ/aOVU1KF9f/uu/geaLd2Jf5I
Xu600uOojCcEVGaeecRzPJzcCCXDnnoaTCLt7hfvOgIqmwZTrpbHUwI/UxzntoW0
aQTMgEr0EgvlN3P9G8TmeaRHMJqS6jp5vJZ+wlWp0hpsGRjuutD2R/Xegs/L2tzp
02Z6mcMhO0UIlOllyK0u1wPoeDZ/MSTsKQUd0w5IVq1Bkc1012UX7tnEkxlMf0d0
i8uR8vqxGb1jFAQqS6QIBGLM1Qkl9Qj5gF3TxS2N/pp5OJprwq5j1pz5o2DmFMNS
sVKSwFI8N3lY0ldaRvXIdumZisx7TOPCMU8YJ3K2Cpdl00TaeT+ZMqXFVpfUGxwy
8k0ljdZyuPIy41F9JwE/Rm7QXvRVKa08YgQ/uCE/W4mG+Wizu6tULjXjD3zZ8Qta
9d/RYoDwCmC+/it7G58LnDHwvvsGiJY0cTC0oB6um8O3FrKfwE9M35TMSFMLTGRU
d05zSWzA27wFrWjnzWJqyyvIHiBxwsiFOhsCgbybOZeg9nNtQwYb/3CfRe7RvRkV
4KcbrVyhQKWWQxvGKLjVRaJbrO6amVb1l9qflhZZcrmV4xaWwIWzz97QSIqLQIOG
FiwGUoaErQPLZUW0YNNxUyolQA8Hbno0MTy6kFfgy9BEZRh1kMv70+GzuyHydQuK
apxBpnFAZX+lMWid/+KUvyExc7qVwfFclj3kf9ZKf/EaOMAkZDSevDvPqWRwukCz
Drn2Smhj+DX2Ikg96Xnz7u7//oOLA4MfKIFN0WGSeEickS2tutDT/UomUSYx05tr
/Vsxqxp5BSPqN7735MUP2evSRvkaJW0u2G67KbIrCV9eaGMs1+F5DqpG3MWM4DZ6
ycbyk5e1ObgHUdc8roMVkj2rRa84zypGGTxKL0kVjB84FgvGlNcXg7LdvJmi4K0T
mXotnb8One9hn9Qz4+sdbd1rMh4Gsrx9t8VisgpTvnY32yVm5GkzwgPOgACsn0gf
R2HF4yLOfqqRVYx5YDGtzjJjhV/V/aZDqdaRJs2wOCWNt4FHfCqGkg5hn6kvVHIB
DHiM/d366cLXaMJAceTYA8RnvupuvQpq808pTx5Tm86FqCBl+oSLKM7dDMyXZjim
8JdyFinblQTmwasAKxkAH3Hv0b5cfLzBVc2DGrkJf2awAlY7FybdFqUqIBNKXYor
yZQREPOyEYj/qvNodu7I/lOPFtmqqT+9grC+gjiO4sRnsOCbFEcvqbT9IYju4ZnL
5B0wCOj9AvatJTJ4FrXkxRhxi1qGl5WiroHB7Ll/weF5jycPi2woA4Dqzcf1oQil
WDfO5XgSRvoH/5xd72u5ZnubQEUOZqjOzXU/LmTVdmDaPl6ReCbL4kzSwU/kIYk8
eL4oLyclCodINSjv+dzDcT2dd+t3A6XvNK/OvdzBHiE/XVV6q9kiico8itJe7MJ4
FwMq3V5w4P0SbRcx1QUTVjxUyVFUsYqghchNtAzyMHxTU9+Nc8mE5+YizhF0vXf1
c3+21FbiJ9KrjqO+McOku7ZpmufSRSRjqLKSC92Oc71KB+5XhCInuDlfFCyYeNso
XXRSUl13biLgjIIRuBJJd/Lx0lv938l18ClaRMlhsW2TSK9bEXTuo9aWraK3MaoP
DQlVTMy18BRQeXdZIkil+EMEHd9xy1OIC/VfCm8XEwb0lHBNA/Ne41R9qKVYmgR3
hxkqqIn/wBFMaTJzqwUe/81hdNXzQsSQ10XvAEZv0TMRRQDKMVammXqcNdx0kXjL
9caH4RWFDXhjQABkpxQtKuP1d3gbidEcuBDwTnAmCyRt9hqUlGlufQjeHQo0WKPq
WXVRTBPNViS/preL83KKO4q0lJl7Bun2qNRpfHPkhz1glulkmZ8NIRvg2Ebd87Z5
11Tkaw1TpkeOdil9WnILQDxmZAmcp5Q1QJ8JWnzSHUmigUyPTf7QnUd1xBNTLsgH
rI5LXAph5luM+KkLnRds44ksr2XlPAsBxx7AxZbkXAQUAu9yfs9TblOi1f8bSmjG
MZsGURJ+Y7qO2xw2QEKMXv8CFBZQVKu84glDwdwOb/V0JpyIQx9KpCXIII78T9Gm
BSPMElwz1SD8N1FRXyaSWrCGx9CRO9hZAjOglJQiO9d1R1Xr6EKUubDfJKFCEGd8
WiJ1FVlPnESQfAXwRvCGhNcNRsx9B2sSwkYtPrCECNrPA1gOKX8DZv+/gzHzHNLk
6dJ7pQFvUWtRjaIdbkLzDYnZ4cRmeEgCqoJ/Dl+Y8dc15v6LTzRQfXBZyqXNqXBV
sktS956r4sHW2SZiZnHsp+pg3Q+PpgL9nrca3XEhUUWmv+n8j6anJNgo/HOj+J67
qIIpts8PmI02coCI1//RxVARGc7dt2RCjKwhpm+sKvF/t7Tilujpv7B3bwF28Uwe
h5eh1eDW7Q8WvgXvMrlB4FkzBlIteBKBdojE5G6Aio/yoj/tNm9pHGhuhulhKFft
2A85wZ/hsh2BHILqslGKH134j91ZwXVnW+J/UnRpkB1iD1E8T+8jO7cdtWoEm0qt
EYn4Mu9uBvnnbnNMl3Fvlmo37Q39HDMNx+sUZWK4js58fTHxB2KWpDPQLsE2WzP4
uwkPONFOSx7IOWZX5HD3AbytbzAjv0wmjktVnNYxUrS5xJwuS4RNqLD8Jdsfj1Xb
8vXbgilH+3PxxONMpOe+SzbVuJaT7lPnEKTMwS0ZFHAImd0MMAIlgccqozhn2LPb
U1+vhoiYE5F+mwl8yShnBnTOlvorMMUcNtwdbbIBbhRtgflJq58TmEGYhAYqdiYM
h0yTrxAxzdE4vNpVQDXqjyV60q0Z28Vsm/GIsE4kNiTtkExxDJylkrrfoi3OHGdB
3K2Wb+BCXuJCFFBGTCry/yoHzBK2QMzWr7tiCdledsum4ewr8zCGe5ys0tUnDUxo
IpXpA+g7HE8Dpb1l2wmb0dUdirISXOsEALHf0tX7NHl4PhGJBplq0CwZ7AtooZ9m
WeiUD2xLUjVKaZWWo8jqc3oDjz3tNXfWIsb4FYdgqV7TEKSEXP6zEY3vJpQO/4b6
6ztqKlGaIrAYEbrJp1dQtTdQaqYpRq3W0aSwKDQlx+f58fwiTY6PNG8/NPj6BpSz
yicR6ZuaIP6fu5COx+immWSq0OFLSyKxDP50qW8Fupq0SAcXx5+euV80BT24yAZd
L+C+i8ZmPjw9KMKQpd7jKxm0+G0FREyEvXtx99xRMPxgwUXSP/kUwRmgJsvayTzY
rEtL8noIQJgL2LKDYGdoMR601nYdKJ/MlnrgCAEh3QP0BjNyb8FG6C3cbsUgyadb
/jzbXbR+fVVMzy/9fSkYSg8jZUBxmx8nmDKv8MEAvmIRRdNwY1Q8q9sprd/wXKT5
EBPF/xVQb2/Eu646naRpPEvBEeBAROjOr+KPm/f2zoEvv8VmLxt9aF4D2giT2FbG
7L2ylhNofL/mEdu1pBgq51kCjycmWEKUAkUNxhYYDO+gW4GGeSWNHtkPacLkcmhG
qRlVHJFL/hHlLeA1Rlzl9/Urk2YnYB55vcZAX+Wqjr1Lk5iLV7cirDl2BG0o+9lS
7HF4mpMgdH2uywJ85NHxnWODYsO9p8+Ati8Vo4Zl0Slrh5snCoAq/DEyGab3WvVO
vM8nLg0D19N+z8zKUPEWTynlJPUfExPN8Xl9kjtjxCnRt4MXB/FFmW7q2VRWpV5b
DyaoJld+PtDN3e9WVlg4QBdXyWiRUtohZn49RGjjCuKv93a9pxbDS2l/tajLjb9d
hUZNupnqf6+gJcULY1fBocgEmYT4eATQJBvAHsT2sUSWbFnJSwikKLBeKPob69AK
WyV7h906JTU21UbKRBQXsI3DbDF3a5svOHEDWHhIC1DYwC36esDeIOPvPylnLMER
AoLdh9u3vbJ6c+z552N/bOvRykJmMj+IjtSljhhn0EQxxTLbj5+db2ayFrcur6S0
+c7A4s5e80gykceAozWuOirAFGK/zQTYeof+M74o4YYqkaUrv94WXh9gxn3NLT8X
myt1JSi3OFJ9mb0PKyZn+PTRdmNicSvCRE0Cmm+XciUaLrx35dn/wnkTCMsg+gez
RkUqMcXKvzy1zgK10hst058jWvI6d27rlgKJ03rC1EPYrdbsAbJpa80Fts3E/JaG
rrCh8q8hcZ4+GWGPHIw0tnZnFURnzyimbu/qGE9501xlnQ1wtXW+6ZAVuKxRsqIr
27Ev9LekqM28EIOL9qWyNvQRfIpUpaYeV3s2TP9Ap9R+xyBUqesphYX024KnEgdz
utAdP1q6QDJ8AS0FIQgsXfZfiA1ut+UseUcvXFzsDjlb9TUnQ9RuPygWFZO5LtyD
jpWSg4FruhMxThui5gHaObhiT8l3AFvACXSWpz7npiCisqOeraEO0pL1Ek/SfC87
TK7tDtUEfxndrf0fwYVE5TqDYDOVWeGmEA2uNgTAWkX/17ZCT6UEU8fMTZFNIjLS
NoEpXtzYspI4axu3FtLZ36aISOWTarebix4ad4CFgPJKuQ1yMiiwh56pvYZEs0hI
60owZxTj9N8YQyGq+fM/wQz2xED8d00LDSUk+zBTHtPB3qPfUWUl39+YYz7yzTfd
V33Qzkmep7Wo6f9JOYP2MUdy/k9O5sQItMWAwI9FlQkGA/UwN9FwsdqQlLJSP97U
eJNz+PxW9+h98nxMa6rQStRreOcHeY3+bgJH8zK6aysV48VELAx+5p8hyFuFE2HH
Sg80DyyC/Z4Ez6nL6B6XHqwj4OIpO9sF55eajzOCPMMMEeJctqEGBFi5T5GQx0mt
WseC9/9TQcipt7Ux3xOLGNIsBsVV7dfmCgSqpaGLiOgCCzUxLg1gP5BqZ2uc09A2
WPWmsbztZDQb8Hr11/8kUVtJO9NZAR2ffQUC2aeld50RHIVPPFTRFA5wGkjKHLdl
+L87IN1PBFq9AD97PR3k5Siq1rGnIO5oc71me+8quDRq6swJGFQiRhWAVm1CJpof
9xdqMg9t6RG5nBYkB6CHiARmeFhECj8w8HRYFbnTPMQ5igzjwSdvvIhh/l6OjY1L
uSO8OBbj7/+PfuCjBO8Pfz97E3K997x1ytKQ4N6ryOkdhTdAN66/RD8aNBTk5hAW
y11IwBMN6E50iDKntQuvc5WLipcoKbL1ZaUHPDmME9ExjcaO2YCdFAvUKXu5U9sb
5ZqatrMBPah6DifUwuhuGRdQkgISKidU1C7u232XKvKDtEK6FaK776lP3MUKBbkb
mMKiL4aVxDgTALV4OAY7cm+sm+OXfnkT1NgU2srP+I40F9DuyVdcg8bh9lhfOsC3
dFsz7Qr7KkIQgbaow6uD+PegeUUA95zLWMuKjj/PO+IBckrsEqdSIWG0BX+cEiQ6
BtBvnocA2HXTXgGfagDNBSQQpN0b4MDjsZ660wg0/WVCZUzFANvWgaNINtqPU7cG
iVtz4aAM5SQTsXAi8ImvD2AQnDwFaW2Q3O9S/eLWgjC8elH+unNgNcBESBiuMzmZ
ZxPs2RLl/tQR15VboswRIK2DfiSzf7bhl1sDaF5En2kIaf5RZddRMa0Oc4tdq1hd
mwSo+g5LGdb341asaa/lE4LAPa1R9ofY/aRDH3r2zqxkvhy8gQAtqQepP2NsqS1Q
/7AGLH7lYMOiMaR1brQNwnRJyBL3uDwZtU3UbnuX36rGQ7B8DBz/egM+BsF+xYrd
EUPSCgMOqWLvLkRmxmhgrAwmbrjfZdjnJ5c2hEKCE12INHKrr94RFkVbyYEBFGFf
iUYV5Mp/uRHnq8dm9wUOfAqzt+g3d4gAMgtAzCUmVOHzHGKSJ7VdaRiNunxm3pra
P/QtufbapwAmYb5HdHwuY2r97f3H4w/zUURQShwINsZZ9XGUFxwyOydeDbCTfEma
c/qLVlpqqDtrGAv1ue34twKp5YxEdfHhlD5qEFaNSPR20FHNpPZaCt8PC8PZpOrn
Da87B02LaV7kD9Xlgi1c9g1cIZAAcg2Hs4MXEawSMB3+lrMzrMvO5BxAT9HiCRU8
nBWasyKZXURTUrQyeIh9wLrUcqjDSvyvmGyDqLIEgDxuAV4XPzrEl+Ow/oRQ4uEO
8dc9zf5+xE3Jr4Z4Eq2WDWm4Fx8LhbhoJwnSll4/M+xocAZaT6WKoCN6VHRFuoVA
VVB8DIpz3FKHXXNytyg9482ULW3StbOVPXsTtTTddeDxJDJTFcZBPMTT5QDoCF5L
BxK0YkYjxdJ1pAmLjs8dRacjtidHnMMHmCCNb2gzb2iGoE9Hzrhs9RgxjpM5Xw5R
68hqhuf7jR1o7/1Zxw48175ZL/Z7zpLYk4txdfT6gxUQMWLsCWwUZ3Cftp2eqO3P
ZmhIoWaQbfkdr0TSj/flHE4FnjIZ5JfmA+GL4A9B8Nyk3UGNP63aGTyROtwMjdHe
0jpE6W+NmM1rTA2l6sJgV2sOFMcF6aVtrBE4yIUM65YX0UScs6rXvk5RDhRMs1WY
4znN1nHInDcQ0Y85/i2f/2uDiAdGTlGJKUnRG2qBNRynBBt+Kju8fKjl4wCEAKqF
N3oH1UzEfudwMaYpl4e4AAcXXF16K4pE7USDtI4SboZWwFTziT7595hPX3iTi8wH
qb2L9IXYL0lgphVYT4egMtsG6rz95O48p6ElYj0a7wE5jdnAG2ziVbNqAjLoF+AK
vRr0PExO8M/LYUtGk4UN5TcaY3/U1fHIabHctkarD2ky+XPkDtxKm8zIxWN6fQIa
KeYArfi5EsAfX7UMcgD3Sh8Y313Yoc65soj34ay3YrwE2vQ+f/PWtQySK8uMxbdE
4R6yDINTjjpf56QldVpkFkdBw+zxLXiCxL0RE8vyQPwyX3fI17WkNWqSVZuQigho
x9g3+idnJdsYub4l0q/eIvQx/QRWjuSsbo0eQqmZptmWcgfAeAeaef/B9dqNXB4k
fUpSChvb4HB+4S5rJ+dpWDnvy56Mlpe0gYwjmAPaoCMm8/zf95TkQbXoLLshk0ei
m/Z2pYZ2rTB55WZd5MUSjZeYX3MaAWWx7x3cv4gfoQX7eW81Tqsq7dvxYqQeucga
NL4BcvLPNC4/wkhCGbNRNjHk6lUC1i1B5pbvOa7ZMJdc4XSAUJ3uc+2ZVMp7C2rT
qXUmk2SOF+bPcc2eBjwU+VSljiZaZx0mkyIUpau1LTmpmWUIS4nKTeKDZD3//EiV
QDEEy47vLyakTkqt3khNtPUX/p7tPZKqGrS8FvOJtDOIbgqQxGajqiKs/F/4pTvY
jmuOKjbGGfgQwF1Xr0vOFc7OBRpnY+IiSyRG6jqVpktm5S+ke4vBK3WFTaeD/NTv
o3iIf2yameeL4HE5Wa7fm23lVy/YOWKQLvk738e4/Zu1s94f0fKQK+bhX0DHZo8E
59HJq4clfEs7GIxJ+Bwv4gnl9vb0YdWz74Imcsl6wR1ddeprYKfnYjhyprewfumP
WnuJ7jepx1myxDxD6beQZ2HMM9qdGcZXkqrHHh0q/zxTi7oygLuNq72Y+4QDHFwj
nTJTmgV4A1znj9OdJdJ5HH88XTLjvmGON/SU38c8S75q1jiEcCmF1gfkbQ+fXPKP
8PNdylFKe/6hJ/ExYtT9AIeobWcj8eGOiYXK4PxFlH1DdXgOexQ/vtVKD9Yk2nxQ
vGDUm/cIx7Cr1awQmXb8+ZIozeGW6SHHbtv8cNPNAKrRtSbpOT1rKAyLO8ADkxcp
yyS0Z8eIRLG1oLbKJr/pQGMH/0jloIEscW8AxOCYIyipWhNo8Rh+LCZxtdN2gkRX
XLsDGkYh+U5RX3JF2j4rLFicT4HWM28nZQBSCUgCSBFMtJ5DXt9Uxy34mgUup3q7
MbBpSuozjwtA5E6PaoK6sihJB+ZM3Lp5UchLcEeWRITmaI/e4nUl9zCdKqSkupCu
cHZSeulOlySoIBv2Z4jLN1PVpIwjqTdUpLbhDo4VuBWaKzXw8V0LsJkiECsh2w06
AsSN2qzlL7tHLa958YKlSEhVzobi1f8SjAcPhVLMMj+zxLjxFQYvVAeF9LHYqp77
fVPnQIJSkqgUwu8ndnqrQygRFWBFZzsZK36kGJYzCuUYta/XJnCOL1nRNcwodjwl
SFt7VzjqnCuJRtXByvDjUO4VpR7ANcXC6SX4uMaMzs/nKb8kKfaxkUhukyFQbgv2
MqGaYKEohPI6uSh/XGhBXqoymMW20daOmyVb33FNZSnl4neKmOlNFVAjOgmtWj36
3Spre8ZF0eZ1vicK5s7OSd/uyfZChvhENa7j87z4tDyhrn7TARwmTDniEmdHmIdh
3sud/M7THQHqaHcGgQLfwbJKCkj4lweL/Txwa+sQqU6c9utt+X49cfCurAw+oqpf
DvCU6ImGZCL+La1CI8jTOaGEc3/2ciad0mzl7LZOwpQpKoj5HuAAfij+qc20f6w7
+62lU5L8maa5lzEsOgtMXaGiAtJGwHwd+iOPCLOstgicrFK+Q9+1u3JiTZ80/IX9
aCscIh2nuP2NjabzdE+vcvNWy7PBtjFAsi83Ld9l/9Bb65gpuFY78huHT5zbCWRA
UyneBIqtNftWZgfvRgjEHbPObudtLnBTFJtAZ21gxlyaF+zNIGNqhIPArpRcj1Yp
1HO5NGbILb9xKiM6zzo8Bdn9gEzCWfgc76rkVDa5OkvrB7hXsZUmEHtxIpNmnoSS
xLtM2wuR428ajbM2dR2hGKNzzh7BZ8NDx+79L7BpQZ1dhSKZcaielJuILPN7Bq5o
f41nH9fm5RebIGJ7MCdjji7X+c1KCx8dV/PBZ+zG6+BF2H3r+fTiW8WvvSpjYEAv
rFM1FnPizrSFX3agVzJ0ObEyohPRQk0+0EzH4K01H3s2QJiWatfx34992OfWIUAm
5oZZxrKDbRrWNz7XPXBMcTC9xPiAoxQVO/WmH6s/7JkeUxDiFjoQ0Zg8x+WZtLYx
CCIy4IEmt+Pcq+r7Q0R5OA0MJPJmXwhgO4xrje4JDr8mSqye3S9V/mFL3eunAMDI
UxCRf/ddfLEwUrhxIrCDLIzxPUjwUrl5u5bLCy8vmEh8qAYNhJ7fQ/jf8+mHg3wb
FRPfYrnmWYYsrrK3sJGNl4jtZVa2weMtJIRMBvs0ABzJTkZoSfoG3DIWy6xqG4Lq
gQfZ/slmaVKeLdAGlDcwSuMT6S5wXWU81KDxfZO09hLT4rGuCPC/UbnJp3BCa3DB
ch7MDD+Tj3QOzdtK7yqhtGIo9xlmxOX3devxgMH6+I+1c2x4GVmVaWqEXSll088J
Kly2JqjJ4gAOILTWHiy3G7bgRsUOtOnfm1LzrQHb8j5vTSMYQLD0oCDANxnPfmVZ
LjTmBmaqMwJYdQqCIMALo+e6F6K99VsQu26ntTwQSzf+JV2jyA0gvlIsKaiMWqb4
QNaAsk86sDcF5EnLpzwyUWSc8+jhP1DvKhw2WGaS2yTwKyjDxP2NBhAgJPLmOuKa
jU9SfQY/Pa2TKleDEYUN7WTHonlhN18ZGpXuUo4Y0pHifICfR7uCRGPzf7B0J470
pvgwgJ1igLL4KG/lB+EQ0+khYr/buBPP+oKedOOOzO9MLzUe+SWMIP4bjTtohRtY
4ppoHqVirZN2NiyrS1DRXFsIJqn+MKFyIafn5PYzAB6oEv7ZcgoP868hbrG+6ESd
UNPsM49296PSrP0qFSUPNgXGkcELPK6uCP4ck4hduXGmEEgIOASjIOsJPlOJg/B2
7Lg79AjC19ICq1hFio0XPLOElA9Lpt7O08AmTPsaHzDYEEen8Ko+dbs2kQkrSbfu
dxm7ipnXfTfGSfjE2jNccLE7xPdrp2N/wi90/oTfRbJ2bTZKxlBjdm2WMlbx9IWo
NaI9wPwC7Umj6QgF0BVg2S9mUv1DRxOvwrXGo8BT6w07Gi4zH6JuaqX9i5njEle4
ShnsYgYQyr8azgPpnMuwILKZaMjbU7zUiBer1v9wS1jvv6Xy5oHPRsbANaCv295/
Y072952IQFzbBCbtND9ifbcVTIiR96xC/hVBWSeUvgLOYYsAgjYp7BqzRAvQOTZB
40yswxTylxCrs8vaSNPdy8BEMb8z+8NtcQpKuSQ43vMnf1VOfN3/PJc6R1Ly2i2S
xDLqrJkFkOqrYAP91eYXrbb4HnUH2Z1+Wvh253xmBIROafor8cg6RhMEgI/JaWzf
3K4oCfmIlAKPsyxba3lpDSIK1126+CZSJ55miUcgVTQFwhvVz3/0Rk5kRUsFlb1d
agIrofZTwRqhSb+pUEH0w7JlDq2U7uZ5Av4vOJFZuVZNuz0EZN4cw0+4N5v7BuwY
QfZl3ZVj0vxGMx+1aMFk5WWNT4S3ZOD1Jh/Y0XdUuDRD0oYmu0iEWgqHFFXE/doV
B6NRqSwKMPdpjkq+gXumB7AJIfNfOrI1C+kMgoos3itqlPU8uHvEJrm5rb/DLZf1
7f+ZOdXMPTKa2uSckrf6bRXi1d9ht4JzE1NvLjXw532MdTFhAsEgKFM003yC9jHK
B/6U9aKy+icwBlPyVA14/RIHX11OF0KA/i7zJi2mNmGHbeb6VKIHIfCzz9LBLYvw
8MFLZx3aW7/UlpRO2qlOLhjIpC8iVIvsgp9DRbv3N4axvJ2RxrHVtVxwtwrvfkSC
l3dmH8WzVfmm7ZPPdVKHy87IVx6EE1Fcjxak65Pi35xx3w1tmjiTiTslmVwvltiH
9o9ZaGWYEqn9Va704sxPlTBv8Uc4hTafETj7PX/i8vpK/dTKRlrrxkVdF0E8tHaY
s5DBaMym2UH92D9uCH+qQdHeIDcibEz/9sFdSKyYotCZR52gMGSm/izIdcYv+sjq
WLAxbJx3Rrmf1GPAtzNLODqe8U+PhPsysaIoa+81wBU9EkYkw73sw5YL/6epNG0U
UZRM6e9Bvoa5WHM+Innhu5gsY5GNO66cikH6t7Afg3yBGJQy+pLyVSaU61bNn4rd
0AYU3CvwcYwI0BsEbe1e7CJCq5d6Bh9YxMUZYNj4cC0qV2R+YeUTBKH66GmNA8UO
OvgHz5HttK8SjSYTbzuhqQjUAIhR5sTwHSGTx/iIYS6SdAAj0xZT8C6PZQJEZ/OB
MwaliDzJGnAVbuyJXareUJVsEyp7sQVfBf7RFzi6nxUebMb6yPErfO2A5MPVzFkE
7J79z0rL2pC2V/ljv8BG7h2pWQMsMNlfnlN1MAUs18IHpFdXtcOhflBR2Lg+PirJ
BBYdnI+wDlBId9hnSl2zak24yjrAlxeTdnAoO+jS5zozPFEgLnaQPmP9qAIa0Bmr
10BQbTT/fodBQKt0DrexS+C+CbM59/QkTPdMSz9oyFg2BFEO/i3kxtFeDLik78mg
xc5w9/HdbaitCkuZ9g64siolgCoIwPqfzLLD3BeO2/W5E1wodonihFwT7bmdWTfc
dcbFqksKUYxltSa7b79XsORmrWthx8S1sT8UswtZk3YI0PbTshNWXANgMjGFmoog
5Yv5AyIk7D23O2iOzTuc0ekpq7T4jV4qLfOkYjiXQXPkkvPCHSMunsMcOwq4Djgq
OBfgiWTHqWwC0+2hWmGC8eeWcUjo0VpN791AyYzyIb1OFAw413G5E1Ks2PvwY9ij
2tZKV2QHOgt+fK62nVhiFTF5Ad8UQ5a+1wmoh23c6HR76I5yqdxVW56HmEI8OgP+
Dk/GRNL2Z2myqAbotREr762TGmdAqKtZfTjx/jRDyPVYMGZv84oN+NUncQMcs2g7
d3B65MxoTI/inTy5xHRt9lnqUB7k49UyAIMUugxLpKsi3FDfmLolvGxoxvR3mXmY
1HvZG8yaRqBXN1tXUEzlZgI581+ypq1UUbizsEEbYpouO34AOjsYlpQErpOcE826
08Bn4UoxfIPe6tRVlBNJLnZe6o5+dYbXdXHSahrH4Wn6P53n9nF1dBiugtH+o8V4
+1qJd2uNZnwd4gKy0vHBCWoLxKAxTyXSxV1VbEkojRPO40zDrLeqyMOI7iJ3ExCW
gfV//NWsHDi/Z1zGWytB1ZS8rWBETCwXZZlb1m/UkMZ+qnZj+r9BldiARBtyzMRA
vuBLbfpTihLEdqhOwh4NWTyxzNFAwrNAwZBim9VqKjhWok+8gL+VVvgSFTq5j2qH
gBReZfbdFppX3BYICcGhgpxQv5Clnja6mvlxLsWNarcV8GyiDRVSesVA0MfvnPqC
fgefp9KrpwmVtTRfhEd0bjEn0i3tx3pJ5wYMnQksQFSa3XfKT3153MEYT4SzAx4J
WZyRVvsZ1jCsln4hNFKDFWcCsA2oPxfRFeFmcubsjn99Mw9jvd6PzoO1QdW7H6pp
+MaZ0caCw+Yonvf+I6VYhB2KN1xdBXbCFg6G+i352ut4MPFbzTIUnbEWGBQ26zgi
WJO9n9cFfEDuAT5uvVvXnZ0XXFPzdRvCN2nNSa2DKG8MAGqzaqfdv6VMu4FmXvhI
o4oTcwAB8bPePUXCXnpzW5Ydm4bjFtajdwh2zVSt86SUPzjBTCZD1BzfFw3LBWXz
gHQ3Dl8Aj54iUD8s7lUhdGdNtlgDMqFb+4CX1/wPOZNVeR+rLUwp5mT52K3a4Kqh
7ZYaBX7QR4XsE6VAljD3leQn+i2CN/Hdg1cP3Dg/Y9WIEU2zLVxhDAtbrLSBiQ3L
osy2lz0Ejifw8+Ld5jATzJdlGUxNT7l/epWIsWLgDivR/NwZERe2abPqAJUYck+M
STsbECLlSsl1Fduyo9s7NHgqfzAMMJddNQNe/4SLv9174bAjGo9FoCgflmXg0Mqo
BmM8S1pCa5tIfyVM2psFp41JNHpMA+4r69ZFX+ILs1hG5UidNJA269HkW4ifXK0Y
L8m899MHub9JWCqd+zHpoBUpIlytQngva19N0IygA/MXRo5daRXaXCfU++RoJMRR
tr558s/txfTRL1lgnueyQ7jd65+4KK5GNpb2GvUTMkPO0AHltOwGK3xCTVaqvIgb
i5nxGd9R9s4XSga8KAWCd8QFCG6/n0kuJrCVjGUk3gatO5gk1OG/8aKW6dROlDFP
n9OVP/1FaGt9oIy37jG2R9Z4dgzTpJ3QYbWE0F8NTT6/tEggfUUacrCTCzrMelLb
8IjLJ0KaoihM7O5FyGwPGWqfA8nnJ8gD5Lpd+bfnQYJQCwOr4/sZBJWHe8LgF3J+
4kqyIzqdQoG5FP1DdosDnWIeeL2gzdpbdCUVkWpJ45EiVn0+I/+XryIEDFjbQ2bV
WlFLMJV8hR/ubXc6wv8IydqdmZUY2giu0UTYY0QidECB5GNkt2uoo6wkCrjrxrsC
oEzDPfW4iXgLDLhQt5WMSYYThxq5UMosUP+a5amMvjYtO29Hok+oKBH7Hy6rPX1W
Cwj8Toqk9y6+/IZt7d2OqwHTLnVYSlBcIXwjkOpIEIIomiGQgZVAOuFCmznVWvOA
1VyRxY8WGU4tHEl1K9aGTKhhh+WKDBgTF1zMwJGZkHrNvGvD584tSYjPWSRld8eU
RfbjQQxtH9MOwA7EmheWUPvVGt9+78krhuNOPflUkqZ7djlWp1Tl0zGUNoEJIHUo
0VLxoV9pNLZ0moY5oP7r1j1d9uQFemoHvDko/xbWB9dasvKXsoQc1+nxUi1OILEy
qW8d9A196u6gFIZXgSPeZlJ/hY0Si4XwHkI1p3Dh5Iz9FCiw4MCJ1sgzVXxE7vPM
UpA5/v54U170Z0H66M3hBu6B+kqfduifwFF0JedvWAc/TuUlAGQ42a0gpQeY2DAM
w7yBW+bYlPud1e3IBSvFWSklk6CVTovfKF4EPF26CN05wWNfrAEtdlEJbTpjDLnW
FPBPZL8lU4/OB2B9klxzs0yu6o2r3u9weHdqLdcX2Wmw04OZAPZCIYnoa3nqBRWV
0N9NWmpMLJZMrfnSy4dSdWJvPERXK4vnpuHpHXgwJ5ppTcqqYKfMu/FG2YVchxpt
oFSsNIp3Jmfv+YHMSTntkbTvGpojk/X886Q+EQLoW6BR1azuKIIKKzeIFtsVEedW
uazIJIqs2/B/YJ05Bo/kTwGT3XYfbGJlAdQvi80/V1fJY12kAPdMr/5Uhi+B0mwO
oVYweAkW1E+e2LILJONWDBIGZzUBov5qfw57qMl2vPotNYu54OsBxjj3xLoOrs0t
QtvqsG0fuVaO6ptOwAkgwKJQTvwTyyKFKX9tsEQInMzEnb7L/jlGXXs8cobdwHul
LXPiEI3vLfNRrUtU1qMJGcwkPNFPDSKCovJ7dx3l7IhAVOrYjFQKUGaTaJr6VVz1
FBctQ0XK1fPorq4ZHNjzqVEdJvsssB6EmPozx0Pk19gtPGn0ae7KiGxH9Pvkl6pF
mua9/4OtYR1pSvEsFShyZvX47WD44O5Pr28G+cb2uLhykWacWTbNiSvdZLjd74hV
vwvJ08i7nFt6NeQGwq/JhQMFvFTzJEfUXYopp2gMbz0XJ6A3MATJvJcQG0UO1v0O
MhslNR803OMdYdIsMLX0GycfyfO2NoICT5uGEsRJhX0z/qhNnl0LhptuTFGstLQq
agigk/XhEa+aMcWetomGxRhpLvThrHlZfLpDGHMuW+ITceO/ggjV8FFvBusR5Q7a
Sdx9mfhbOP0CBD1Xc6pFWQzQOqan6GY9xIZ13tKQhhB0WY21bUHaYWTjBriLg8yf
Rpe2i3mzf2hvppPhxSJOOD4lmDxSR3YLJ+eVvmOC8DX5Z10UGCJo8/Rh2BZ45N2s
N0esR/ajUQvgfQCobMGp6eYe0an/DzyS5fLLfzWVbYzETiPCqJze6wjb7yqpV7DU
gZpqlkd/N4h23iTx5N/FUMIaoMCpIp1gm8n3Wbrbmi0=
`pragma protect end_protected

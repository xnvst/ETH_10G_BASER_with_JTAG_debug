��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO���{����<��_��Q�پ��q��vN�g�u�l�J�.- 8N���i�/�My��
_��
�S�Yˠ<� �%C9��
�V�F��Yv�� .Ǖ�L �C�i��ή��nk�	m��s�<>��;��BBG���H
G�'3�Gyq�]��{��#�[���D�7�.�H�pV����+�5����ےv��vح��,�LR�����DO��Ȣc��^?[_��!��/i�25��1��10�݁d�Az���#=G;�BT�����a[=G�-n���dM�;3~i{������!bD���]>��,}���D�4&Լꔷ�@�����F���H�҇"4��/��h��e��1���$��MԚ]��~Z��In��a4	���QB�}jӿ�Z�O� Z�?�W؏j�H���n@�kȕ�C��B�t�v����!��ʔ�6���*l�{�^��S��f���X�T�sr��Ү�~����a����I��)���0O��*J���3�����X�ӲV9�\�6�����ڌc�����r�T\�+���Vr�M}��a���-^�{PN7W�¹*�@4�ڕ����|�=�ѵ�)x�~箍���kM46J�ՋX���@eΐ��NS�O�b0'��4�(ѳD��;���d�j�x3��{7�Pϻ�˛�}��ޅ]ۦ���\C�z^㣈���H�k��0�F�[��O�j^{N#b��Y�O���K�y3�@�+�C F⁭;%
��t�4�`��EfW��ty���'c�6�h���dE����z�� +� �~��Q��}hX���ɓ��)�5�i�����Dß��S Z!�Lڶ�oÄ'rd�;{pn4�/l�T*��j �X2.d7�Q0O��<sA���э�*��U��zO�W���DD��g��Bq��&	��	���X�W�Lvv�13D��2��D�th�<?m`����2�wE/v�	S�<A�F�Sa�'���|�pc���l���w��`��]n��\������a�ɢH�K�>���͞Q��ٽ���FЫ������n.��pv�)���г� 邎��O�|r��b�#S�U���CBv�*���א��B��������n~�l�|�[hu�t���!�� ?���	�7?u&���Z3y������,�Ԓz��-�l��O����V$���"?�n�����BB��mz	�zV�i�N�x~-�����#$��9��b���3J���݊L���� R��������ʌ ҕ�e���������������(Zn����
4\߁G>�L��;�Oi� 4Ton�e�������a�R�� ��E��pL��jz��:�f�z�{��Wu^�<��.�T-Y�H0�f�-j�������[�&����B!��ڷ�o{�t(��v�5��e�p+b�Fgʚa���z�*i6�4v,�\���?O����Y`�cĎ8�~B��"<a��-������f$h�qV����7�'����[��0�����qa'�tk��q\��[�@�z������M.� ǤZ���1�YpI+!��?9g G��Q�mV���`Lˊ�wn0q����S�4�	㥎Kc�1��N�������FICo�@RI���^F��>���w'[O����~���ϗ?Q�#�̛[��{��k~f�����5��փ�<k����|��`4Sdz��ṇRq��Z���K
�1lA�7K�Bx��藀����S�J����*+ԋ�����J��O�5�������v6�։��	�u���aqM#�W:����
�n����.�1��(CÊ,�A�k6��$�Ϲ��tQ����.�V�Qc��K:�C���Q���q���z!�O�b�DjJn�虅� �s��1PY���04��5!�!ƃ'L�bմ�	�kؑe���^!.�� �A��Uߌ���a��G>+�^��7L�ئ[�n�4m�ܨ_/#�P3k	L��cCPh��+��N$��!M�9A�}���Tq��M&{	QX+�:���W7�I#�,_�Sα4�n�]�B*{����(��154�;�ї�2LY�ir)�ny��H�6*0˪P��I,Z7z��vi|o]ɳ����|2��,�<�Y)!f�t����%SV@��R��uu�l���{$�9�R�_�&}ț_�}�r��A�Qy;��T��A��[��WD�zS�f�;5��� D=	I
Ϗ���L��y�Yr��AE�{�r@[�(��?�Ӽt�:�@L�>�r�>�ӳ/�_6�+)b��w?��j����,�֛L����(��cN�f���R����,�8�$`w�+O����h��6�M����k L�x:u�)'0��ƣW�B����z�R.
// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:30 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mvnBZ3FSXi+veGaB6dKMKIMAedxl4gmv1ljWds6NChmZccnsgBuqzeDDcfl/L8F6
bsgRDXxQy37a5MK3aPThg4OFXhI3zsERNVQnxH6+E3bBEgCYgLc59tedUsOI6icT
44jAzBoQGG+FVqwJlSaQmnFkPfFjmDyBUPNnCZT86FM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26544)
drNXk+17WK45MjsSc7B3Ctjx4a8I2rZ9xn3HWthSnu84/vL8CVZ1nHt7xMjmi7MY
bL1l0rbCeFtRByp37AG3pE/UReekGZy1Jaou2q52bfhnhFNO9X6O182LdqUwIpSt
Uogsm4iGdv9IJkRf18pimlluWVfxMcpakMfpOrBRIyBYUWu6fEbsyoxWqLiu+KxD
uvWRN58DvbtaWW05CC1n/QSMIK3h3bafRfWEX5veZRzypW9DtMKxPnevC7qZrJtZ
KFNYJ90mhpbH8bXNI3GvhBJhWLOG5o+eBCllrDp1xPZtEUEaIN15PPQTClocvbIv
7RNErEh8iZP5Q9H7EiH/FRJ5hHUmMCnY40lZH912v2Ud30BiVolPK2x/mjsqFmpV
JgBXtndzoWhVU/NoAjAGNp5O3Pe92I+cjCHqKyEIgCBVvrgFM/mOfMbBTUcBkRTt
TliApCZ+Fc5DbTvG1pC6yUeaHOqtUpo6kOXvlOGWkPMFbDvMA+FIgN5QRRbzDxPZ
8q2jFp4cSjmPRkiBvv2w7OktdxYHnfWbuABGSP0pwGpWk03PWSY9SW4xcmcgYveJ
SNGIv7B49NCxjdTPCI4LoAY0OUK1Yfio7rp2yq68onJsiljrqrmK9j6VQcGQnMnx
tFpq20Bw04cULLF/T/Q/bFEAhbxKNyHA6+n/Rlyk2MDCXJ6FMOQZfG8JJbO2Qk4J
tuCPvcoh8aGTzRD53C2dJ6pTvbEVuyqzJ7xzCgMa9ochUyRyI2n7S1bgaUrUgfSt
rvuMXL0Ii6dJACIlkJ5qmbcy3eqzTxbfKRRiy/SCvXd60PWnKbatmclhbBwqSiay
HukB2Vhgf6Jz8ZZZVQXIx+sHR8NL3djPkL3PHvPGaSUz0vdXLAh+otE41eNBhcrx
X17yYK4Hga8IE0b4W4S8hf+tH5BPl4IQVQFjDnrgNvWpgPq0qBobWdYPqmt2U1H3
NzjTztcYyRXc0NrCcp4c+nZ1OiEnIqPxkm8POXlOrOj72QqNOfpCtNxqOJGXhIsz
NOgA/mwneb/zE3tU05EQD8y0xs2oVQcLarBpVU8t3lLkEmoJK48Zv4sapckHPMRn
At9wnUUa53KF5nimbfvks9Gxy3pfvK2bhCCAsmKN8TNZR86AryegSsnZQqkrBwio
nycDkdkj4NjQvvKo0q0mBoNX1K6SvW82V/rIuCl4hQ5vISI30SlP5uYnFHK2gkVJ
UD5Z8H5b0i3QOCvDqcfktFcxtw5o7yD6AHSfQyR2GKzQegzEbubWg/sVM8mRvTdM
S/LJejlKAZrFqp8FEw8wVpUNX7byMHSSddIQHCuFTyqxbYySfEynlYp78D+WMNBL
krIfvuAB0x7qgztNa7ROg8nngdhMHKXYjWJkbdh6FPJT0Npi0RRAJOIispEh2qgN
Wpnz67jAOhHxUg53aOfoiL/pGKN94HAz94yE1SQehKvdPUMZYqr38lOz1CBKOJ/1
H2RK9hHOQyOYY91F1e06M57X2nnIxwb2Bs40B7wd77MJlqL9GXqHmz0pxc3EiV3R
jAeBFtloZJR6qT1b+1pvLV4gvqBHpIHmPuV8DTFp1lWCPLTq5vINA0oQ5PnBNBww
An3tB/uE0iHr1KxVQx9I2DsIcRtFhogkDI6HjOM8DSzPOdG+TtW75ulOf/dx0qeP
WADOgm0DD5+VSuGKIhjTS8TOyDoEzpZX96IGkgYfjncu+GidUzQ4BnqlwZwD7Wqp
uYaL2aZaLSx2FgGyQbJHGDuqBxv+0FKvf/UW06wwbea1OmVIcy7wQfqgdLpXYHYO
e+ON+h4N47n4M0cLfTfCQ4JLbAQpcejSlfn5fFE8Vaow/MUEh6WXecmujfwFc7Hg
yxCY1ga76OeZwQ0MqcoZ1v2GxXIdbnDFTdjNeqeY9fpSZxP9ZQzyG56EdNEEbdz4
+B19pWgjYJY4P8oPbKKpdzj5/O6ILPoPRexG0sE1MApFrGAFp1FDaL1foReqz4qe
/XAecgAFUnQuJ1spkhkpWTomDUJg1H0lrHruVUFeEmerC77Y/1na3xjxHmToGgAN
FPFsgCTg4FNRyjg3LmxvRHiVQvUX+qEvlFfwWrhd1cPmd1SDdAI6s/XEMEMulauz
ypSLHvgHpEh1ZgPhC3guY0ri2WVdOx2nq/3piN0GcjWDacVxoTPqI8gUsZAt4Vkp
bSi+mDFD/3zCAPupV76MIR+UIOqUne4kkbpxkw69l5Te0r5ntbRr88PY7EJbHDtH
y43sB84DSaCNnLheHp/JeEf0qTtJYk/PxB26BFU26YcSE4aOIxQHV5uS7dKo5iyH
nXk4xZEX4qG4D6/qbmFMyOvzD+fJ6L0gWge5vJ3Edt6zazYvgaOu8RbH2m/67V3l
uUz50bkJ06oqscI4yb+10reb8VMEci/KVbZ6eY2XRBWWhjVh1ZOa28Hz0LcgdXiO
EpfWb3RCIa6GtF+DY9q524CYxYfCuZQE2hVrUAQ5+mTER+xs86AM17jZAjSBN8SF
07zc0+/0hWN830r2gZtvG1J2cySLP94x5sao8MyXzVIViLSjW6AHLxhVjdRPAMoN
jHipQ8xJkTLBHNq9Ltj2ata57w1da+q4LYWMQahyEuWozMlr3fpb/VEHbi79DmC/
pdd7V+uX7caIesFECQfisXxghf6a89COjYVMp0ibuD7raNa0QMr2TWV55GTuwFhz
nQyyVNvJ4S5kzZQakcqh9dCSpTZd6m7m+9MY5+LEjz95uCLtVUpLQ4eBcdyw+Dst
NWrxX5N8PYDHuSRQrgEYn/gc97fYiOe/2d4/VJbO3quWPcQBjdyTmrzUgzdVDKaR
SuHaeQkQsK7MBfknoX9cR2yeJiAyPL26rlCueUAV9s05blgoXuh7L+UwMfvYJA05
w7KTljTnzhtxCZ+v/uUZ5VGHmQcm1ozmb14mHa1WRm7tDyXAcVyOeZfFGl1YwTeK
CLNN7wAqKn1iVPt/ZD7fNtJM2HmmjV0SaqU2TkkneobqIKjiaInde0ipavqL6oK1
PVj2xIg/uTww4XzRCzixQT8i8kU5jFXQLgImluj27Um3lgQ/qNR1AaVAjuCOjFJM
zfpJxUHM6ZggpT7LyIgf9OIBfR0qxpEwBSC+zGYlCcOb9nlLfH04VvTCN1e4SN45
vwLZ4bE15DFUDTwsEybPHusgWbMg6T5Id/Iv+uJH8bi3I3Ysw0PCVFwr4jZpNRKW
FVs327HuNf6kuX6DgZ3vfdli3gr3QWcOhQxuswx+11I4dyvV4MIDlRUoc6B6TAbz
EKZVfILoQhYZ9T2RfrFrWuoWI+agHnaeTnYR1jwphZEZJGaX8vX2DOKSe+HgG19w
KcQtOZmvORsc+1N+xA/6H6eldndssssJ3hs0Sfm8Ier3ChTSXWvZUwIpB1vcNxk/
kyIybFZkXtiXWpO/+K387GpVKBUoMy28ydV/d5Hcx7VVAUcVztY/W6I5bdEBLApp
EEbnYBsmsn6G7KEN7MX++9j5X8q5/VpxzlHL4pBAH8Lw8NhhjcSk/hlmtjz/GTZ2
reE3B1eEBip8YgoEGNRT8bG4zoGqGnC3inr7gJjs8WsRp+WYGpCzynBB7NSPM8hs
PEiA2tIrKh4Z2cOXw3MtRcDcKTkrURxfd3Ov8Dk0NoZngYGTnQscX0MZdOvu4hqs
e1ZEtzlSdR825HUCSUHdYcwRwyDiUwUc11VilyuLD76YxuZV6FF/jY+XPw0OraqU
8t7lSnBIRbqD88LGS3+/3R4oJo+AzsTtIklNACZeYSCM3G0et20YuVQ9MMQJmFXK
sKoBSJ8IJr22mwVd22j+miIpOK4o30u5lgRNjQNyiR/VK6n9l+nu7dHB+AXd/N3d
NSJ5AF07jOT+H970ZEOjNcT2Qj7QD1xnwNEGbr0OOULxngtVG+qzH9GBP0yoj4Fh
ld1yfuSiuGW6XIpok23Wz50QbybUDYRVL736b1gZ7Vq+GZQk5xYT0ya4uyD11uR+
cALd1f2LJmzQBfaZVG5HpOvyicwhU/dGYP9BMbyLbOfFpYTIHxxrAfp158wg1uSF
/TxUIzNOrCAeZSIZxCnpLf6QT0JpCZL0+AtkoIZQgeT9SYK7la4MtEYXbn5USLYc
LTggZjb5+w3kOmTtS9Agv8YHZjTICypppNiPpW9FV1hA1LjevxxBoRZA44UNzWrt
F9TcGn5bHJF+smLrtYWiSCWvSZZKHgpoBZgW0/5EziQ+Xfti0qPKA4arCdpENYsx
eydP4Lg4e1l5SOGSJfhb1PHLxC9mG6931cBN0wcpfQkuJr6Ee+XLgOrBtzWpdbsH
c62K/h62S2/V36qBJDqwtjHFjWhsvy2S/RFJ8dJ7L1Ozm5MyBXzf17KmQiy/MvjE
LDyztbmNez9ml+vMjJw6hw0VfJ0cjHfa307tQIYuvFxcRcT/hwqwS1N+z1BhjWBL
I7mEYJVW9jbv6ae0FRUa7VycH/n23QBTI+mIOmRxNI5kQ/EaycZdb9Q8FsyLxk0s
oJBUMMANSWcyKTck8FTeSW9EFfxar7fAqMBl0VPOQFC+sBUTrHRpA14ZcaqXpKwv
KobDHX9jKKKZqQeqrIWQtNWdqgpfKUhRIJCRjNN5urjFcnWK2vLAKQLeHzDW5CSU
538J9/dMD2UtIOnxt1v2saEKHxwGUVO+0Jm0QXNZhKjNrwvnBHvpoAQeXd6bUcdk
jnBeQJ8w9XipUYl3KW12GIlySbpIJ/alSjm0AaQH4u5Wp7YU73++AIvjCLH4wd5A
r1KKUzBb39O1dtpDC5oHBg1xkHi2iNfL9OUQfy0OiLO7QWTcrGZA5KcNrM9sS48+
PdRNVe50cR5cHhUABw452e3iQEHzakzHnV5Olter4X4//JLn/2CWEyAkuVEF0Xvc
9XUWUFfgg7XiojuLS1kr4FTeReC9MJMcTMyxWsbXXiXfMo0gH375bI6bia6Bxh7A
vY3RXFmY+IcNyGKYqoOXKRVqmXjy/w51BCXl3JylsWv2XcVxM2ELUZ3ipOKZGQol
h4FrIKXkOxRQSYlD4qnFdrT2QUNyJY9SzvveG8V8QlzNxuSLJd+vtGUh6E9QxVfe
fY63oekEPlJLZewMpVwhH2AO0hIhvepEJ/piwXcUz1rpBeFGx5Afw/nlcD/fV9XY
gOt6bIA0Js7g5vyIveAt7c0IPqZzG2ZnYRCWE/sMlSgcX8Nwc5gUSM0b/WTF0ScT
vZRBpQdjpuvaIjMg5j8Y2BYuTIm0eG0jUuAqanINoEVeSyb6L3qPzYPYpZOZ5J6D
m+Wmkez1s+tDXpfw3qskhQGBhPjqz43kHPPc0J5grRUNr1j7F9s9v1drFlTh+Jhx
QfEc1HHFASDhkKtzc/5Mx0lALIdDp+m0i+7yvC+4DRvnmp6gQNg42b2nu5Ck2c4u
C9HSHajRpMhFKFvr+P0hWnHwHaIOmiA6yiV8ktY6wQyYPvB8yhWgAg5Ua/fhgbPa
fSb7PUiq2QdKkxblUoC5oTQwPDF8RthDDiFKtD5uhaKIehSnA6F6pf73SaW7rBPa
86yw46mE2INv4gce5UFpvyDKo88BXo94VlZVk7lUlBIrJ3gpmmo9R3yQbvqfu4A6
V/ughz4m/U5ruJaxNjMeaw45Au4PvcnzDc3dPvK7bPvVbJ5kiDMUfhbBlAePZPZg
bFQIs7NLV+uaHxtB2Kjc+0/xFo0xttYMvZqwFdUEt3yvB3dkPP+N1+RZdML5mhNm
uVoR6robtycAYlGwsou217CT0VYFq31WCh92BFm/sCggUtN5ALsuZ6xkycpry4Dh
9WFd1gO8V1M+ROxySdlBSPx8SF8nJunSQtXxQJO4jsN/Zy6ylzTwMnBRZ5saRwd+
Ai2Jn6g+vETzI4REjdYdfnwHq4JfxO6TCrNCbcmj1mb14JAocgTxL8hf61ghuGuO
uMIZKk+27T+S2ghA/RBgmaKmCTBlO4sNpRcaofxPa9nXndhkY/JoOD1kc3nVkzCB
NIAKEpyQiojrhPtJkKoeHPrNFuhvYoWl6OmoNaD75pO0PhCP62lIMknF00J7u1Uq
w4IBazPf1ypGiVFABqAVsi0Rf8iAt44p351zECTfQCniuYbCJ91X4+FoPxXS4uI8
jXRbWGv0YLk3a1+h47tNFIWiyx5MFOKekxgjr/0/O2P6khlKpM9e+14Z4GEBDuz2
4+bzRMCPwieF/0IfU6GkQtWRD9llIq02jWsZTl4gcZElpqtnktmzcvi+r7CuIDOH
bHNAM2MskHB9ZDHzi4PcX+KPM/G1pfT5JkoVVhRIVCCLpDlp2IJBsk9ZPcts2JPz
AX1dAZU4kuNbkAAu4QKLOM4yCMNs3CRCh7MzUW1TfiHwEjQChCv/1IBZyTOZKouB
4vXDLwvDp3VvvSBaYCReGfhykknFEUPa+inAoCLICROyv9DoflHTmJfKy7cKqgKe
KLr0QStAB6dpeaplDKnyUdYAz7afitIVKcduWk6HP6SPFioKHwZ6GYxK6UZ64vXd
a5ZAY4IiQEyu6aGNaQ17c2x4oXFexlkkr6EnDaaKsM1vuxq131jXUHcX7ce1/z3Y
/deBcXpSJ6EidNiNw26rYUUTipLlyunSqzVvDJ7PGuxyV5BlC2mJ/xekMCcqSM4u
mcS8XH5uIGM9mO47/DiTBQslzTv35Ltsl8v+viclXmBINFnW+0JAERwhqo7BR2me
EeWmM2RZdTnyausijoToUBZx1ddjxotV8zntZIfFhlXUWOybgK9mPGSayVtf55kl
qR0mlwABcj19OM8aTHYPqw2kbnygtzbeGERJCFLxMNcUKDE4LZZfmyqwCo9bIrZX
Jnt2s0fCuurrsdORoXBkqZAWJg/m58CAMopO4yzpK73atcbKding2Wzwt397Cg3y
bnY74UhZmCRCWjjncVJZwFm439Ev19+c0VTWfpdXkeFp3W/sU6x5H/WRKxrOPZoE
K6r5nvlx3PcdCdRcgwcwWmZI5i9f5JjO/QR248GSUZUBDQmfJPHKfVLp/nmSRWx4
MtKENO2NAQjZ9ICngcyjM9r1UzB75J51G+6XuIRgP2aCcQbP0HRBVc72sszzZVTN
mRkH8dY6p9rdEhbM/fDAT92s4TjhULoLjtApoPqSSqWgUvawfY0IOrptG9cJCYff
ACxY0mXIB9dhfe4ssYaVL/1X8CSPxIlH4Ic/clgZojXpqstCDSchUssTkjVeY6H1
QikSfshN4wYGaESW0w3Tdsc3q3k2rnUmVKrnkUChths1sbJ5ReHFN2wJEP/s1VHA
pmgxjrNXW6cgDlj3Ub/ttNikMrXqsz+2O/b7+5VXSKIJHR8YtupbsWXti5UyA4eV
vaTSAKaQw/nZQlTQR3ysOPhNHFPq7LTJLNoRoK1j+E9kTgaf0d3A+oOAnsd1JB/o
GYjMF291l2UItMqAmOA/gneIqLzZUvxMV9EWNLN2vpb85auiNaqXHJyVLjO5FSet
tN1lDiRrAy4b5dA6UJCMZ5BxUWmyFhEw6NxfuBrp4dC+czUBUg+vU+hktgNidKHf
aZmOyAg1++s8UOlpG8yDTIi3N5vHDyDAAGVMcH8sY8aCUrZBgr8AVUWlb1ZLwWBR
LvV0UZdKZp6tl/AYRmV++TnvHkOuA2eyjrZmaXXPANnPjHVyr7E/uBzhAT937gg/
uiDZBZyfDVOzfFbbBD/+jR5vyPNusyCCZP/iViVu229cU3Kz+nAcqcz/XvyTtf0O
GwAbnihbIHi7oGJx3O798bgb8ctwA9w3oSVkJCQzkGMhjh7GH39ehKNJ6Kq4uK9d
7hfEFX2SY391WHfL4uZ/aYD5ayLbzWm85q2QHAQkrH+JhqkW3Bn7J8ZSCMXdkoCZ
3Be5v5uMEFT+tN+0FZPtDFfljJ67g5oQ7y6HH3mg4/k3UtKTB5dgEOv8RTZQJZL0
7Ckod6+Nrfu0mDPgWNJRuI1IBsGoyo7AWBzhlQmu+vzXH3nrgWZL5ihREtnZJS/I
i5AGnbq1FM7oF0eBAbrytdwPPuvQsnN6op1CMTYNDks/e7g8ox8ugr64y466ds6c
Vp3eis2MZpOUDBJ+9Cnk6F1GsIKTGgWni9VCfkKiaicSYKx5GBNR8qr4NWrCuIAa
pqOIKu3gmaOCeiCszAj9eRjqlbuTM/EOuYdIpSYXPGAEK+3E4mDbk95I/brr1oDu
1LSl2XGfzxWCr8y9ZDDSN1+MeUc+HlUskb9TkC48czZ5a7ITUOpDb/GVU3xl3Y0q
bC3Wcy1BWsdV5hq07jfyMHhHNBNKgjJzabQ1cjty7Cdys86YoMLLnwVm7zl7KieQ
zlJSNtmEIzt33Xdqd7MhYhRjX3a2yjPw+kkP9a3wgkb6Z3UnsvAEX4ZTyAkUH8Ve
gTVfOaWTof3UBqm2d+5VvAbBAFph1+1EdA6vtbXcx/+a1jis7lwL2xK7f2QRBVg7
HEP9+Mn4noEI+kfuM7rZ4KfkR5vks3f9PJ1Hh7mr/uYhup4OmqCKDygR0ORiVo7o
jvSIdoZof2L6kUwvMW26IeIoNgUY8CCwfLPckkUL+hM9UWkyHFGIKsBpG43BZTJ0
+5JCC/SJrqzuQp+kuj3Yr1CwDT5B8j+KQyzk0RpQcUDdyOJCtJ4lbuFnjbQVM0Pa
K/x/wFvA3XbuszRXcuYf7gEMzRQ0VExDyxfJf6E+VMRbtND4Koc2PvnZwp/l9+kh
+gTUX7XOvhjqs4dxsDo+rNqWalouVqMmp54ugy7S8a2HNJ9AESrDw5/uGDkTfUMp
6pdKhjnzzjljwuuuJKSox6LCLS6cLlRokU1J8OR2l9WxPCBGEmLkpe+vEOi4RKNi
j+ASa2aJrGtZPmD9NAWHof1orQi8Lz7tqokWln6OR9EERg3n84YRq15w/Ns6lX+H
XZRPFzbgbEmCsQf7KgagSYOVkh5UgKw8cVg+MToAg8sPNrUY8ecd9O2z6wXL1Ovd
KlXy2gzl16i91I2criK8+K1SvekK5qUdAb6yhpiBX6hFkbNcBGaip4Ae7qctSVAy
V8nyydP64QLU8/gqB5Q2ImaTDD/9boaIyQGqoMM5+lMScgvwWu4+mC53FzJWnlne
PphPUeCBJ+Jfw/JSd7KKyovrCWCttdQpVfeIs+CW93q0S4t173Hzxz4Jw8824vRE
P0/zjYAyfFesR6MrAvhYJfhzg9s1JvoQZ8TpFeAoct0Eydh+ltUYpCu/xlm5fYML
3qmMoHkQz7PKHFWAGm1qm6Q0QaJoIvSOfuosFPJ1vR4euY+sl+NKwP7QxwrlbaDt
Ph8WrajkUayUHNw3Vv+Mp60n1BQxme3k8XTcoJD/qiFEPONExfeb5DI4IDgoyZKi
M8eoTnqPc/1meM5wIlrGjzx2itJCDvXwzPcRb0J6ZClgrRGZcgjLlJyazeDoYySU
oZ2dqUdIGwLVJRfjqy2r+/tZMRkYzfttyN1MQi7dTpCt+jZnfaWQ4F8578BoNC89
HGXJe1RvkJ2RqtfT37qipaeRe8QGtQXGENxXZrFiTRqpbq9P0ru4mLEfJ8FIDUPQ
DySGeZge0K88vx210A8TJumSGnNzTpk75XLHXGTYm49EaFHx+tQBrxspxjgCFOiN
hT91yyOb4hZPEbQ6FNcEz2vL9CyvRyLxtD9g8dsvtCNpVgrOuuErJq8tw/uPMOsk
1sF4gdA0I+3vmjPuJ1VLuw6KarkG4vUavIW+1mIyQhwntLhijh7w2+MTd4bVlC1v
B6u3i3sVZIhSnrCVpCgkFblFkWl4iA+HXOtWFwXLlY48UrjnNuzShMloXmw4y9Q2
BhX9mxgvhQe+TF2oXtx2Mk9Pn+Dr+aZo3kgY4a0vPKI/9hzAdgX1WE3BjCd62rd9
0eMZRJ5aP/LWF3zSVwTlqFOKm1pm2KW5LtcfMnmOI16ejxuqlpxNFzwFTHAxcYq7
i5jYNHhfvf8OjbIrupgVULzB2mgBQyirF6uC5NLndB8QK2FNWxne72SO8Nl7HqaR
NPZo3+eaQ6a6+1pGcz9j1DAiiTmoxtChCOCcKOxYIhsD576+tuG0IXILZvsXqjtv
H1vSJau6cPYUuA8EqguMda+cnSxHrdJB/tOnDewRDZuJok1qfaKRqc1AH5ju9Haj
9iwtf0h2XLWvmeepA/IksJAy/3EyNfvE9whTh7sShNgPzf9B8MGrcSgCMCskOkll
mMrl+yBaypdjy9XNFyaXcB9+7t53W+p9mFoVttw1vMjHIbUjWBTdgV1SEqVURsEx
nUZfB8ZycaHLH8E2FA5tEsTHLJ/6/afQWcRC0Us79rdqlQjuLoIbKR6LfZB/Smwf
5EdWDcSPuk2CU/5lNTdCN50n7Y5texUl/FuQRyO4nN+ohhKfc4O1bSjn6dEEiTAh
R4xJE6R5iWNO63UtG9pz9xZD/fmIP4BXYUyBe9AT2cGmhzVTRvzLEU0LYjbVSUla
kbH0kHMvKk4UQbC6EoBWGDUGtNbhxWkzYQpDaaoWkgh5+z9mBsJ5bm0K7NgBn2Hc
WqJ5wj5OX2uMClVu74itlnt9KfnrwuxKI1xXoinjPWNZbnWGubTOlF1ogRONAs+V
Vda4pjTeQMGkRPCuta1bsGHjSQ44o5OkVH5sXZzIjFI8oi2LlDX56ySXJpGv72t8
dTBnsK1BYJKfcDoaS+On7c7ohHdhOTSag/mOw1iYbmccvI7N8w7Y1wZJZim2n6jy
PzpJi1tCIqayBrwdQzWbZ/EFwAJmslq7tLA26RS71CLVAtzXjZ8EXDjjYLXa4V9g
NVOcESi4pnhJGzEh3c/8nB2C9uz3PFfGnrSnQENY0tB3YKsiLBCkt1Ne1RtWfA7a
25U6mDblPWaOhu3oB18zaR/Pol8JEwcvfiUV1uZBjDZnpZJEA+xKBY1Y6wQC1njc
b80fHXOguvGH8KXDNwiA0HEvMCftmNlg3J3RQs0rJeY2KW1lHFRuCIr/pBL7sfAz
Ebs4qY32HsDltjftSFxyxdgDbyuPsO00sIakaKyC69zynN0M9JDtXSzx64NNUQSv
TfN0o01Xhw3lD2GrBXRXfEd44NZBsfYzXqZfKVs2cqxIMu02LQ+f0KnPia4cTy+O
9uY95cqahex+mKqCUnQU63vizWUVMadPfJrKbMwCbfevJHIKYaTA+u3hsNZG9YsM
kT2cTCvXCPH10E3Wa8hC5LoJ2rDjFqBYi1xImNsk+XKuNno5gnjA+TStd059C7oL
aICGjhxFvBe2jcpCwSHgKuQDXwu25Am69gSi71o22zk/7Qk1dmmsqhxvGv/TUqrO
zkkd0R/9GuqFj3TmOp8zZDmrLbzTmK9snXiI8KDSoRgIXyb7S5ZuTfUjYnmHs0Pq
9KHC6iBVzxoWd+BXBsCZEQOVDTFwwFBdrCNPRoDdALTkdSl/YAoLAxXWjLD2ghRp
W29T42uThe/E6wTfb3uTeMbqJFEpDBeQnv+ev6DejAgSINo4VdLNMoIYRXM5wXwk
z8XXL/JeCMq7EdTQdIj/gcbheeUMGJu/ml5MivmtnjVPiUCTYwTYBm3VZPMAKDZQ
y+rQgFLKTliPW29O3rLyZHFUJV6RSpvei2FCp2NIFgJrRavvDNJJo+vo0i/gy5SJ
6bM1/bArlbWnKWlAGELlGz7ZcAgINfbaXfEcBYM9zmLjIwi7o19kjFlIXT5TQAyy
BGu2TXkhfXGTmSBVxofBbFU4BD6CChlXbfHFp1QuEdppWQp3aN5XFCa8D78bNr9m
a6yPxTupAUxrYKhfOCJSQnjExL/udNJEgy0BiCzks12ZIZ9J4/4x/7Q9lor2LOr4
/LfQfz0fS0CUdiJedXf1cjGGoxfOiXlj+1f5jjd50fZsGNJQH87bZrzpDDM71Izy
rIrB7j0JpIVN8yv/5dhc+UN2SKfO48iKsZfgiAVZtt0Vbe6I+JEzvCLscFfxPLg4
fzxxJE0hVDKGBiIuW9N9gIMegBxfdN6ibUr1c3IptK6302//0obtav7R/aTxQf17
C7mvFYreCjIOWAh80xHGkQkJFOQnUFIvZ5dPFyayfLRdrBChd8NaspOgP76SLu5Q
Xro60NpPTEFWkW0qZf9O1GZusTR44PTCBrL04wsg0DP5J/cgGG2iLMkJ7qVORvr8
Jlp5lgOu20WPfSbJb1xUtDoCC9u4SbcOYOc4pQ/3EkS0VE68/n8omUQOKqZmkvoX
MPMYvvs84zsv06gYX1BkgrAfUG87V060qgBfsMtNDI8yz3c4st1gmrqBtBICLtkH
ts5ZK0QAnU+4TR9SNcHloFqPfSRng5JucUCor1+PCBvHC7U4nnm4k9+2LrEOSFLI
n3zfMCN0EU2eX9LgCsCHLHdKuEJNZA5H6BjOGqh4DEKotPDsMj8eJiRckEWGbFJ9
sae6gdoizASZuyNHQOYojjKZA6ZVL8DCUHPO6YrdMNFvndaNgRkH3YB+wWWRC4Ie
t5UZCW53WUxR8bZXS4KEE+ZoVm49YW+kun1sn6qral22+QN8RGLJWqaq5T3NXc88
FU3gcQn84MvzxDLMPowg1I4fPIPe+Ok4s6Edjxa0Ex/ncbb2mcagr86QuSTKBZy2
Ei1Wish7Hc+GcpIq0oO+yr8tIjjBC8fcK6EgcOiScE1bNkahM7rA7H4A3WuQApMK
4J+1BpusIBZS30KeNfY3OPy1sdsXD9MkwhtIxWrNvOJV8PCBwqjQ6FDaNe+XU/l4
Fpja3EtfAy4KAnkKzmx6zKIOpj0zte6dAJSpQuQxb5grr5F5kYBM7cYFkEt/jFFV
ZzOkiNKNLXrpcMNNS8GKbA57pxzKg8zs1FnlBzY5NkXhGTeo4GQpGUopKFY/E8nw
aZ656+meI41oLcf3ZC+O6Q+518qpwLlVJ1Dj0NmX2rKxrlqq2ogxSBDyRi14l6Ut
jCoI0T7ly8Ym48m2O3rXz8RjvNFZ6EJpT/xYJzD5/UOPoB4gHsvFu2PJqBC9FzJ3
QtCsEkS1IsgjKflYzhTaEW1Oa1ILxb8u+wxJSeono2tgmMiJEH9dvgKYmgNiY7J9
O+S58axYeADQNK3mt7a6T1T0Es9twYdHda3gCi5PFwhcfWRWboEUsXaayUJD0h22
gFtd68JQON17zM39T3GU4ZzNAXLNDMbqlmKZLbuehxC/GoyFW94PNvdDCbMnOP26
MWO2BwEQYN2N3Kry5Vf8ktt7dMGAFVY9JyLkqZ8tM45JbGPpOH7gcnqRwfY0GS/O
4NzTAvdkrY6RucgT+Rr3vyndIo1Z6HiypWB0+RE2KYQzI+4xcDQmnhML9eUy7shP
W4hwSDw/5YRWupvTzf0aAr57B6GuqgX8y/eeNn6qZzgGZ1/wi6cbKdLpGTqpvqVG
AU4RAHKVM/KLTzTQ0n4Jgz2kn6JajfVuAGQ2M0MF5196hLr0O3yatxWUHaib3qwX
sDz1yX9Ix/69ETv+ehsfotNL4I1TnHQX9cgsCsYENkS98Otvsc5mXh3odBkkxHD6
EQBaJooDltJUjbp1uIuKybH04wvIsUCk8O1YLSqDz5o9vUYOpsmxiZVyBYEBASvb
6QP7tk+UKiLGP9ixyhHMCbor7hcz5I/M+WmeGaCICenWn3n22LUgUxdFSZXF8dhF
XT6XKTC5SnEIqJXO7iEyh9SHDxZfVefwQjVGyg4nkR927FJiKStnoJ/xU1bLZ+eH
nSXAUvjKNelgWo5uhzkSwdUyqgSwi2yv4u4QQSsrKgjsnnz+joWxHca+9v308G7a
nHLh9fMaM5avnlGGh0zfgAVxPARxQZ2hM4x8T/bZMuZ7zJ2f0PqarC6dbE0fWgCm
ZU6+3amRYNkb/q514m1KLpCHFb9sx5MHwOREZ+21EU5jzEctqQ7qPhtPhA94+rbm
VL4Y3BcTbnobmV8+RPRHy0CNbuQtAcPCXXY41VVGcrF9ycfMysWa8+dUbcN4rQyQ
FgP8El3MJLy0kNuoWrzB5vED7HQDBPC5MNB6Q9hlorBmXo5/fhp2NM+nLrFV6UTy
flrK6Jn+Vy2VTdjislYww+PqK+oy+UZizm+T3vw6iAoB/1Lgx0B0nlXzRqQV32bZ
oPG9+zfNG1kCx1GOKpaM/EHs3Y64CquniGyKbGW3Sk4Afxdnw+C0yGrsdbCKdfkG
hZtVzA0IwKJJmn6JEXdb0d1T7cZE2kdJsXYFhrpfsRSe6ryXahRcWA0m8gah7Z9u
bTHaeKb8k0QzWutlU5CtmuQRL2kHJo1goQYeacozf3blYf0ZH5HIghn2+HoRVXCu
vMmNi2BiDClOfxAzgIgKYea/t2XzmjO23UQ8jIEJWLy8FumYonC0/NDI3lIV9UOX
Nln/F97u55mhAs8SvVXyH0UMIo2+jIULanFPuw8EwvQIDJk5CKyZULgj8BRTOA/U
vVxx2r8p+s2rOxYZ1sWDiLfLqlHV9nfLTbd78+GGm22qrXq/asnEeAb6pI+Xc85w
PwGB9B4fM95MExVyx+9J4OdQdPwOt58eMPpvc585BFe5TG2HxKTGfMnidFldNKJT
J2HHU9qFCozUZdphJ6snRWdciQjGghKYJLOIGRR8rhOWzWZHWz81cAteVj+4z5NN
YOcCYZyotceA4bCugGJZbdeKv8EosedvGsl1i+nTWm6azrPujUwbS60Ow9+FnXVB
r+Y/H2pSHZfmI23Nu0xzpn22INaWkN6myKAOvwBEUCqjoV/eM1THSHY9gZOthn4r
T7/NsyuzTQ9tS0OTUjLrCVCg0pJuKcvFCG7Z0Iry/lttHeBwnGCacm8jJFB3eFCI
x9Oe+pcA0MGy0d3+vs2f1gcejS/2OE/AMkMa/waXBkNmTssD7G8Jx/zUVPNZHDzm
2CRH+/YFxm1h9ujYYXvY3aMNCUQDUHu1A2S1yKaOTOkou5Slv0MusyFL3G22yBGm
DTb9+HJtp5KHR29h484AOaZF9bYNND3Wxfy1SY53ughkgcUoe/zTrZLrpUqWu2yD
b8Zjc55DRzrlSr6gQgX+6dquE4DizYMMH2K8+YsLkyB4YfxrECBoxCAPJ40+SoNU
jKqiQytIJ+kA3XHD46i8tGMBLoV7yXwoMwKYnRslVcYgAKIa06NN3n5RR/whO8iV
BTuaz1U+VLtfGbYK2yF72zYUz6Pg8IIrfQkgja+59OKOuPgWfg0wmRnwojT2Idiv
tfK8qZLfi9phIERQi47hyNxgUvoWZbP8zwISjTpWw3FV+3v96TAdGiJyohQSuhUk
xWq9qvyBqHpKSNNdysJkuRRtJctQyEhzdq3impMHxkjWznIQcpASFDw0OZVJq6fN
l5ivpJAILK917QSAhFcS/oGKJ6EGyZP13GLOl2XKWuj6raoAdUgJHSaWg/LwiewE
stUz1cH7jjUwP2CfwyFYaUpXNnXaNxT5X6djdU7ALP3+eBkXaUXQPlvl6iRqxP2G
wS7AgIQysJpWfhIQVKJgFxfEt3Ld8ax1o/uWeOXKpsLHbaZQQsJeN1I5LOaAYoRe
LU4/F319Wfow1F/aPYO2elxMDiFmOfbDTwlS+FrFsyWYHFBeVmsOMruNe8cOUrHc
sHW27MlUmQafaGXGYV65OMTamquf7m/9CYNzM9DAnZ+3KCrzcBqrFCFjffsNRFFa
1KjQsCVnJ3W9RWp5VuJ2opW4nOIOZ7xdc500oqVTyTniYm8fuCExd9qrISKc2GsC
IAIDA7iwfH7s7SU8s198rxlTJiUM6Rw0YEIN43k+6PrIVTtUGhRMuAwotGwTHkC3
yWJh2yoNfW8YiB9tJ0DFJWfucf/MrQ7YbSGCynHM2whYFuHBLJRhtbPPZiPi5g/P
YV41YIBptgBA2byaxMl8SWsNyShQD+fcK3x2nVBdWEIyZcZHkrY1xjgulNQr8dLh
dYBKAcRFioaBDz6vF7OO5WJxVlKomLULGhh0i68YHtkIh4KWEr/IvqvhIaP5T/s8
T/J1BtqO8S9cP0WtaC57FwBurjgBn5FCo/xmMeVltf/vOOTJMLWHdSVZYYHfAgxZ
7Mj2czOXxjEo3beY0xFCNSg8ZkpFEuBahGUMvI4Vcaq441Hcy7rh2fCwsg3XEd7V
bQBW5/C8ThRFN2Fws1sDxdCTZJ7dHZJtTxgK3bGtd4tuGVPu5Z8wBEECWGzjWSFN
quIqilVx4/ne9OL82oSnn5sCQIfhWp3tRzXm9CxWvwIkTfaxf11BcZc79RnPtxX+
IDraM9saePMQwBcUc391dpsqQKA2XVzGlcVt8I/53ktmg7K3SuE6uSX4Zp+gEuge
lJP55P80xRSUPC+6osDHOQT7OHaEh45wjRb+8PC695rViYqrodxJCcgGN4nEG+5a
m1An7scfoTrohRWlg+addO7q/wB/XK1QQ+3Ouzq7G7JzgSsETX45LWzL+NtPvSfE
S87A3ShalZ1Zmret5seY/J24ePoBTocJqhTY/NGUb/gy8pr/ou+OCNPH4M7HFmtc
npJcw11tzc1IkZWMwFcH0kd8XT25ohnwBhaAFVPSFcw5Ckho33NBOfDEvuSuL7c1
ugvCJQeqXp0KvKDEx8/cEdl4qIxO8Q4Q/3LK/SQKWPn3+D5mU/8YKK2RbxF+BVcp
W7USMwT6/l8dzOIfMuQTYQUwTGscM44gykRWm1MHQDyygz0NvIrYHkuzhn76SyZ8
o8jo1NQ76y/RWb497tQoveJ9xNvrpYTcCqneXPQrHm9bHNe5tWBVZI12Dncv13SG
1bhGFEOlCFLxmYUeVyhCYJXHLVkgYcRu1AfbT1G/gzD6jQF2Oq8okwouZrJI/aET
8K0J9bozEb/1SALsUUcZB7Ysy+2+ZbHDvXkGyEQgQfrXE3yNVhwWkdxek0sJSxm6
G8gDgvJBf5GCH4vk5cuD/bpCHHMYXG/XuJiFo9c66DAUGq388us8nJ7H0i1cOjFu
+5o5OiMdHKVTDMdSUwZVS/JQQiULwbobt35udQT0cs37sZtjscqxAZCdhtElxaer
+fI4gKS4vbLchQpvM/T0F0nP7uX4sSQ/3SIXdkl726iam+mJHlQXTykmIOwOeo6Q
UDKqWygPNmxsLCsiPkSVAthqLeZihzZob5U8jTrUGLvSW42o98eipRUD1cXrc3xP
kMNyKxJq4WwsSHkyiOgR6VPXAgrIqP8utqjcNLmXKKNAUk+q1rf/9YoB301e99L7
04YJIIFC5bu+cF2t0cz4oPuV2mSMxMR4ljZ8tF2wqTPSimABVHC9SVQhtIyDM73o
23XTONreDWCulxsWkvCSY06dFlWGeFWGxAZI0WWFy2lMhLrENn2xoVhOaT1hs2TJ
kePi5AP62YRyxLJoEZxjj98jNcgFSeuFniAPyV+IBhpF7aIpu9q+6B7PONYCNxvg
WePiXr1O2kU0NOgoqKUETgvxmf2+fh1AdtDs00UW2erXwU02FY/Xe/E+dHqoJ58d
hfwzvoInvW/qLjQgL/mbIeAoVwBBAKqfY7NBn2cPLmoUcQ3PEbaKQbdqVBdK1RK8
vZMywWqboIrytJFgNtHXYyplaE3KE9CZ738VUVD+s85GVB/6+LMYIhfwAkoWXp1/
MFaIXhwbRWVBKrEPty/ybw3Q563YiO/XUp85/FpBSQtsBHc8TYAL3mNAnyjCyZ/K
DS57Z6UZFm3MaGO8PDIkIWGx/uQJ0iKnp/Pg0sPRfYvQBUgtewET4Xc8qE46+W5c
omW6ZArZgmUWZXe5oGuLkzblEYpuDXEcjxRXhsvjRQPLUKrec3p4yU4YVAGdViD7
oRhjbbxfDeOYRKhPgILxhQ7KcGcye/Fl2cOygxCayQMvxFAOc2nn1cquri24W2bT
1QB5lmkYjjZz0fP5P/A1ewLbdshODQYd/jc6sI3e5k7/4O8zTe9xJDLZOwDkwTzO
TizazslsYp1d4oE8gnJv0+hBybFCyZUXH76Jq0niwdg+fnw/XGaeD8/l7Yd93NX4
4B2jiOOaRSOuxlj2bYp/0HZWba2HaU9ivfUYFE8FWjt92+WSmBgJ+upL51DmtASd
Iz17b93hjgl+f3rsMW2X9GMM/Ez7chKBO0xp1NAT8Ic1C3JvBXU5Iuil19oHIFeR
+A399MlDzhxwlYsLnWJg4wnzxS0KSns/W5nMP2uOxYop16mAK+dw6MS5kyumy9d0
1//+mkznvyi0tBeWR/gQtgoOJIlNSrQHE49PFVqicnIkrQC+y7jgyf6+kQ47EVjd
QctWoi9NS1ZsUuCoQYsx4uDP6uZx1ANyjTPndYsZUu7+qo3+OCcRyMzzucUwE55d
KJ/c5a4b5pcE8x6CYtPirC7j4X/eUw56APGvE4jqOVZR8isVAL1DW07fC+TpY72R
zDULrPup6XqfRSBq86GwFYivzar31tgwhejqzGHOJctlnMQLOhvAZx9JPHDZDhAu
L2j94B1z6Zl3QC/FQLZBzc+dIrPLWnBktPilePLnHO1ScYEX1LDBbhOrOsLFnuhY
iYeAnJrf28/PNHzwFyooECyGaQty+gOX7217oVKkiZaZI4iZmAw/c3B9mz2V0PFp
nA9wL+Exo/Fuw3h20z80oZ1CVF1cQ1JtCbedWr348LCsdDhntNF9oTfIwL3NYDgs
Vngx6xCojAam7ue6CXDhgPCGYSFgesoBiw6b6wHpjnZ17M4pQ3nYAKHYbnz3Qszw
Z9q9YOLulaJiaCAvGpi87HGecl7RtBk5SVXQDS581Kp9G4/Haz1pRWOcOETCQVkw
cV5r5Weh1/NVFWO7IQXKzo1iRZ+4+BZaTVHhWBcpuGAQwAMrKCptpCcvAmwbbNj9
JtmqjGzjeKdR9hknwQRQDJGO9+ZNB08xcT38n+UXdlOrB4lllFL2B5xMLn4XD6+s
A+YrjHfJc8/oSCe+chdexIDnZXFfXEF/LNF1Klu3r+hBcdbXIYMyrTbKsWCdBPuJ
e86mO2C4I6ltMxvZaoSWxhFOVytVjBgreXya/b70oD9KKvgW38cYMcVz87kxkzpi
k0Lj+uUEbr/0f/6XuL6ltuKDbIrMFLsFDhs4/qLuxei7HFOQkvFd55v1aTWiGwNM
9EW4BP+xE40+KzQyAn/IzX79TK16ebaxrLMkoXU/NZYWjFXf5xUqQfpFD32o+gAm
TS+X3tnHrvuD9PQHdOSY81rHJm4baGtysGlkRr1+fpbyteefgkjniQLG4kKmEGDX
g8a3gmHPJhO28Sy3ECLyk3EsJRSNV23DerfifJieemyykBJLy5C3WNpwz3yvgmQ3
mlzBm9Saq5PUFSo0iRiYrva25nk9YopsXL4WH+Uu/DMY2VEEfS+oW1QhxjtMtPNJ
8yE7yBtL9cHlzfwvMJr8aej0GjWY+ZCuXDJgmJCwBIUODTdtYq5nkCdXP0CqG/jU
QFTUmQ8ZZCSpLzItwqYulcHZDfLnT3zeeZIUcIojiCBvYqH4zstCUZsw/AhifV/1
sOnTIfc54CXZrm04f/UnyfbuKGwJu6liYAxBIHV1y/ptW6Wb7jTt1/VJwTJpHUKO
KCgsjIY9teusjqrzCDrtFcJB+r1znLgM+VHGvtqb9ujd/AfnQQNl/cUv6FzDCdeo
+hQFAnG27nlEyQZ0CHotH30ZlNOuKZpqn+K+4gV1TuKInfPlww1exY0n9ZCtXJ8Y
AsR6e2+nVd0Ccm8qgdZXkAMs5h9DZBYSb8pEw6R1UOC7JpxqW8caBYWRA9PTl8Jo
0RMQ+tiYhTyR9z78fnqpH77ZzqJNc+E08VWvMGoUO1WVNt9Uk1EsdwFv/WgxbZm5
8NzrpknTNUcWyxDCq/vnc6PW7kjUzQ68Z+YeP4Z5PWmegn244JGY2W59GjQHLhl5
VrR59M6ER0NVOnXYNRoeSU9Jgnexjm+iP338SW/U5GvKaibJBImpgLCEqp4kmyPu
gfJru2TH86sTTdbvNqu834vLUtCOFqH0JmFM7e1sg7AI3Ax80v7xh/HOPbQ1Baup
ID6j9dD6qd7rw/FoBWK2aV/EJvPyaSdUNulag1K8itiCipjSU0gHarfwUP3G6jdL
zZtItwR1SYJDe7W7dA7N6Vtoj7w58lOuaI4jW+k4w7SQR4TvKB/yCgs7jXHC3UnW
OXNpgwmFR0Lhiug5SlJIsbSzMeqeOBSYoFwDb3wwOhII8OAgYOu9wlgt9U6kRzsb
gzIf8LUFqxvm4cnAOlEqDvHysBPhOTbUcDKbyzxLk1i39GW4vAIMg5GGcyDsC0eS
PeWWj8q9GBHOy+bSLALnK8o1ImW2jugB83iHAz0ts3BNa+dvhvypf63kMC7lcxBW
dNOz4o1mIOKdR8IJwOopWcoHV8LqFCsAJL6fdPFN12ecTJI8dwLsaJzmd7pXA60R
NDJtKIl/toKAmlGADIFxe0jX+dkRlOuVcGM2YUEj1/M0F8xRdD4nvzDxCBZC7Hyz
h4g2jehGV1aWKFSyUCgTyIVDp1jNr40C+iMSacRZMm7AEmw1kovo6WgFpjQvi6sj
rFhb6XOy8NgbzDNdYB2nws+mCMVPRXsHWuogHoTx+ZLmrBd8bzdjOueQtBciN6/k
GUf0E13XMlJPUce8ELras8/MXEB9/T/daWvDqZw7mOOTAb6Giu24phBxyvCLX5VW
s4FR+TAWSntbuJamngUdBVSmH8enE4MvSNa8amqmS9iiV/ZuBNlXdKnRl3+RmAOd
LjfwYx5YDHjmZD734/eRQtXXbHZViPSf7PCjjBHJ+NSceeUwuLyRCz0zuygU5dy1
eENDxxfxiLGw+Mr9/6ZzFO5rF05HQWNDqiUp+HmuOxo77BfDD1Lz6auM1SoRkdv+
ckznJPcsVuC8PKxb0cqGKVyNTlMJt7K2LAA9nksCaQ0xsJiG6l8MLmVUHEW90xrb
j1df5w3sq4yY17yAf/e8RQHfFxNlutapTRfttflc9E+7gxbhrddkNk9dgNi7zI68
hJn7uHfGgQD2jZfaQ2jDeDFolEftTZZ2l0hOw7S3B4b8f2JToQnbEqYfcaNmFijR
FFFdxSwPMDqe4YzDu4o0oTb1dnGbZbFOOq4FoEpbwIALyoKGHSzqlNuPCIgosYn4
xdc7Gnd7sWSKC379lwBxScPN9xIx9azEDr584bShcu9w0Bj5AYxuoVpKVEebfoGd
FXpkdQ+qM2gONc7/PfpaNs6ulDnTncnpgQ6ChSz//ftyPOXYWD/rr0FG0CWe+J5/
KVgJ06F1fFy2Q8WA16XGdDHJeZZSMiw4O++U/I6go1YNnPjSSuKJqWZw9jJzKWVn
RfGqFy+H3D39+06v8YLRF/QBJ5n6En5Eq2GoczlVF5zm3xfCt3lpluuyh4Ar7Veq
DilRVXMyK1s5AqSztZBi+BD8zjxqEZzk+yQTH1GsaFsxw/nghHOUwJ16Jv3kPxO7
WnoGkL0XMfNVrJwqFGt3ufsD5lSLGBlKASIAddZmpKk/Ed9ljx9zIAzAByk0fACu
TWnnr7toTjupBONqO5tFTAivoBcyfJzvY/0oEg0rHD9OPigqyTrVdfSOFTCDhRll
UqYNa8TJMaBWvIGzbaZGOveDoIeoRsjY9ziZyNTbCEVYEvLwuuiHRE2WQSdBXoEK
cAdi5SXRWIK5AP63TM1sHMEYQNXOQWgbWalNu5LvBBSUWpNYQUywDzfKJDA11Vqi
sT40IFAT4/aPBAp1n3mA9DKCs9rKNcqokQ/0TD1+5aPnP7Uz0nliQZdg4Rrk54d5
LkXwoDXV0jHLm3G97HBAfOMhAxOMGuXRiyiekQJxcpN94HvCxNpIlxCIiKOT9iMi
3hAlS3bT8RfxvwD7sLv2zzvDzZMcXt6hS8mOe43T8oS1mlQmJ7IHp3UXA4nTwqKQ
Bosg2BCUAHw91FQAlH0JYGjH6EDjziPVm/2F/hS7ou4qHpWo9gGkAd/K1TLH+l3W
H94euqMNUNQLS5eo63+az+MD+qywqA9Wqr/gNBiEnj5j2XUFUTkN2sFQpOA6Jo9K
pC2RJpTBAtu2E09LSDumenvuWnGl7lskYe9KGDi4UDEoG2IKc2lscIQcpMKOyhDJ
PNaVrIDJ1GYge8YABZtRVilMBhGfKIOE/vj9mDVGqdd5td5P39xIP0f2TIcOTyFJ
QnET+0w5BL6T5cw/2SNDWTGUlan8KxD3J+fuMbcEtkb8nApmttqpdqRBrdu4ewQX
oQCqNOr9Kl9794sPNC9+EjN8taJ9gl+APnfH4sXpPEbo5VoXFEdzuMnRAXjSVxOa
8gIJnZSULyKf3J2Hb+1YofsnrxHVMugxjMwM/is+EC3orJ80kUSOi+JxhCuHw6cU
oXM1jZYHNX3LD1k6jaf/NVBoA6S9e2m961FVzXmv9EcholVWEuLF8xTyXNEjVz6H
AjxL2DJ2PCV7avQVIev1GtQ6eed91/d0A9CRriAURWg9lkvpfr/flm5JgSj2jvYg
wFto+zRBqrMKVD7Ec17G5g/yzoeGsvWRh4Wgd7g1Cmx3m4yiXUDJIrGvQ6I/PLMI
Fpfb8YNgxpPta8e3P6uvujng/bLxEOdN37bGC9smyKm5y4m8a4DUCdgK8bFqJAKq
s69kFuvPo/TZ538AHNQAy8W7QgHGtdCoSfIeyM+Vt/g+Dzv0Dz2pMqAeJ1MwEH6E
UWrTAU8DFyDIBbp+RPcaZR96dfzoToKj9nVzSMq9zKy8yDLXYAw2cjHDCybXz5di
cT3m51QkrHMX9AlKsPpy/cfqj9dPhH0kKNG61kYeKQIELXrzW585T68HyFYE3rDv
YYAdNwWokVpsnuJHz853ZUPmdNtU/VFHHZjtQS0rG8aAcyOqYwJofeIEU237uclU
2XS5biiIoBVtAmfZi0xBt3sg5mYzy4W37mGMMRLfcwK6tSRDp95fe2Ztth3AVg+k
Fu0MRBz0GIOudE/sizWfwD9IvvcJN7+P3NH2GrcYmd1yda8/7HdZoSt1ITin0TuS
ADENlSdl/bnNuQC5OeVP90jLwHeHx9qOnYVrgqDX1Ydhd3C2RYyaQUl5LcWzZUKF
a6XQe9tA0BjYIc87StvqFN+SYJs7KgJrbr5GClW/69IIl6jXkHj0iA0Z1blTTfbj
AL4XbB36DLac2Sm1uz2Fviq69v6CRggttcTfDKj4HFmEPxYOS2XZpgCbQwu3Uj3T
JREC5Jtw289M5TSqFBzxYjRp5N5TsGk8ozmlHS2/jCY01KWNJEXjvY4Mb3bZ3DZg
m5RxmZp1vaHzVu437CX+nrpk5VqlTC0MAY1cKvzuQzvHh573eJsM0fiHAfT+KYMv
RL0lTeWG9lXf6fiAHukQjQ0xJQpE508J0SXD2+jWogYtAqKfqcwtpxO1VFkwA5HE
9Et9HuO49ZFDHu7g40wKhmQ0+UDxTm04ShBhcPimV037UvDkY9+QC/gaTiZRTPwG
QQXgWQbcsv4NVOtwzYj/zI+1470+tvRDSdyPuafhRud27e6nQ79A7nup5lto73is
vM+/+lEFw6STCakQnpTQvC7c49m//l9FQl+wCS+YIw5owHM5ExgleyyLo+2orsYy
c97ioF+cHljCikQH+DUGMOXJF7cah1K3Q0WzuFt0/5333A/Nb0NiJ8kxWXsEtZuf
mxib53MkKmwRmE+T9E+GmojrHI0/jnCDY5mLMfyrP4kd1dS0EC4v9rX4Umj0cTB5
L4wg1HUouIIuDBwSAT7BrczUoDrvXCiEtm4Dpkufm4gnqwuf+idXmlQ4gi1Y3N13
zIglhz24jY5OnIJevWpk1CKRwxtIYZ0z7ZcCqf7WtBQYfLp+EzNgPIu/UfsSrXyD
95xj4H594vtaCsvFqqFsYkxQGhPwCLqKJBOqPxjVc3ytg/F1g1VCECLFiWg3Tw58
NW5rRHYgVbzQVlSUph7kmVFN3hT18clqCakmLG9w8J0DE4ZBT2QQmNLTkHsVT3OH
AeDAIZKqIC1KsyEN//2BUXWdl1Rxju4PMC52omwJ/9gKxVQcn9g6p0n0dgRoxRV5
TRc5Y09vw4vks0NxA7Jr36ojGTFChbCRZxhdrMZWXKOTU2ulhShJbpvw2zSZh7AZ
AlrO+eTVY/oN3rxeDbkxvja+qc87Tiibox7yc4RwnzEqT+4oHbWKsuVTqULwFYug
lI8zG56uy5DcEnFzUXI4NX1QbW9+bNo0PhR77rs3ZrQ2m8oScvng+T/c/Q/xIWcc
mYXNO7GpwBzY5TelvODONrt4leLUZONOcgr3RgfJR85ipM7jUPSXbtzq9w5Jo2O7
+G3c3RDWY5v5hMtst19MNSXD7r+Kd6Jg7Y5g667Uo0xAD7+2EfWay0N50ut2FL7b
hJUXG9jSAQbR2cF4y3glTEhng4R7/FpFCR0Dm4Htlbm5tt18vaGzbv+KFXtM6ep8
lU1p+nPfx6///E23jt0AoMQaHhD6sxU2e1G7GV1d2Ei6uEUpQbiN9Dd8SUV7MfJh
lWM9nWlenf5rKqq4C9oZglfM9bQwe+ORm3QoAxJ7+906sWWkjRAbbNsNnVfUNHtt
umbjJiR+ny96FJnRxB1tZSTWCRpLX9Bwn6EZYAYd8dw2uFkO7ncA8u2ZDz3+KJ6y
KrxlIrHa06dwc54tB9PBGSdPk4XnY5pQs8aWsla2/uTLkJJMu8VX/Uqtp203XuWl
QIRP9wXoejNAaSEc4WlJGsI43Vu/GfoMFyG3aTsdkMV2Q5mybTZ/8QYiQRrd2kDf
gJjsYFIb1qelRG3FjdzDmckkPDOUcl3U5D+G+bNNH2rtyqztSm0HA3hxJkRZghlL
4CHjghoa/v3Kq9s5aWYqX5h4+SFlPsSjv+gE9HZryqnBmmpQnC/cmchsftamr8zb
au/lYel6wcyEhsjELg+pANv6InEkDb21cEPHQeyqdyxRP7++f4L4gIgwR8OxnYr0
DKJTQwNMIHRRB0/PP/dLo9joO5FzY5Am0qX/9p+gsy2aVjJYlAZyT86OPcjVH3Wo
sfL92hOvTKAi8v1aLFLMuDQ4vDcg2hMEbfUZ0Qw9XtyDhwy0dZK3DiOad1BaBdAl
QQiRgr8ZR8BS65QRyQGKm/qiL34YPSVed9HfDEgVAYSqleNsmKG1mOyv1jrbQFiP
tPeJf7VZ9w9pMkMBuRJrcpn+4OIZR8k8M0zZGOd+J6MnBDR/2hGe88R7nTWYxYgk
IjIA8hEGXDG89RwPLXpzN/Ziuu+B+yI6SnZLHr8gkziUbXBGjx49xMnLiANEOgc4
xlcNTifaE1Yz/4X9iaxbchd3JZupXVQG67KwzoVAwhRQobIcwJ5Udu9Lu9MHF0Dw
Sv79VdBqUklTWc0YMPPczdAM2nnP04hW8E+bOTnP05HdM06V2HkB+xWDbiN1LzF6
SySFllFul9n/Z9uS4Mb+8LYsobjsaTt6vu6sEcr8inX8YaEMLTI/23P16BZwKouX
JJJv2RqQ9q0ZOzoD9iZ4LxktKDhmrwaZP1oyqXv3LYZ8R9y86jComiDI4NJ8d0fg
KzA/Gkety+WavWvdzZkYKHedEBP9JVdRxdBEPbIuo0E1E+CH2J3rzKl4mlM0QoXg
Psz6hE+PE8E+/wtP9ZV4h7HmceVbsxDTb/ML+QgR0/80pIJ0fFqXzLpVfweYRdxI
/bez+S4rbi7/7EBJIkANcy78NJ/AwpY1npAezVqunWxtK3QnEAh1tjiorlM/WZbJ
anJV6QlGHDz/gEzqqypyBkr16NooUw5fz+xPPrKofNAL2wfJsWEQqLFunevcBA+M
MBliJWWXTw5BJxb0knvsBsG61NiPKP6YU6BOvH6lkcjr/MynoWD4IY3pdcoZrlnM
zsvMTeSiLYml21hRJ0289flfaxZIP2BCFL11GGFOH5j3qHgJSbqjng2aBBp4oEZn
nb4UisOFwarU5Z2s2QM/gIqxYxBO3bRt4J2TMp9kVpHKILHnKg7FeDWGROCNH+Bu
+HaEZrXyuvomSm5dSIqF27g5T+KOmEhllJ6b31PGSaUpL+5qjbcdVRmTs35celwc
QcaNhTZojn9igPN8yloyMPcPtOAL5WVl3DwU6VjrOVY8HvWB+sMQekDf2sQ9EVqC
Lp4O/RiCka2wEyUVP+Byx5k+nEi5T7YG8l26S93A8era9diHdvRti9JFn0PEmi0m
Y8lEicLDskd2c8GT+Hbh1uvXGUPsjjZkfU64NolZf87riK8A/itXsnLJMfN3QKOr
OA/fxtN+SH/uRvFYh0/WKgRm2MfnmbvKmVVtfnlkQh1eAfqlTbFeyTZv16e95k11
2C3WSizHZpysyLZ3sVvbCsCI+thrxbjX7Bt94dfC0VBPQp+oGMgnLupVCre607HC
Aq957QhJYRglePkycLgH7s8vUtBtdcJX45I04Qxnx3rbbZLPHVrA1wG9z49UMtoV
hN2A0c4rfWGDX536dDS4ZiaX1sA0EQOLbql3uEn8peOH7ZVlWafYHy1w+qe46y49
MVWt4C91iYUHQZJhkSf567odWYVPAqOjUiyeSn5wsldOIUDj9wf7zF9HYJaSyX09
yu8wfXmpVbzF0IqG7gNJvmuzI4yVAIsaP0uNjVYh64VXi5GhRzC/yPb4XJt/GKcf
1gt/Po5SQgVY28k+QVBUyUbtL2FGkwWiBpSm/VvGq2GwZ13wqYP9Ea5SgkJKmthq
/dLOHgXX3uk1T10+/QYAGL9KLC0Zg2iMv/J4ODHrR0z8PwT/UlIBGYwub2GHVbb5
hBbjCaK8s5TACF5tvtby65h29WmZKwUvG0icLijuozILE1dhQ67QP1c42j2UgYJ5
YSNAs/bYvMP45J1b/GtYDbLHfe/8Bwb1d+8vY4i5L6Xle5NsHRDSHvQ29F+Fm/GP
ATs0dhg3siapUIg6UUc3sZ0sDH26A46QNCXdujcPwdsGPOozoJ9mXaG9MrbcStKU
AetPjNDtfBFVrF1/05ghvhrW126KT5iSgaaQaiZY98mRkXNk1TaMYXMflChyhnd9
foJM6y4YXtoqKQyLLQdwZG6y4g5CASdtUK0Xfh6FwK7NiiVRXqUaRtQzmGiO5Fqt
WOgP/9C03WRKn33nGCSBMQKkws+fNRIW4L8Own30fATmaitiOqTyry6yBAiYmmXI
AGbt+s+XVY2NhLBQ4FiAAqKLgHp/6mNuotx2rAhq0cOdjM7N1FtTgzoX2eV7Mo2h
Wk4K664rZ2dVGzrC4KPyLqnK278/ETGquuEVGseS+C1fI6DceL1klbpuuumS82BW
hZcl40C8xDib2zNBTpbNEgnr5cLlTXk+5ixx0e6hgnJVJCukXEJ1YpL0rXlBg4c5
jA2uW6yY8jVMPaCxal0r9/BTV9BH0OWbqDMHkYcxckKuTF/T0IHvSJ3B7j4sHZBB
YW8YViwTAN+FkNcJojPN/n2TOer6NiK+0MD5cNZTExdYDmLLG/+ABFV3AtLuyg/B
H2LrlMdDo/6NCbzqV5ktwGKHv2X/CXD2dQbaKCrQUuWXDV9soBabSURtS2cpjgO8
gYu1QLy0v108FzsNslmKzuVT7KzkX+/kaDOGSi5tcq8UiuaFXtJWwJX574YfFjPC
m3PZmBJDz0w68KK85LXSnj8ihzF1LYeT08vJ83x/5bTalk1OssWaU/G5hMf7xE5C
k9Jzzp1f6kRgNwv1E6OzvUBeZ/VdqBxMRoax2/xXKHEx9BqMnEAojgziYuUCJYkn
T2EaBgfkDEC7v2NWuy9sY6PagOo/HXIDTdgJuveaVvoVdcv+4JmPXICpI3yElYue
psX3FhkR7FpdqZfUuZbQoLsAfav/c5WdO90G3jGyPn3UgC6l8MyA8Avva0WivnX7
qNFCq7M7EVXh+EYI3E5WD61CxIDktJLHme/YRVgFD3qme9lXTb77eTLw/Klw9A0k
PzZ5SgMaaDj7eXD5ujsMzJsrsPZlgsJW+HFQJCwAjW71f3ydsQtjLH+ZNWKcMpRd
aOs4UZGjf97NbVyEk9Uf6BGKGQMrvnjCjugTDJ/sFBAB6e6uNujzrNcdyWLmbi9Q
jFUcIRZN2eVJojdR4EwTzkasIVa6QtEkv//KkZgFqc0krW+UphUDKgc3xGNUcNRC
yCWZtHvxOrsS6QUaqj/n5qRq8d0Cs9Uwt70zFN+OQxt0NT+4SYSwz0Ojg1l0LfDi
pNhJRPNczJQoTDAY1m6tSHXjsw4oWGlBGGrmYjgoglmntkPVG/dHh1ZJBt31ZIuW
pCIsRZqGl60k7xKcuP8lMrFtq8WLpY8ImJnfFg8LiB7wIdgxddK+v6lnHoMG9DOb
s5bCI1cwKeraLkDv4EyCSs23DunUoPMnPMk2hmpdWpCl5yxDDrtJ4+OU+Fli3NTQ
NASaBq9ci789DrGtPXY/l6rn1TQR+3CmAGtgHQymV1Yzdm7Y8qxRjqtkQSN5fxB8
bnR5KLfVKnqFRZr++KcvUzsxM6Tl5ysVUBpTkR0tIwTsSE/62FGgcRhGAnC6F59i
2fi1F4dhnJ05PsuJGKTPYzvXxpTcJqn2l4ODGro/NT+gpITqVyMWJQqpkSaQVZCI
86SMk3FrYEiXs75YMO9cosRYCbYox6VHun/SUnXjSbsJ0BgjX5+qoZvazOKpze5+
FE5BaAdEZ/IOSb+YVbUFJF4yUtjyAFSYqStnAGFLt1l0I5n2LENnfCGZZLLI7nxm
NVchPONqTbmo6gKfCTJ4ymTDARYHh60bggPB8nHVfYGArJIeQ+XESa9LfuhE7coW
bA/j08CSHWmTJ7qW3sTu1vf9NMX9SyeWAB6XzLc7/FredjsCIG5j1dH3t8/fWWnE
OXIphkP7Vexl44I4jGDeG3cMp5JSBRnKEEYuG1IsTcyoF6QxyBDCVnB/BGBmdjFh
rOEJfR1Ukp/nDxTJNox2VCoHgLubkOYNq2FJjbM35xbTUrf+nwYF1k1RFy0yWYFl
lMiHiatMeNNKwXBwT9MOFul/U4fqN3Wxs2efBm4PbmowHRzwppgKFJuJ7mh9QMbf
6t1xvsxgJGx/s43GJWATYest1WX6ADZjPDljZOQNEynDUtr7dMcr2K8fBmb9iqJR
UtnshQAJatsdvfX2W1+mMf5H55Ro1JHe2N1xqKPrqnJQ38mXgMytV02CIYXSDB4F
XXEFmxjyYr6XLMr934wgFbJpS0IZSo89LAL+XSu/PUmRblwy+3T/hDrullwuqWJw
ZOKeAFoQ8YPVmQldFaEvEpBL5qhhgIm42qTbMCIQyBMEkeXSPoXRgMeNmt33daVK
MfSvyyqPSGyUoUM1LkGfOeET57x8b8Qw9r9ilkxF++XiftX9OK/eFi09zThKV5Fu
mZPDY1YEPY/vIVBa/+VGgsjlpuQbgCz9QGMY+EwdRNb8Y1aDTyMmMxcWgIvEMSyS
MzSeI+u5lnmCnPIXBeC5+dUc6SofW1JnSJQXOYfOfB2xKUno5NhSkX3gcnpi5D/G
r7VFOZHDLsn0dlORXzumnA2esJgTvHxCVm5/Od+JSIH6HizlbmoW5OmD7K/9Udq5
UtdtUleBr0MRLyx56B65s34aIEaZNqyjXl7dboOLbXMcxQWZ9bplemtk//VrxMEW
cYVcXUt5OenuoHLkHRMoKPOjkrg9qzWocuMPcuiJvgIN103cJjmBAfNXfG8NqO4e
WElNkRp3dR2cWT3PXDGp8SX2cXqE7XBv8y3+d9av+yZjagzYJuq4Wr4W/b/qln8U
nkMx8J/kpjWfWGZKOy+JmKvMSep7//a5ocCqW6HblqeXNKkRTIxCyzunbgr4/BAY
cgTU0rVZgpAOqmqhDLOfgj94qfFb7pn/cPS/bsQ2ZmBH8DLQkhSXddx0jSsdLlC0
XG+JfKwBd82+UHIegAc/ygAFqUiLLfzPgd8zGRgCqnoWOJo6gz2fxry1HS3H6Nun
08QcLbItvu+py0HVpE0uaR+kSD3fziXZR+TPL89uk/WnFQRugmBgXznl9oj8b7y3
OuJ36YYhUxgkXfmifPobqDGKB1IWDyFBhMnOJjiljVBAq0vJPhCgdF8rXY0RSfF5
TE6GcVij6KfpETNlMSIQMjI1gp7fGYfldc//O+l64duUJwrKxrIs2Xj07275a9RV
ujr5KxbZP1+a+5na5UmMQ+K+s47ghfyF87Gnlv9BYEseZQ433wUtocrlB9OnTp9c
Fsrv0fNcqzav17ldV3l0VuVUil+xapE0q45nAxUE5dhSWwg0Gsa5QC5+obTx8v3t
3H/ULLcmlFIcFI2p8eKboCPCcXXy2zPwjzevcWWHE4TtSpCY+ud4R1j3nCzCB99k
AGbAwHWskGt3wDZj9KH8IoipOtP3bJSmqcojlM3z45JNxI1esHt/qADv2ycj6GTp
8HfIzZnUIjUov/H9/H2PSEDC3orA6rir2iEJDATA5ZASnmxeZVnxZ3LinJeUh4Wu
QycpTeQQAre1c7h/+I0v59nO6PsvZ4AWHv+MIEUAH//+n5m8dxKuhvLrHDJwRRX7
yuUHukjEISsTDAFmOJ0eVmFrB7wINJ7VMFWohIFNR9T/P6ZVAv0YOwKI1RnmF4qN
0SiqVWGj5H+zCcN5YhdXr+OWCdFgLThXkpf+c/EfASk/CRCPIlcNXr1V34Plj3VC
OjdWt/ahTkDfz2lx9YBKAj1cTnK5ysHRtUOmGRUwK9hoDpEymMkUnSwDzl7b4JMr
dd+LekmSkupTZZRGPbnnoNIXU3uvQr/YyWmFhgeyoccmVxcPnevKHGAIv6dbQgr2
GkVJAthc7OLY3Dp8uxRrhuijxJEOxe7z7NbmDoF9R6IXzbrTPGle4UFlTFL1+Qq9
58AiW5fgKj1EVDxljGxxYoyBoTL85zUugRLb/fQ5y4IQYmPcifUClCu6n/j6hpvP
YepZ7o/IChyveqGlSnAZlfeoQHWzPq4LLFB6G8BUh6HLBsD0HLEshYCU5txPeNHh
13BR1SJzgL/2aBONZSJ9+g7GCTmMAoouxbKpPfutwwGMOCI4yOhJkqx6KM8GgwLv
lKWhi7SuknhBeyMngM7JZsYru+hNkVS5344YQsmSkCCUr1jYd9BzDLFo524gduIH
9SNj0xtvNxEkG/DS5E5Bgt35+7TR6H3oTMTTysphsAmgnIURpAy+nwztKHJSrRr7
9Vt/XQOo7/Nh/x/Pi4Frw0KTECuwjQQV9NWHGkefl0zzGTp+3QH9Ylk0jnpkGSVo
KQcPLKocpnOMNFA3cK7JiCJsyhKg1QdmxCMYNO4R3z6LJ6Xry6mMcj35IS/jQZYW
/l+ar2bpg3UkxjziB6RZVX5TXqAj7sQTtefejS1agvbFlhAAeXFsivz8LVFbjWPR
BWTdHc3+pNm15Kxy1PNbln032DpidGMDqQlQ7fM6dFGDRfr9OzeTXOiC2u9blgMN
6jgZuLz814KV6kp1nHwBajmb/ZYaUZnryYhj4rNkYqT/T26cUwJNivCs2PO/xkQw
iXTYerEHCbFiO5DlL1QkhLJLs/lk4w1itJWvS/6X0oXr9UREmHPvBsAFK6K4c7O6
+nTzLDg8FcCjKjqX4PwWlekyelefoelNrch4khXP42EDcEccuZMW3rGF4O0nLKEg
0cjJrD2QFW+jTCKIhRuPHW5/TEUeSaE/pOJs3sci78eLpVQU0rDxalbog985Cfo5
9fh9S5Xpowz8nX4a8o3riTBZepEv53R8SWnV8VbuizlA2tLeEnruZFWGVex/ViX3
ofeWfPOArBrnO4kkd1W4dQEE5XBSG45f8V2A0oQwvVWxonb22HDsy+SkvBVoItBn
1/sJG46rEtSKoOV/RDUq7LEbdctzq9S4++tvRJ1PVvFqQO8TEVCBon1+B7ilWZlz
eoYk/itB9EF7x1noqT3lQND9DfS/BTf5fVGY3uBfs+G6AL8T2Qq+I+rtmfXltt1b
2DyBtyb0P/zIMbfOEjiGwfqI95xiD1Atsv98apfE2/BwIR5bQ4HDDEHyQsbY/D8v
2Djw5dDhGZrtHebZuYWMwDckz0raGl939TD1Pg5E7smZmbEpeie8z6vdeUu6cveI
aib5vHZ9llHZsCxNn3QoPaGLF917nRYb/DrDLbHtyV3o16aMYkq5jvXHK/oBiGN9
UD5p1g+SHoVoUzTg+DDLjkcQx4BSD7wlX8qZbnicVyOs87YsjlGH1f4UerXXgGmk
RGX0uiE8xbVN7gGIYHynAcTKeCo6EI5GvbfV371dAD+RMqKl0J5OrPAnDmAAmmNT
OaoEky1Dpe7qr0glKDnGnLbnEO9Nwh5NfOV26Z/QtJcO2lLUZ8Rc/tdv1AplN8nQ
TdkvtDt9nCqZkDf0BxRDhxU1VMoEH0j0E2EnLwi4P/X/SdfZnNWcw2QtvrjMup/G
Dsu++R0Ylp33zf5220s3/jpu9ZNtXMyJSEeSRySkz9k9fE6TF5p1h2t+ceO1xveU
VwQwI314vjealt9GJlLBdbF9RUlGKCXqFMnm/TJNADBnGluP9wsofVS5fJqG0EPF
XSa2YV0cC1eLjHiplkZci8RhQrx74s+aZipKQPzEQ55dJ4VD3kf1CNQzdQLnzYjr
JA1psTEbSler7bSpgNPjAi8KYMfaBh4/oleOLROsR0+2QGp24WTiVlm0pd7d2CbS
iCIJLTmjJDn3iVx919A7lWjPXqq8n5w3nlWaADsph2D6Tk0v7eQsO+b1u6PQOlyR
36j4pEvgoALAzGttWxFQv5Dn2jBwkA2zVwNBcwUlXbunZMR5FDThDpoigHeYjbUH
PnZUVF+wKwhYd4XUEaZssNPc7QavGkpQSw0infEa41Q4hKtjkLc6NrzjydAvWmjo
VPf7sS+aXnLl6zQAcnwjfGNPOB68AwmjdXyfsGE58q94uEtw1TJVyRBdt6v4fh77
EezQuls4x5QgejJ511XY0YQveJ8eYy2G6+2Bl/R6FMXjy4sglIRyH2IisiBO8bUi
ydGhs7kKwtm0fKqmEJualJSrlfmD13HdknZ84Rhbna4qeHa9ME1blPeYShWxrKOC
Ot8rfgQoGDFiI4EAn3Z6TMPAZ0sr66nPopS06RZUGu3/aeUemOg8BDQTj02vYmUf
/Z7dlKRrnFzeyxBAKJ/+CGjFQCuRtowVrGd3tuv5Y56HhcGfWmqvT/U0uC8EzlzZ
EvYCm8R+NQKU856+dHXXOjzCSi4D9B2F0vxk4BVWcBFO69//1bcuuGz8+MQN/bwT
Ud4M7+qQVe+cT5DA+3nykyGZ/1g4rxochnk6ATFGwh/Hag0cPNKdbSJ41rjj6JLF
MTMH4HVCqN/cFmVkGqjVQE2OA3jQn1G38V0s+aHAQqw9kKsNfXPQSzAj97z7afpq
PIFGnSwvhFSdWhSjMklhk8LkKaNlZaVmDglUXhCmd0AQXAB1gxGnp9xyQfxxkZgO
/eQ2yM466VDT5gZbl72I25ljV0mGBTj3qGh3KNwHHgPBQg04BQ/M/0favhtky+/6
hLZ7K/FOFm1clmxL4sPk4B9RPGxVryDhVN4ZP4FPW6LGe094Cup57uP4y1cxEd9q
NqOjJAxLwqxxE/7rMrLZqhv05JN2/LHo/4cMkmk9t2su5MBMyaEJxzn+eVaxTise
2HZ0GhR5H8QVRRx3sG+WXRD0TCienWfVHLcKSgCnub0eVEVfvy442nTvCCQsurgg
vWESTOTVJxZnKc/sHgh+bMWOmNkS83VD2tLeKJMzLUEirzz3E/rDGEIS/1Rsy8u5
x/LFIXVYWAIMYOUqEJF7jRrObsCmOtB6z29ocyvIUSbO8r8alxsRs9L8ec8PLYeK
ZVE1dZO/Sb0Ltw4S0JvMxNITeDo5quAsbTG8ZMQa5ko+Bk74ewIgqKr59AWK0TS+
tEzq4VJvdFUJiHGAEa1adRiISPMLcrPzPUeotGcC1U7BB2XO9vZEO8uPQZM41i3F
trSCm59OsdOndFPvq3fuNzHvQfiofbmNrEwUmSQFP7eCJ/wLw9804SR9Bw9bqDIg
Qo4AdBWPNqbtlJC/GsQEc6fJrO6SQwGe1WRdSxBYnJJ0s25iLEpMGZ7XcDqniUzb
nzYZfzAtWAhTGzqjZrAt8hdqmJw8m6Cb7PYeB5ctctlTth97hDqSiD2Vo6hxLblo
rpOuY4VgTiWIDv8pvLBvx3WaJ2sDNT/Uji79a9+v1j+46lJD0rO/Cz6WfKYAfVsT
fhNc4TPANXX9v6h6p42KUBY0uhV31nl+g0GRkaLmLJYKSf3u6Q0rCnSsJQyjG4Tf
J7cMve1TkfdO28PSazbJhqsrnn7kdyHgj6bMFaPTQuY/CuZLWOoG4wO7aotK3Bd2
uBKrmhb9VNgIWS7IfzV3gIANlFQeeqlidhWW5MECnn6nDHG5uLD62iMZ6CwQRLWF
eVdMhc6GLR9lGXiZgv5bDnjMO3HJBWChjg/ldoOjFdwv2sPX30xV3QpArpMjaP6V
0w0FeKWmMkcVBNfLX0l6C8qjidRlIlh4CiqbmirqJACMwEgknUV4ETiBZ+fOTVJM
igMT33rwetDMHkrc3P0HvozTGjixL3mV+vDlKfiorgQciW5VkLPdwh/fG4fph2ks
Bir3HXueZFQGG2Koiym8H2AVxOePupfGUmp2+qcu/Oyuc/w9mnisw6wwJJLpVpZM
AAXjl2+o80qsV9QMtyf8ExivIZ3rO9ArhaJMnKc+Me1t1Xj5L+Vhl7fbd4/1bzDR
CixGlyd30FqZ22Oo8i/zbKYogqEoroqxpv2ueAgUStsY485GhI0DB1bUEvOs9XkJ
AqGfAZfFx+ZAcy5TXOrNi80+TQ+3DUU6dpXrNBANSigQfwWNeRYz8K0VMSnsSElp
+5g+7Ysj/pmvYpE8lkphCLqctaZgYvBsmVkwRLXLmFQABPM9D7AeB6MYmj1Jm6ZU
dVVcNFqSL8HjJMlQhy3BdNxTLb4D22hb8+vwN2H0KS5oNd3YBtPoblSxE6c0gfCZ
uJNHwhKxAw4u8SQEsQTju8Z/ZJu7V5c9OwHvvuketA0c5XAdi5X02yEr0FflE1Gz
L06UxdYKINQTE8wxZyzNIzrnIY6tl9Fmf7t5aTMJlRtcxJ0fVFvCMUzFLLS7wV9r
I1tleWpOv4Ro8ldd2ozPDX44dAWqAxIcncZXro2xVkxb76XRt8BaEoqeWYrjeetp
qamWISvjCbkuMTMFpjeNqGzvf1fP0rEeo/KWVtQ8gwdzlPvXcVoWPD/tKbkq9vm5
J14jZPvVRDigI+d+skf9KpAK1+g8NC0js0ConljiZGazspq7vIwyvBpTHhmbRLi/
vIwRX8LYcaPmWgWtf28HHrfBGQK6EzUx3Qr3TbRVWIkIMkGS33LllplBVW3PnGMm
VtAn5Plm57pk6doIZx3PG7os6MRuREkzXqsx1s5k6NanPD7Kc3H4/oXd2epOZGW3
sICV96S7tqCMFGhOcGmghDyCzloXNsR+evieZ+LtAmYWhty+vgIly8qqs3tIuBjt
6hRcsGx4zZbAiYTt8oRe+QaJ7wp/aPyzblLeoTIwQlrZgPISOgnBzXz5nYhWdbBw
Jz9Ts/IiqV3n6VjNI9K8dlbra3bXHCPkvhXh9vpcAXR5S/nWHrz5iPkoTdUJghNU
Yu+ZCVjLHOW4pePDO6Kln1i3h9cFTzVq9e5HIarchX4VPbJZnkfWLI6OA12MiNaA
Ww22+uBjg3+PNNGlcjYF/3MEJATTEPtarWTeXnrT9oWhlIun0MfKZiSnLfQXZ0At
OHOEQJV1WOmCpIzQkDLDMdBuuPzikp3Egb2dbjl1u8456M9AuXu7/thQ6v+ke1zZ
`pragma protect end_protected

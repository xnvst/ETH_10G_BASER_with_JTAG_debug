��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡j��-��l� �3Wʴ ��ȟs�/�\�Kڰ��n��T%�QjtD`�Z�YH7�-��;,z<�x�PY��7S����>)��fB���.i���[�;<�%��.��C��2���؁�eDxw���+Y����b(�OĖiƈ�֏Efsg�����n���>S�������Kx�"� ��q`t%�f��O�+<����=V������8�Z̄���W�����ӽ��M�b>�� �������
x�����e����Q�>���e/2 ��v]yH�)��A��
/����%Pq4��#Lv����Ms	�U�������?��w�ڮ�[�q��/,y} �I��(-���{���$�R�����y���0�!Z9;3�wS0ַ�P�K��� �6��YUg�4�$;��6#��4~KG!W0+B��+#սnQ�a}��s��0ǽNFh���CXJ��i���#��q A�p��e�{|4�<J3S�� ��R-�#Uz���T�����p��;U��}�C�c]Gv�9#��Z�~�^��UQ��!U���X�z��B�S�P&F�i@�v�M���n�+G E�]���X�������T��ė~�Ōu*v�ۍX�_@Z�dNn� *��ް�P^`*�D��a���1 ���9-'�8ng��
+��է]��E���\��̧};=�H�W�2�I:4~��f���\�G�̡�7`�@A�g��DO����|��p�|�>�֐�}����E�� ����Sg�$]���
K2�C�J�xh���{1����$nB�2���Z��n����>wm�^���"�Ko�r�Nj}in[DP�I��|�r��|�����}A�z�uQ �H�5s�'
n�H׾L�.�x�[J
���5(1���~��@����ΰu���� }��7�vh���S��G��R���p�b��- �zLM�`#�D0��:6���]@��-����iDG�����hx~q�)��+���2)쵗��nJ�\KL�H�z�#%�gs@3��u���oe���h<L!%;1z͑�]_j~������q�Y?�j�T�[��g�F��Z0M���r͒��3D�K���II2��I�::�!��ԭٜ���^�X`�Q�:<0c����>���ɻ�k�e�3ݧ����`�7����'��zd�*��&|S��C�gV�n��1�AV�E��:��	<���^���H���v�ԋJ��K��e,� �s�^�iXL�D�+�NQ�u 5n�uF�y�|qZj����H���Ǐ��b/��1+��q q ������k"��j7W �n���d#�������t���e
���j�u[܉�]x ��J^D���#��k�W�&�oN^�zxk�	��:he�?�X��)>������@{"�˭��H;����������90�@�F�y�U�9�m�N`)�~�j���le�AI+�o�X�2��g9�q�;Q��� xX�o� �����B��W���rߙC�ۼ�%D�4T3�)�;ad���_���lt��V�[u,>Xu�H�Q���N����NDR4s!r�� :<��^`��C�1��n���h<:
Ɋs)�=��<&��|�{�ȨYm6�?b�&В,�j8i��P����	֤�ʄv6�߆�_9��G�����*~w��C�o_�bB�8	Z,���1_D'�U��{�u��6
��������;%x�癑߾�
�ـq��ښ�V`ϣ��-oix@�.����6r��wm��@ ���4D���Q�+�<�i	P���%�O��Ғ�6v���G��d�%Y�s����>q��t�;����õ�}�8�@�&���=?��v��v�|&q+���Ɨ�D@�Y���f�B	,�3��vpHV=np7�SZ��5��Ȯ�uU���?v #�Y*�cc�Cx��3�"�2���g�#�Q'�� ]�µ���*I1Ǟ�HV*âZ���@,*Yo(`�����Q�V���`��?!�O}u�#��6*!f�p:m���Y�p �£�O5�Z=�.M|�[�(8�j��'����S���=���p���Tyt��	� ���3���p_�D��q5����A���P�xqV��7EG/�\�I-Q�EK9�ݽ.�Ԟ�٠��b� a�l��a4�{�\t����7v4C�v�08��do�2�F_�ofCHP�qD+mCh.r��F}]����
�E�%���Բr�n����������3u�T�z`�u-#̃���́�1ַ��6�)^�����9�@):Ӎ��5�`v�/��{��ӥ`C���\�6����o��z���̅[�5;­ypHe�d� ����3����G6��f������	����x��NE�t����
��ӔaV�_��Y�\H���dŋj�L��f�zw�#�����]R�ae�T�)M����8�:��Q����$dɃb�aKYՖ�8%2�I��F���9�֮fEb�n��G�H�%	Mn�m�9�'Ļ�����zGk"�� Bٺ�E��}�	g�xKH�:�
��L����#���]fm>2�@l��Ms���T�Ae��Ѭ��o-�T����u�����$�<lB�IS@���s��.! �r�B^�J�`R��4����`j,��a�tc����1�Ԕ��
��ݭ_���c(�����_��f6��{�	D�+{�ƆHJ1��O'��} 8Q����Cs��D����q0A��5���9�R�(Ȫ���T�&)�M]��zԯ0��K6�⚴�[=CM�ǻ�W"?�=q�v�����7�O�e���/u��X���#6Z����.�	qU=B��K.�	�x|cl�[��+���wfܱ��^�����y����?���;L�p�D�c� �Ai�[w~� �|�vU�9tB�7Hv@�� Z�F}>B�Pƕvq��0Z�8a���Y�`����Kd6u�B*�"�F�����b5R�Z�l�n23{�[M=�J0�rt�Pĥζ���eW�u�ٙE4�Y��j&y�5o��=8�xn;�	�(���� f��)�n���]I�-��Ct�.��~�	~Q*�`b���U\��|�S�L�!��>��3|��
�d�<�]O%פ�=[gR�{=�{ف�F�K����Ӹ@�qsŰ�>ŉ�H� Hq,�{�cX�N�r��m�sẈ����T���A��Q��}G�.�Ь�!#	I�i�|M���Wǋ��׸���j��	6�@=h�}+F�U��T�OU�����pֱ!�~B�~�1۱���Z�gM���,��b��M�A��4A��<B������qG\�����A�vu�S\�����z���b�o�0S�;�Hg���Y�ZR!'�8�(���678!mV�'��+���A��U$��O{��V�F�	Z~�GYn����w�$%x�+x��
��-�}F`�D����D�}�i5���f�����L�eU�託�V"�f�O��b*�)�&�R�+���$�O��Z�cs�(�ԥd ��ma ����X+ζYh<�dC��C�>z��k�H��O���_|]$��}�����&��`����|Kb��B�H��J̐��R���&OM/,���U�j�7`��Áڽ�I[?��qn��(ND�B���*3��ic�?I�c�kC��KI����?kG�g�&T�u��i���7}ʏY�Z1�
5{��toc�e���w����?%n�G��i�d��GW\v:Z"4����%������
=L�+o��jm��=��z�����֫�[��M4)��?�#9H۬d����S��Qa&)���M�8_ʑ�x-Y�"�A��_;e�*ʁ,�m	����f`�KF^�i"�t�M���CqJ��dh7�VX|�����b��gY�F>K�t!?3�6A�@�b?L�*�S��_�§n�Y2�#|p�4�%y��п�-Xw�	��~m���~0����h�MŜ��/��N%��ђ�p0ds�
�mр6��±�Rm3��^8�"EU�N��N'�=(�o��B�����>�@v7�ާMF\���0��m;o}*u9�t��.;x���C�W����|���9\���]���Z�|L�]
H����&��Z:��v���dw���c�뵓�	�E����/ci8��]���$@��ty�CSB��El<��Z]7\�`ܚ�O��$o�
�B�z����p2�����A���_`R&�:��'!^� �X�?�7�H�iA�#�AF�Ʒ<A�£�p��6ǻi)Ȁ�	�3�G�����1fK��$K�hQ�\�A�:FM�hm�B{vt�\�^`����o;��ߏ�D]tY �x�T�L��"���a�tޕ\�ur�$[�Sӛ���ПXQ2�q�蝝F�>a>k��Վ�\��?Nڧ��Z��;'�/\�-��%>�De2��Ⱦ�3�#2��t`�+;e�o�X�OU����ٝm�:J��Y4����y�)@ݘ�ܫk�EF���4��Q�.�#�H���b�EfF%�M�z<�N�!,�8���BcE��~�˺D889��I(?�I�t�n�|*�7[��33n�C22>�[4o�b���@O=� ���P_Ʀ�Z�A(�cؠ���*#A�U��v�����8t���TJRU�Nѽ��˴�9%}�,��7D;.����;�0�X��ʗ���f���$������MU�S��fL��<H�4���osɯ��*L���M`����sE��N�-t}I��8�Z��\,X��aH�r�RF[�+�x��3�
�n��@U���֑�*��8���7��~1���jT�����6�ՆaWKK$��Q:m���ɚiԏ��o�,���j~�D����3�qR�V�]�qbQsm/A�=��"f�Z��=��/��<�2r˕������WT'��[<�H�X&MP�;���땸]VY��(r�¥Ӱ����{z� ��0nc�Yt'd\{�-{�,[uj�8�;r�˲�� փEV�.;�������)��F��~z��J�Ø����'����ȣ����JvnY��r���$P+������wה���c�y�d64��H4����Ur@3L���!�X�I�M��!�y9G'-�D�6�2d�����͚� ��X�%����E�q ��ni���Q���Fn�����Xi�cSK|c�������=��e
vA�ǥ������P�D��,+1/��p��h��6s_�8`@!��o9���۳G��G�������BQC� �<*��So�<:��H�
��[Rq��>�Z��!)�,�,/��%@�6�YV�f�@�9�b,���I���o�Z����*B���Qu)xEUA�,:��9%a�زρ�}�^�ϩ�_�R���[#�,1nUx��N�&�~L�b���>��4��S���66G[��M���;��ݠ~~7U�U�Uk�Ƕ��M�,��P�������<UC����˪N��V�.�r�qh�?�;��J�)����]T�,疙��=_���z
9�2n��YmO# �0;�YJ���O��$<�GFu�v�}T>9�Sc��"yϯ�����[��KN��4yI¥�n{��c�	�9X+ K�>�aC�$�o�H>N\k	:����wu���"��!̯o���2Z��T��y�B.���LJ{^����f�l�os��"�Қ����������x{n��qv�+I�ɮ~���movx 
2.�豖�ht��%c7�q��t�٭�S��/w��r������7��k���_U��$�pN�z�:�S�f�Ul}����|�q�p��D/���#�������>���I����Y��;���W��]�;q7C_W)s-I�] йZ`{��C���G���*�X�����/m������tG~����<��bM�z����z�S�!��n���T�f��I8j��.��i*s'���x%�Ѩ���5� g�7��ɹDݯ��)����t%7<!<H�u|Q��m��~Ӹ�0��7$b�Q��[w��kk���L�3'��C!���	�I�����1��1F���I��6>�G�'lL�8 ��N�.�*^=�68B�x2�E�5��I/�DLL�'������_'C{�o&�@y��i6*oGp�A� �٨A�y�CY��Ȭ�9��O�G�4���Y%���X?�Y��1&�v~3f~�WX���%G��܇/��; ��=�*�ZH\�+��mA^C�/��)�ޔҢS�_��̬�%ڤC����g�6��1��(T��-W�Y__���ު}���?o��HS����w��ँ8���c{�J��K�-A���_�����B��2Y�U�xP�"����A�$��h����/M>q���A��	(4'��J�R����	Ѩm>��h�#��E�Q
%���RN��%sK(R�7���H	�-��G~�,N������B�Kj8wy-k��Vq,��BWܴ�8V�C���S�C��)C�Y��>Hz4-��_��V�E�T�Gb��i��!V9�*lx��9+�Mj�#++%;zJ�a:��^?�Ա���:7ˈ{&~����6]��v+����.�~o'���L�&i�GB�ݑ<��$Ю�g��� ���$��	�(��H��3��ʿṭiĘ��Wh��|�A�)rY�X�ކ��N*Ǵ�[ ��NJ^�=5���s��8�G�<���1T���w�ަx$'y�$p�m��A�N׸좆��dȄ03�n)�_h��}�������d]��-����˲f�z����	����F钭��	�vP2�_��I��i�Cγz��g�s�zl��:k"3�|�0R�9��Dh+�=:�X��3 �K������x�� ���qJ��hd�wGiaXӪ�s�3����Ga�ߖ�����}wL{��\d��f�4K�;,	�Փ_:�j����g�ӷ�Ÿ��-Y �-$�sR��q����0Y�2�*uA�>�y��]:� ielY��#C�K�� K:	)c�҄��DZo��-<^H�@_����%H�/�Ӕ{P�e+��G�Ÿ�H�d��*��\���t��5�<�m<��i����`��������iڅ�7.D�;�>���L�$ uh�!s~�9U.�����k̙ŘO���R/!s�CN�p��x/��+Yf& �<Tbڸo����l��D2J�5�4����5�		k�ǚ��&���E��7ِ��������O��$�q��㪞�-���ʺ  ����س���Jm���!����j{���\�Y��M����b3�/?B&]�93���Ē�n�u
S�Π�y������m�o�A"�Q(h!`2z�(��J�g{Z��yq���1��9|:!)IDv��Z��� �7J��mMŊ����z���<��j!�Xu����%#~W���̜T�p�_���7�@XYH?۩�z���x������m�d� B,4v㱭ئ���c��4hi�NeS�E��v[���/Z�N�G�0�呇�d&��|0,{��}�)�x֬ �褅
	q'm�%=Z�G3+�V�J&����N�5�hl�����n �7��b��N��t���@�q�Y%����PA�,�G�����Gw4�e�:
���ͯ�n#��T��+S9v�x�JZWB`�15� (ՇU����i~�C��K�-e�}��2��Q�z���"�����|� gxE�Hi�\w�:�b5��ͷI,�Q�p��V�x�����y�x��裧}!�䖇�FJWPd�A>����C�1�S$+�W!\�i��SU��KO���p�)"Tv�O+~)�c��]|�<�ם+i�K:mx�Ee�_�j�w��L18Zw��.*�]X;���?��RL����I�����H_O�YUt�U"�2���o׀�1.S�I���$rio�Pe%�o|�Z��O��������r�~1��n�����[��<uޥF�S��������B�%(=?�.]��i��`a��lZ�*�b��C���ڬ4wE�ٲ��!���)����J��I���8"�%@{�N�w&�:b^��I�|��;��HoCVIB�p����0�JY���S�[����+/��,J=��$��\�"j��I����Z�'�tIsuq�Tb�s�	�q,��g
p6�iTx�O0jjՐ�T��*U�;16|%�s��I7S"��o��A��/뮅p�����!�9$7�����a�����ZM�W�:]�5����Ɲ;�T�+{�����Qo\O��ۉ��-�Z�s��=���9�0�3Q�l�X��3O�|t�1V� ���݃��I$�ܱm$���~Fjt���S�Y�Wr}gD9(�tRê�) W��pb{蔙�A˩���:���8�R���K���JG����� �
i�yl������o�pfx�<�����E�<i�:Z�\��e�ъLo�����hʹOk7Ǥ�����Bt�l3u�$�'7�LB+� ǯ�>��G�1S[�em�������w���dGy/I����.܌k3�cO�I��Ӣ;��M�?�	i��$���?{�}�yt^����0��X��۳:]FQ�UC9T=���{��<;a_On�V}�p0���[��,B�"{�����H(�KƖ�/xAl��&/�E.\�Ƃ�R%��s��c�R�~�:%��ҬE��Ӗ�yHh�?���9U�ԯNݪ��k�5��X]�3R��������Y�L]�?ts�x b�R��L�[��y��9]�[�}˛�J�:��U� �/	<t��(�#�y�C1P�!8p;�����:��}_���Pu.q1�7�n^�
��q<�������'5���ˮ��Ӆe>�ZXX���i�����;�Z���u�"�������05{���֛g'Hܐ�H{�G� LM�"��r��z��5�Q�E��	;�}���J�`^��F�a��\�d'��f6�=7����?RjY�P�������������)���B�3~1�.]D$?�êf)��.��P%�4���d�"88	x�N�U����ȕ���q��
����K�5v�|�8@H����`?M���l�v|0�h>V6_��q�9��U�D�+I���q��ҬA�r��>
��p?���(h����n�R��>(�������4-��/�f�a
��_����Z�����|L��t���!�Wo����^?�}�����^e��tۃ���/l�vJ�U�[hX�	��3*ʀ=����uq���x=oۗ���n�bӍ�2R��%<b`L�
�*�?��q)�Di��j�\�H�:�5m�hdt����:��wD��v�D�u�!{���gǴD4�����SG����Z���b�STF�&n���}O�S��bM	�zfy��V���\��¼�����/0z$3�û1�ݥ/��/�P�^�����[��x�i�T��7�l|����w�@ɶr�Dba�{����r
�0{ǧ��W�O�N+5�(
79o��Z��ơs����I�"���lJ_�p� It�S�7e_ŝ����J
��k �p)dz*�����i�AH�7�}#3�fɚQ�i*pv\LR��᭔��+�>!H�9+=x*��/�u`�x�[[�e�,�Hю1\o�P�����e(?������u},���=��L��
Uw%��1��t9^|��V�1��0�-�6���k�u�7Ya�Y�R�Dȷ����,ƠbV���&������k�K�����G��|�!�n��W$���1�k������$�{1��Y�Q�Y+�M0�J��ٵ �󼈏[�bƽ�8�t�F��R��MM��+o�(-��L3Z�Ls�|f��W��`���併O��ĥ�"�O���-�����\D�Z���Av�m��@��7�&LpQ�V#��GNTx7s��pY�3߆���J�#ܡ�����xJ��X���B�\��2�$���K��	oG��kC�6*w���v�y;��*�z��S��'?1�w��:=S��$�(/Y9���8�g�\��0�'���]��vX�rO�Sb4��������G����j%~s��g�i�xǠfQR��G��h%xΟ.��`
B5v���v$"i%��I>���5EV��-m?�����[��ܝE�=� �W7��d�k����<��0������e:(a
^�շ�@�Iޗa|�@�P	4�7p�<��0��!<��/�|���0%�Q�U��<G �۱��*i�?��A�cܑ�O!����ӱ�R�Z捈��Ke��97����[|1�&���$h� �-߶,3��t2`�&j�+�eHh\�T���� [�����$WЕ8_�\�8��`	���y|
�U� �,{��Y�w&f>���&��^?�X������N�8|���)p9;�d�$�h�����`0@����! ��"tU��x�B�����?̴A$��� �~�Xd�Դ+�����4l�[(��U'��p u�,�bn\"��ƞ2̫0U�̂Og���Ǚ)�L���hץ�YC����q�!�d'<�^̵p��d� �x��p�P�b3ry]��^pF^ay6ݓ��+,e|��V��uq����36C�ͭ�!�@n�#!n%��\��U�S��4`H���W�n'��f�6�������r4e^�pպ�?_��y����H�K����6���C��&��H(.=�F(����?�Aq��w�!\�	���{x[[m�B��]im{�?.�J O��ǘ	|6�K�wo]��g�+�ɘ y��d_�
��`�����fK�\�f�"Q��`oNSwġ.@�TnO}}�`*�Kx,� p;�v�C�o'�dm ����||��WEn ��1n��|��pw���{��T�+�Օ�p�����2UkPZ�q3v���k�z�0g���o�qi`,��L�
hk�H�]�z��w�`��d�A�P�k5���Ķ�b>�i 5�} ��2�V�������� x�Y�Dl�L�h�����,��.�pL����o�v
G	��	NͿ��[�/o��>{ß;ؓ�,'�V{�i4@iE�����Gܗ���Nّ��IeӰT�AǏ�.����v:��O���u�B+PҘ�ro�S���U6l���c~�oQl�1'u?�]*[@[ų�y�{�Y��+C,pi��7>F���w8�1\����IP�+�����5������������� Y�VY���|+A�MZ�|�0Q�4�[��H%@������V��gA&(���D�R�4�ֹ�ƕ�g]m�?n�h��*�/	̻v�	��| ��i+x#�����Qz�A�,�fzr�`����l�C^��-s�0:�J��[y�M۩e`;��?M��;Mz䧨�ᕾ.���k��d��.T�aJro�lX�h}G��6���%!�*rif~��l"\��4 N�e{2���b��	aJ8��f�ܘK�R4�M�!�h ؊JYKf�=�'Y�m�(�OM�o']V�<<t���d&�t-E�`a{si�M�_��L����p���z�<�@��J3��^=6`ڵ��O���9�;!�-��}f�D|[�l�RH��f�Y� ?C,m��#Fg3 c�h���&����`��f��(��x6���J���Q��װL��=8  ����vy�k懮�t��ɕ�C��\��мL@�� �Hxx]@"^��r���޸C���d�7�֖3'�\fN�̀�m���8HT��d0b�R6��v��=�����r�b�Y��׹JGl�)��q#�����}�x�߷؃(���W�����~%�nn�$�l�狢��r/�b11���<���6X=�e XТ�bd���-�m' 6`� q��0�*PH��������ޒ���i��������o��lZ��G��1�CԔ��&%�Ռ�v@a���-���E�v��G6��Qֵ���bV)Rn��bhw�2xz<���WcY����8�#��'B.-����d��*!�F<h���t�I�Ѵ��k����
����L�'�I�2����	9��%!���"��]	�:�sAY�s�&�no)�Z���v0������D�[tk#c7�=�{��	*1�r;�M.�hS~ 5�qم��p\2;H$��ӻy!�~Z�+>��?ȴ��+ho��S[=�
�f*�\�״	���8F�y]�nWh��� ��X�WD	�c4����%t�_��#���׃�nV��y����|��1��֐iݪl����#��������������/J����/?	
�ߗ;�~�l�|�>�����@w"�q��
q�S��ns,����[c�
<(�޷*+0�Xov��䈖s
i��� �s4�N%��:M�f6oǽ�\qbkyv�-'�-��
rm���$��I�{� H �>@��i΢�>�� ӥ|���QZ
�'�2�4؈Q4���<�wk��R���M��a�nȕrc7E�]����d+G �OjO�X�+�Z���9|$�-��R�}g(�1q͜<@>�wCN���#nO̅d�^�L)jBl,>���*����sO�V5�]���/%'��`9���8>�ࢯ�~���͢�����]�p�o��I &��xË�!Ȟ��u�B����U�k��^�d��lX��UjKZ�v�}<���I�1z&�`Kz���H.0����[>��~��Poao��s5�X$�.-�î*Ph'������U?�
C��#X%�dvmMku(A�R��%�zU,�Tv�,`2[�͡*�U��`�N�V��R�:����fFbǷ��s6 ���H�Iz�5���wZ��K��]q�|����E�,� ��͔�D!���(���Z��d��\��������-t���9J���Ys�K�Ho:=Z��C�f��
�H+�9�r#O$>�:fLf{ C2�݆{��P�%kK��C�����tD�ʞ�8�`��=;�B9�z
u��L$V�=�kAR�c�"���p��j3�=�<!d�qA`Z.Ԉ��Sy�<�bS�$k��'�܁8'O�mc�y ���ݤ��G'0�.d��eG��՝�����(�zO��P�o�w��n�����a�gg�cJ���k7��d�ͽ_�٭8y0��@������uҶ�I��{?�uR��Kʺ<9zY����V5�8���,��.C*�6� f�ꉉ=Nޏx�8�Q�ȌSAY������& pX&�o*��	k�g�f��>���k�%���#��$�s���
�jj,,��G8��f(�H˒�F�↼�78��`'��sktx��S<��L����u��if��������ޡ��:�<��1 +�OC�:���i��_j_�F��|?����-=����� �]��:℘��*�$g��>��u+_!�o4�Xs�ŞD_	G�����-&�璗��q�1s�O�U-SOg�K���ql����H9A��bL�(����KG��3�iiEt�!Zq��O�oaƉ�Ǯ������2�T��ٗ��d���3\��$��G~&*�F���0�pFדh�,�,ڙtV?:"'�M���k\D0�D�yX��/b���'��L�O�Y�{��U��Z"[��]ގ�޷�P����N��ꗬ�U�)�:\�ܞ L���yHJ��m5}Nz��O�%��V�cl1"�q����G���e,�rF������j����؁Ld��7�H��>H�����}V�J��,ώ��Ap���ǥ�����=��k>�*�R�T!�f3�3+�ح�C���`m��ъ9�{���6����.Ȏ��=�w&3�>����:�`�iA؇�HMC%�IH�vĻb�o2�g�3.b�.��e�{_kt+QD��lRHr������l�eW��j]����^��� 5#���UL��GxM�k��7��N`���.X9�V.������H��M�}�-��\���n">����T>��
��7E�u^�p���_������7\�gr�����/E3y�,CGUnt+)B.�:��qS��}��_����8��'��p�U�`aM�]/��4֡޳�]:wwi"�at������:ec.��3���R~�l!ޖ����s�8�\�7h1�7;o���0�K���i׉�aM�'�� �)����K�n�u���
s.-���r��@t�;�\ڨW����js�I��J�sC��1�c{Sea�~��̉ǈKIr��Z�:�cAp�嗐-�Y���d>��Þ�U��`�@�u���G+L�
j��-�x��	�0�5\��*�n%�q�6������� ����=�ƬCvޗ��su����� 82s��4Dp?�^r�"u��j+R�c:)����*�+�����+��p��vI4ӹ,��m�n�2>,��}�ƾ#��M\8c�\�KAG�o�Ȇj�2�(ƺ{Y�"Xb�z42�d
~ܷ�scr�>(>�T�L�)]Go�WE�b1q�L�� �I���:p�*��{����El��,EH_HC0�Z�*�ߒv��]L�c��q��+���=[x�>g`S�HL�q��X��+ӛ3�U��5OP횪�s�s�v S�5�������=������0;l��/��
��D{�$a�N����&�V:3
pf�>�@�v�����Nm��4��n�ɃP�kU�%�P�3�8�(9x�Yi5�a#������������ >i�����ǂ6=۝���q������1�y����}pW�M�Y��\�q����C��8(,����ƴȵ��K/K�-}`3
tMc+�-8,c��Wvx2�0���d
���1Ζe���R�W�3����BZi�_��� s������S�)&���d��$�̈́�+n�A���.�J0�!�eM"N����3�x�����,U��J�G4��r�3�����5Áw\�;���_��T�i��%\T��t��M��g8��yo�JKU6V��o'�prT՞�����IU��M�8����;.�#^��0j���Z��`~��or�'Nm	���ۃ�-�`��Z1�||��R�������J�ՠ����EV��d�U�"�(	����S�����E>&��ZI����4<fV���� �v�o�+�z.y�Q���L$`�$��t^�%���:����
����j�4�Fϙ�tr^���hS��Îj�o��M��;&�ͮ	�EH���]���rv7�Kƀa@�3y��ڐ�,�{L�䪘 �t��������?[���ċy/�-�a�ӝ��ḅ y��rd�[����t�m.C����)�#<�3�,����a8������0�0�)��D�ɜ��Z����m���]�GۮJp1�'gj'ؘ7vY}��	L���������s׀�_��ٽ=l٩����p4�]���x/aB�ƥ�˚�̡�WׁD��Vh~�Ù$:2ȵ���3��>Q:���7 ��Ͱ���������Ķ��Ҳꘛ)z�R �
�<w���'���8��cf� 8鷆�>������t�	݋&�,-G��FSM{��,N��'��m�7�
�m��x�N*M��t��J���8��Y�	��[������������1�GҰ py��tɽ�x��[��}�"e}�K=A��کRZ�� M�v�\�O�ߖ�*t����u�7o6�ō�.���ֹ�� j]j��t?��x"do���wm��Bq�݆�ƴ��:)�+0k��-�כ��V��~�����y�"*������,o�/�~B�`�߶�EEb;��b�N�]�~��Ыߢܦ�N]��x�^Y����YC}I�03Cli
5T},m1������.t�?6�.��,���I0��dO�SZH�;�����:��\e
�G�Wޢ{.�p�T�<��Fޗ���[?7���p�E��q��-wx��|ο�;$K^[M7{dP=���<ss��Op�%KI�s�+B�9-Ia�u��./�t�y޸���*�pM'�$4�<}%wl�M�.E��y�V������!��e�/�3%�����+���n����m�o �b�^~����\-:����b�.�le0�����q��J	�<n�5mF�\��3W�"��s3�8m�Yq����z	���4X��, T署�E�q�+�h���xY����t�:Jz��]!SR%\)ٔ���,L�d%D�c�z�WR��pߤw��-[���7o),y,�|�ë���
dZ�N*I�f��dw��e�N-���o�Z���
�{҄�`�;S��4���#�ۏ!�*ȴQ�}/�Â�5��p���g�G���&����h!��K��D�)�F���}�G�ꍫ�"���R3��D�xk�~���?'`#>��GH�(Zp�CgI�YpZ��8Xr�,�̈́Ik���A7�/����<� %լ��I<���L�$B.M��^�����S�r�ahKW��c�M�:	Z�m�P @�U}�nUJ�/L�NjŰŏ3�3:��������u�ϋb��N�I�;{%Nk��W5���hٱ�Y2��N�a�����D�ǫh@kא�Q3
�\|��k�����B��hÀq��N^�d�dN�>��������6�ʳZq>`�x�@ƈ�}�)�Y�٪����s21;��M6Aw2�gK���6���b~#�8R�t�H��XX���_e����1��b�G��	���;�_T#��^&�*�|����D���=�]Tfk�rm�)�Ή���l���*�DŐ��*=�g��":r���θ~�����7T�s1}��R�H;���p��9b`��t�|�e/t���*68��ٮ8"%���=;wX\M7�׃���݆�� ���g()uRz��G�c�H�7�)�Y��xD#�Љ}�ˬ�x5�jЭ[�_9��GB�����n+���`�i�g�4}��ԤV�i���qr����v�P�ъ�[�_z:��$G!^|�Xd_���=���9k^!��_��]~��n���EOK����K,Of�A�ڵk�I���N��y���[�o�;�"��y+�]n{U^� V0��8c(D�˺9�%l�� .;X_�p��Л�-����)��8~�괷N�&%Qb��u���1��#��M�SJj� �L���6�M��(S*�gńR��X���'[i��qa������Vg
�=Z�{�8��I4W���Ŀ@�	�5��Ho�
Aٔ�I��a�Ta!a�>ld�/��b���KI.����x�N�eOV*4�=���aS-`��j�=����	Q����_����]�vlc&[�76�3�Я�|���X3M�/rQ�{\��}�u�RQ�Zs)]���>����*�w��:o��v^��W���(ުS��|� F)�I?��9�aJ�m8ES2��6Wm��̓*�<C8���JF��?fF�}��䉏5�9E6�U#��ٮ�>��:5���6 Uk���Xɰ�W(~��@CuKU!߂5������8X���k!4)�}��bU<�f�G֠��Iy��c���t	%}�V�㷧z=l�̑s���_T��7��)y��3Tq��Y+���,�� �'1�K�,�%�}ѓ����f�F�c�|�5�
���3�R-cd�ԍ58�$LO{x�Ob��9�p��a���O�>�K\ט�����*[�����,�� �o�''����c�i�QbU��}�I�l����A�,���|��B��/�<��<���0�[1�.�R({x�u"�t��c��*��(�IG��?��y�^���$ �<v�?�	����J� �����Fh��Ϯhc8䚺�1���F�WQƻ{��U,�r]����+"@M�V
{���8�����.1�둯{��:�!�bτq��iJ�ڈ��r���K�d�?����N�)�J2ܑ��_����G	�cfOCh 	-����͖��	��.�՘�i�P&��H�$���2᰽�3�Ѡ�.`:�y`��
cӥ�Č<��_�8������
����QQ��1U��]��){#���:$����lq*�:�8�����Ns�c��Y�P��儘�h�Q����(8�i�ӽg<�N���4a�Y�R�ꙹ��9��s�l)���ϔ��>[R������ɢH� �~�9��wպG�me<O�CT_f�r;�؆x��q���<'Զ[�:C���%�����=�EP~ǮKG�	&��A)��1��ǋr�����C� E�S7t��Or��\9�$/v�o�&�S��R�c6���=�ڣ�%C�e����J��B��&Ա�JGޓ'٢��������h1�(��d�@��I�}�#���1ߗ�u	�o��/8*�p~��ɮ��"��H�h�~�wsʍF�ţUϿ�~�,��ٍ@e���� �2�Y$����=��Q/����~�^��ڱpRJ�#�K2�NL��0mXC�g��JӸ�w|΀��¡�}:�����3��;���,�Q�.]�I*�B��y˗ ��|��5��Iv[�>P��IY-)����/�nh\�]����s��T$����TT�C��I�W7���E}Pڇ�@R����i�����j�.Lm�'+ҬCt(�!�}Q�mK7�l�(_�����&���*��0�#e �/51�6�E4��e��_�ej4f�q���b[/�e4�����a��VP-1�N�>��@�2�k;��=�a��Q��5�a�����8�'���`_�#�t����ހ�l�<�2�B��.%���.G���Qv³�z��^�w�<�fy��J�L>n���eܻVt:�2�~{ٷ�N���K�N�uSY��A�	��o��~�Bgdq���T���Ѕ�6roTX�qgsZ��/���`��;��ދy���u8aqF�����A'��bS�bm6�O�'�2E����Q��	���&੫��+4��ɒ���f�p�Ts&��4��Y%!ܝ�ց<�N�l0'Tm7XJ\�gn��1Ā�'���<��, iK�/��jR,?��D
*��<�B�Ϸf�i9��/�b'���q�c0	Ӥc����0Gur�u�;a���,�&)�w}Ssb9��'H����A�!X>@9�La�		u�Mjj�V�O�?�1��9q�0�3�s����˕��4���)�.�<+��d���������{�3�KK������5��ި�%R�#MhG�����mQ隌qx����䱃H��8B!�?�����n�����d�y�EȨS#Jg	K�ʆ���,�?���.��y)Bϡ�gZ�X�$A���#έ2	��{#T)9#���U��4�����-�J9�7�ϒ7�+V*o��(��"OS�y����wQ$��������g��(���il�,��O�C�	V���B^���K��9���}wd��
rZ�9P�;���Hl���^>�B9^�~�'�$_�B`��.wUm�֕����s*��w q�^�\M��*�:�o�	]w���˷�*M�2u��s�*X�2 $K�i跠���N@���e�@�E@�`ì~6�A��kL�Rk��n;#��}���:����<����t��;��7��8?-���U�;��
6�6*�Õϣ�)����..`�{j��\o[ LVF9ݛ��hx�r�{�<4]�4Q��^�^��VUP�_�����F�=p=�(��qt��x��]߃��Hf�T�e�i��!4�cZt�V�ͨu���7�f�Tħ�:�*���@��,�i����y��{�&��ɒ��%�:�W�p��8��IH}i��9���Y8�%<��+��º�((翺�����n]��c�ͮ�s��cR���O՜���^µd�N����d8�%S� ��5m������e0{�W�'ȡ2s���\�F�Vi<[���Ae
д���l`Z/�9 �9$�U��u`;�B��ŏ1V��#B���1���U�qs����o!/��WQUL��{�!�֍�2Z:�� �!�xͬ�/dB��+�]�s�5N�*e5�l)�����ą��iXj���4��Z.d�~��g�x,>���/V��U�8fB�'����A�f`;8!Jj��C�'.��-B������Oź-,�˚���o2����*M�����84,م�3V%��Rr�	�&61u��'�b�	���$��ͼF�{ �F�h�&,�c,�Q� ���ٺ
�|4򠇺"}X��Q+�v� �R��|5<¡���l�A7a� �E��z���O���f�t�vw�����n�$xb�S���������|�wSLJ�!����'rL�=XW���
��hɀ��k�M��֑��@aݐ�l�~7�w�{-�nO0(��KAV0FR�YH��̳ϱ�q O��[�Ax��»){��Y��?�]q�n56��ڕ@j�;v�u|���I���^ :��Z$��B
�b��BU�8J�nf�C{�uZPV\$�\��N�
/��d</�SI�<s�sx^��:��Ԙ�|� �) �b���x�t�H��c0ƀx����}��u�t�J4�LPc;�;�%��L�`����o#����F� va��'{b��s�r,�� i���Sf�R���E���^�Y��:#S�nA&3m���S�a��ݏ^M�	��0��5��Ô��yy�d$|��>h����f��yT��PkBSC��<,�~gVj�WB�������\h�scyT�[���uu�z��~.� �%rg��<QWN��}�&y�(o<ӄƫ���r'��V۵�����d�tiL�/��;vb���\@�H5*����Q�[�~rM<�G����!�v�����v���[�p\; �m��� #����/�QH#�T�y�};C)Y����/;!��ŗ	��GHDva0ܿ���_i��|^	�D�SV����.���P��/��A!����^�����D㢄ե�ǲ����N�HH�8-S�����N��-	ak��=��`��X��w�����c|���E��i��D�R��0���N�����*5;��È�y4��|�M#���=�1�1=Or*�Z2�6ߑ��i2{}�B`+���Ir��j�^�n԰�U�F-ٓ�u�脐 W�7��h��(7�M-��IIc�_�5g>±k�0�{��3g����(6��}�uXC� �H�2=Ӿ����Z�z+�1����iO��+�w��c�A��sKF�X�BJ�1��!�'1"�#�=�8���] �W�R`շ�"α�e��͟2C��>� ��b�[�a%����*.�Q@|����`n2k�ҽ8ѕ)�o�
	W7����:�]�u�>�SܐN��w��C��WCq����?K���_�	F�r�?T%q�w����})��a
�|�)J��8MjX-�� 3s���e�����A}��1���b�ӓ��|�-��ڼZ��#<egV���p�O.���������Ch0 aANV�
�	6ݲ�@8%8gQM��͘����_=�A������B쭖�9K��'���:�g�H>^?'��Ǚx�a�a��\]����	{e}�AK��Ȝh�/ &"h�1�ʢFә���:�D/�#t	�?/6��@rOX<\�RLU��M[�W�gɿG�w�{g҃�sO�T����AN�J&�v~������^":1����m-#�@�b�gy���8����,-ѹ�J̚�����dB�,� S,�P���:`s(�<��y�&	|��ͥX7bsd7V�\ܟ�nV��4�N��Y>dM�*��zTH���/�����_����x!�d���q�d��A	_(��\���2;67�X̏���ȝ�ֆnƈ�o~���>Ȳ�}�Ez���-��j����� ���DE�}7v�]u��e^F��;��	9S5��O���Zߊ߲�glxo�?"�F��p�)�����;�nlF	e��2i�>�4KQ�l,�k�����>�^o}^%�Ø?I,S�7 ��ʮ'i��O�
���S�J;+�-4H3��[�q�$�s&�X�3��Aӛ��D0e�.^�i��D�:�l�y��
ۯM4p�ޮY(wF����è��"5�LN-��'n�	��uP��6i�YNC�����aRU�68���W���c�;�L�����3@�[�'y�^)�u���F6���c��_*y�(�3�S�[׿�ߑ�0F{)�C]�lsz#_{6���6cd����m�Ó,A~����E�SF����"��]i@�]NN+C��.@( �a%�0c�T���a��V���Ȁ/���L�"\l�t֧i��y��]蓪6��n�G9G�Do�j�J����33(��)jD��.�F������U�AJG�X?�� ,Ĭ�A�~x�L:}N��' ������xU����e���D^s��T�������wJ���q��p�&u*v�vi����%��}6�����Ќ8P�g��k2�	��p�� kҖ
8ȩK/.�����o�8f�
�eY�{��c.�\�����<�|���F�W!���4�/�7?v�{C����yt�[�PR�%�����M�Ճ�A�pq 6鳱�"���B�~����� ���J�����']���I���`ym�ӑ��|s�-l�R��1��Au ��W�ഭ�]�#t�L�l0n.k����]�d�����;v!{�+'t8(��tg�3���6�W��E��F�Wo����=�"��v2 |9A��mH�hZ6$��=w���{�'d'\��:D��ϩ���_���
,9��X~d�Ɂ-�"[�Be������k�N0#��\鮂��˖�_7%e��2�͆���h��t���D�:�oH�:��M9Z@KiT��ݠR6(���X��hƮ��٘��B�S�y�ru���|�^����,����\v���{׭��w(V��,�)�k�-C%��d^`�$_Z�M�mC�ɛ��'�m���4|<Y}�Maiӄ��'e&�^���>��rv���  �p��*=r�28�<c�<l���q�:X7
�*k��4L�ON?�sB ��:y��I��ePW*r�]=�#���J�	�4�q�I��I�ډ��̢�k�)�@\����W2�c$�̲V���R}�`^���[	�+��L\��c'�ِ>Կ�Q�\�Hs6�e�7x2�sa�v+�,B�N��E�/�dBt���N<�J�MO �|!k�
_T�q��Gئ��W�It�Dol���5��
����T�sf
�z*j���Q�j���!��ŋ���%5��t���;�'�
�8�[���:'�("�k�� ^8R6��k�K���шRE�W��ۍ���o7(�u���b�Ԟ�#k�QFn�,�ɞ����ҷ'h� ��;�W$���� ښˤ�1�9A�c�4��><��m���$3�łP��˓$Y��/ *|�)����`�Og�=6�x�������;l����x)�P�����0� �mہ�}�`n����j��N6{�P��Ə~�Ƈ�~��Pؽp8�a�G�P��\�`�&��x�D��D��i��L%j:���o
��u<�8g�*����~{O�F�V|���n� ����>�`��
p&���!�{V3���d�ʫN޼�+��QT�I[�C���`lҦ�N�Y���V�g?)���D�b6�z����|&׻�}�>O3��
�۲w�е�b6�FkO�A����O���q�)�����S0�F�]�9-'���}K/�\/68�B���$�'Qτ��e�K	���I���ɛ�M��ͧБu�p�]��8"��:��P�b�.tp����g:AIr���u��+���������dUq�t��ڷ4�!�6A�	BT@+��, Iձ���u�t~�P.6'y�q��ؐ�K:bD�qY��Ns���F/�<�_M)O6��X�M@�|�t��Y��ؐ\ R���'��+�i%�J[R��7�������Yؽj�0��wT�E�������i<>�k��bӄ�ˎ��z;cڦ
Eڣ�?/	�>�A�u��%��}���:��(j1tsK�q�~|��W�������S5���#����2�ŖV�x�H�J!��5�s�n��O�I}Y7@V����ىR1�ȏƜo�c����s��xT���U��|��k�=�sO�B��ɩ<8�'[K���`!_�a���5��.��lʊ�\��*��{�7 ���&��Qé[���sT?�aؠ�YyLL�M��M]�v����"��(^�v�[8����q����o��]�]�.����L=��L����Z�1n��<y8�����ؔ�
}��߮E�� �ay|��)5�=`�?B|W�63`}í�Qc7L�S�w���H�>CG�kyï��_���P�ª�t��3��@Έ��(��
����+K��qcb_��������8p������S=�8��<=�ᗏ6M��_�k�C���q�S�ɶ������ 6����l��t�'��[M⿀�r����KMA[���	��h�]�fR���������=w�sC���l����4�Ѿs��&����^����*�Z_x2 [�J��K�%��~��ao��S�7{kfS�<y-�c��!�<��u&��O�Z����K���� �4����7ͅ�%�\1p�Kz�+�=K1���5ŕd}�fO^d����A(Jw��lZ�G���z��(��n��Z��Nr�Y��d�J�����~��?I1�gۓ�6r�k�a�OI�rO�X$�)��jP�ƅ�;�3	q2d����]g���/|����=)�̤�$��a�*�"�`�ϩ�f;;f��j:s ��:���wU-RV�̇�|fUț�& ̃ �a� }����!��\4^�0�cm�0�J�	@�ۡ����v����4���C���_������2^�e�c������WG�����*�gS)mNs�V,��Q�E�2چeef�R܍n�^Zh�[Kk��Yz4Q���m�#�X=b�g~tP��r�5��j���_Y��l�F	,���|��XU5�����p��+�]s�X��~�3'�yэV�Sg����ћGD�J�,w�vl���2{U@ҦE]�U�;#.�K�!�"8���j�%s=u�^���İ�Ɉ���3Y��"�A���>�^���f�g,Lmґrj�]k�xZ�0��������H�8O��Y���_i�$-Ђ�֑v ��%%u% ���f�0��&``��<�"��F�:���{��D4�m�E��/QC���x�� ;ջ�<���&�sE|���"�P�"�L�qj8P��&������6r��M�<$3��&����}��מ���o|��#x�W��:%����f��x���T�!J�%J���I�R���
��8�~v�%
cIȇ;G55��z�u�?Xd��kEkg'4����v���&b+BB��8~co�S榎�"��w'4�Pk��A�w�(��@G#z�֢������ׁ�I�����1VG��/�Ķ=�E>�C�:�1�V���:]e���Ѳ?��a��ff�֔�}I@�T'�sۉ�bމu��g٣X�5N;���-	*�Bf��S��"6�o�5���s�}B�%���?�|�9!�BJ�A���V�_�0DXe��h�$ǳ�3íF��>R���.���)Ui�k��@Y<�@ae�������g4���k]��^���>ʁ��l�O�����s�l�~9��`Xd������s��!�xڜ���z���Py>�ľ*�|_y��2!�Sh��*/�n%�tm���N�����4X���I�l)/�'�n��?xp��n��~@P�Vu'qBYز}iL�,;Nѿ�_M&1��7�hm�Ѻx2v�&Pst����xE�%:�ʖ������7���蚶�X�X޹��)�:<��΁��4��- 'Eb��m�cWL/ ^�K���7K PIs����_V�+��-�,�-�b���!k~r��KwBS")��9�:��go��L��#H��M�q�����J����H��,/�y.�k�~��ɑ�N�CAyh���ʉ�P�E_=�p�lÀ�$1MK}W!Jn�;�B�?��E4:��:�-*��3��� ���5����<���>�̴��E��&.S�~�>�\m��e(u��K��J8A�'7���0)*s��r2��N>�㴠$pt�����i�v�:ɸ2�A��U=�i8S��iWJ��l/8vP��%t��Ъf��ѐADLV��[��\�EoD\������[Y��,K��ϵoҸ亢@��٬��W��i�L! Uw߷�?��)�q�T����.�c`F#�r� ����P�����+��A��*\�K��$�.�j�y�W�*I`:o�`��
zpKޏ40�%�k��V��/��b8]y�����BŎ<K��1�%�X�pgc�=��c���X1��U���U&
^����GҪ@��>儗e4�:�x�X��C�&��\@;$}�����������d�f���a���-6E�-,xϑ�PG6#=,V���o1Ǎ��/s��[�����Hw*�]�Hg���jΪO:t؊2��wů�Շx�2�NAs�@N����K�q����T��?�?�\�1U����v�~q���P8����:��e���N�/���nkE�^ы������iq����\L�/�uu񡠚��U�����lI:ʧ,�F�p�n$���ۗJ�:ҽ+�*$�>��Μ�A�+NV��T@+������K2".���sLZ.tj��g��<�`2i׃�UW��+���/�r`��I�;�R�L%��<�c{���F��"��'��Wޛ��y�T����c�YhI�-�L��$�AO���J!������vR���A���^���=Hh�Y�J���~�)�G$N��=!�Kc�o�
X��t�`�_i~1Y�=���W��7pF��̢�� _f� ����8�l-p��q���ׅ3��T8�URt�������^��N��Y�W.V�1o��pLk��;hmY��Md�7.>�2b��}+Ğ��b���D��^(�� ��8"�~�tZ��j�%U�53\�3~���Rv��9q8��S�ʪZ��-�2*�0#�Fd�|�?�Y���eg,�]���_�e�s��p�>Κ��:�8ŕ�7w9�Y�y]EI��*�m�h�7n>	� ��sJ$I4��� 6�%�1 2tҔ,Ǵ���j'�7p!ܓ�g�; ̘�y`�z4�∢2�Lyi�W�*s^��=m��A�x���h9#��;���-��8Xn�k��͓
�w���J��S;
�-�o;TĤ?�jqZ�ŴԂ�/��L�]�盷��a�G��^ʬ�{��|yf�P�At�w�)Xx�\Y&�x��>�d�	BL���9H�)��ȡ�^�v�T��eS��#�V�=����_p��sn�)���Q�8�D��������n��0����#�����b=�j^
b&��vf��P^jq����H�C���E�qx�-����\�Ep�U7P���ˋ�ܓ�82ق����&�º��GAӊ�����{��F��LW�����r�x�1Fx�����0P�0kطz1v$Cn����M;4�S�1:�	z�bB�T"��& ��1�4.֬2�`L�0������2��N�P���W����{�S���5/�+�/�ը>�܁�%����O� ���Dܤ($mwL��\�BIp**�x��/� ��Q�dLF RA���"���=|��멯g����L՚i��w�$�<�P6�vL�͏��o�]��f����a�/#�Z�U����v �쮞HoN�R�Ŵ��"��#�<���_���Yg"��.�9���� �p�
C?'\�����Ϛ���u�H|�-U�R�u��T*��U�23T�A�����)E#Pk�D@b�*Ѻ��/ �P*��I��'�%�;�$�R�qҞ��ه�4�5�l��u����߯�5����5�*��߳�U��I`��o��v�g�Q_X"��j�pQsv���"�jxBx�vF����$ե�x%i}ݓ\?��]��z��3����6�<g{Р���v�����n��(�1C�*�G��,�n�<r�?�dq��Qt�6͊��&�����\�C��?����J�F�F�%Iy��ѧ]�lYVr&4�����/�\�0ec�5�(�"o�kb_�i��2H�U��uNf�=NpS�-�?�M��I;�G�}B��;al�_�?���BK�/��B������!�_�
>�j�i+�ǐb�e�s=V��,>M���
��ک�?Y��N��{��sv6�03��D�n%��8���F�ŚX�rL;U`������^
�Hꋜ;���g��'f��d	ru���H*���J�1�4vP�Te%�9��<�3��-����v�@0�tluJJ��#�F����<9>�)&gS�{'�
�)T�1�|V/���)<ld&�C!x�;Ɋ��M@�K�?�A)P%����Y��<�$~�7�[s;@�4ɬ�z�%���p�Je�Fe���H���7��Ƶ�����p��~\�����/B�Kg�����d|@lM-�:S[���r\����Z>�#?����km׀��.[ة�,�DڠC�[��W���\�/��+|�3�P�u�ۗDݶب5ᐊ|� �b�r
�4<$/{��F'K `i}Ρ-0J��Z�cg�������
 8ɇ�)'���*�������[{��_�KgC�N���h���ظ��e�{T4����w��f�x��_]�I��ag���r���9���W��K]�v�j�d�ה/����+8Ft�]Z���� �b�T>։��&�Jh����"����p��V���%s:s���SZU���͟��S#v��F#������i�U	u��hN^��8R���q-0�c9e�s���Q��X4��VB�B��f�?�M��Ùt�J���c������^R�<�̐U�<",��2�`�ӗz��BB� yS��5���y���ق=�dk_�q��7�mJp�v0�l2� �D�z]@ڡ��TK�@�-������hh��\�[�D��q\k7MJ��yux��<ې���u+�sa))��].�oT~�%�&HtZ�N��v*I�rJ�xq~�����D0�p)��:x|�>!a������Q�m�SN&��K�<�|\��o�[��QР�K:c��
��(���G>���Ƚ�pxg�+V�]6�l�q��LI�U)�a~Y�J�:n�Ÿ���E�A�?��/����ւ�M�HRy�E�G���F��G�ٶ%��	w���T�3-C���;8#Z���l�W`�
�]�D·��տW���W0�J��\�k��)���%�VB�W~�z�׫9�ѻ~}v��g$�"r�*�d���|
�\s�HY�}��Tl+󑄸�C�x���ǅ{ӿ�@Ynn�\Uԏt�"qE0��4�2yb �!��t2u�.��:q��C-�L)�Tx�K��m��NǨLli�\7�h�t�jM~?���F�y���L�3ǵBH$j�vXz��*_��+q�Q�P��[L}����M�3��Bp�6ѫ��^'�ٹ�cR؃U�������7A�!�����;_��l,����͍���"��B����;TOC|�x�7�F���C�I��6���_�����
��V0�I�J�.F4Xwx�|��e�dгE{�_(wn\���]h��"�ﭭ�g
�>I�Z̨[���Ǝ���n�C��J*�#���s�8r&{WDU�𕳔��|��D��y\�33���D+�޿I���/��Bjo]�5j�"�˫���|c���Pκ��+͛d����7t��j�R�X*��] '-�;�!q�>\�h�U�͜K8(��������cE��)3(��S�\>ՙ,f��SQp,k��-�2�������N*<�j?�6k|�M�H���x*H���Q�r	u%�,�$P��p$�`ww�݅@�"��6%�;����[&{�:�s��X�63��N&��>NN�(���51�hj�e���������K�\�QE�� �C�����ɱ��#t����>�s�)~�ڒ�۷��|�!*,AT��=��Y�3���+��o8�Ny&LT�z�i%�鹍�T-��E�r�5��R��ʑr�d�qāL�L�?�T[����� �����e9��GJ�j$'���O9������{1��χ9���1(*����z�^������_e~�J#"��@���~��+t��+hp<\R"����X��+I���ag�ziB��d[<T�ZE��xj:1=����C,O/#���(P�	"mB[�&>���U�p�o� :��],��A1�{���bQ2I��=g�v��+��%�8	�}j�_�eSŕ�������S-[
|�FV�Tʓ�\�M�v���>p ضZ�r���vDR������c���j����B���ܮo��̔��2a���]����(] ��/{sʬxjխ<�&LzI�S6�=�M:d���'>w_��&��_�������B�8 f��l�K�8��2x�l4�@oI��0�ńB��0FG��U�ʳYI��,�\��qD.���[AU��b������/���M���&?<#�1��$���8�4�����p�㻧������OUQ���@Z*Ֆ���m!:�Qs{%B�юS3|q���uId1���J-A��Z�t��}��m\��_��ov�a�a��]�� �%ݓK�Ң�mg����J�~��[;�h-���ѰM�u��G��iuo��ڂ� ��kMA�'ȸ;�im�Q�m.$O~��C�ռ|8y�a�`S�������R�����"��~��q��Ut}mk�&}�xJD�ؐ/�zEQ����5��P�BH:�/O���T�骫Q<�����L1e��$�^IV��j�6�X��jpO�6���:�!{F�ۊT�TPtqMZ~zVW���A�p�♴�� ��ir�#�(�[�T�M� PijU���}��5���i�s¢���4�6V�G���|��ɣ0��c"iT���'J?ò
�8��c���R�����ա�gCan�*�'��d�׌݌j^	
W�T�}�Ż�A��ӊ%ʗ=�;�Y估�Q��ԍe
�eL�ʕn��^m:�G_Y�c�r�,����t�F0�����Ҽh�۬EO��W�$q��1�b�/�)~�J(�n��"6$�I�g���� ���PG�4���P�8"���j����}���wH!������&�t�gq���Xb$T	a����i�X���__0��xI���Z�&���	V8���R��*�%����I
iR�:S����u������t�V�#���À�ޥ�h=��"���q�ny����9��ۏ9�������<<����^u:S��� F��;�_z��}.I��=�R?+�/����o �5�=>�	���V�Zju��+����QZ�vĜ�I+�.��
�A��7�q�Hw�Q�wB,kS2���%��/�2>c�kJ?}Tg#Y�ړm>}wɊ��-$>FO��H��������Un��ce���3���t�툳-��vN��$f�]���ً�� 
�b�
2��;�*DWci���:~�G[��)�O���E�n_w���7��đ�=����KH�~)�M&~=A�q�׵���x�����7��9��L��9���-vsɒz�V7�����\,�9!U�Tw� "�;u�Yrꭲۧr0����O�>�ѵ��AOS1�	�_��4y���@ �!����	��h[��2�u��>�VQE�.�騲V��ȟ��&L��oe�X��˗i�}W�����@\F����:�'�2~����R���W�����`)<���^�W�Ӕ2Z�a�i�Ug�u|��Xm65H��=?Y���������ۋ�oE[7l�����,y�{r��*�|Z�?b_�^e�	����%(D�֧���Jt��G��-�"����6����#=��#�ƫ?X�i��zv��R`��}�� �hG�����'|4���&aǜ���[$��
��L�;*@�����8��B���Q;�6ױ���U�4H
Z�����ϗ�r�}.�u�cl�2TԳW�t���8t1ЂC�ςE2N<҇���d�J@�:�Fu[0��[r�O�f��f�3�a�XlB�E�~qw�R�|��2���*ع�Ǌt{�]��O��Y*�ٯQ����k�]��Ʋ�6�˒�)ܒj�$��iQ��8h��S�ʐ�=�Ue���JCy�1ѩnd�&n�yp�B�N��n�|&Бb�
M Oۇ-�N#�3�\��Y���̠�JY���$���o�`+��R8Х��ӱ$`6�i���*�	v�t����x��ك����Z�e�-��՗1�u�;���?�)Ŀ��R�Q�r;_ʦ��븩�)	�6���C�^L7]o
fl��I�q%�H3&7�l�Nc�0�O��M��u��!=� �:�~|���a@���L����Q�6��ů�ߜ�����Vzy4c������p�E�]����)�_�#�5970�;
L�B�&Z#\�Ír)��Q�d�~�R�5�>K�A������ ��j]9�s�P��iiho.�ȼ���Ɋ��$e{I�B�Ԣ,A�z3�o3���`zzC��O�Ӷ�P��QayW*u{۹�Ί��>��l�%��9�4����	��ͳ��w(k+oĲߥq�n�L��A�H������b���jJ_���J|�)�[q
�t������N��t? L*�K�,L�_�P�з����U���qWI&� A�{���|6��U��2U�B�_��r��HY�5R�F2J����@�u��X�Bȶk��
`a�����h}�+�d��y�se�\�mN�O�_��w�5:+*52�ò�^bI`�_�amO�Ok|mc����9�;����q�o�{K��tO��Z#��5M(�K�?�l_ھ6�W<�ʜ�"�X �es����ɔ�ѯD-y�����h����-6v
a74S��n�N����q`U�g��8�Uө���b�H�n]���C� ��@�e7MM�����P - 39�3�O��Ƿ���<���`6�$�w
DP1�.�(�����_.� �����u]�e�RL����֪+!��m
���Q�=�RU�s!d�8�����\@I,��+&�|���eY�3kǕ3�([ѿX(%��<���e���L�KۥŲ3ԕ�m2J�)� ���x�QJ)�GW�8��9�"0���$�I_2!��,d��ml��dJ���t�0&b�.'tҔ1Np�D����iEj���oA8�f�6w�UQ��ub$���[��m�^a��X�c�a����U��7���5�Ԯ�w�vz��)Cᆐ�{JF)��ǪM�Y�J��F���ɚ'	�&�ǋ�%�vUMx/@���|���B�9ɺ�"��Ώj 9C|tgGP	��]�I�5�U��l�!���'}Gt�[�Y�?2�b�'IV��2W��dB�i��=�X�����e~�<7V��bе���X)��jM+�����;K�+j�B]Z���$�g��%�yʤ�.	�!'��	�s4��K�Gݦ�/O+e̘u�Pu%v]!C_6���|��G�2�Y�6��E��B�n�]{�2�Eֽ)�,�iu*����G�N�8ƶ�'0:��`
�fJ)ж@��MM����<^�Í]��W�����o	�{�Jk����AYP	}�<�Ə1":��*�L�U���7��k�����r�Q�0��-ƿR#�?��jp�]dʡ�&Ђp�tRS<�b` ����u8;	;~[��J���-��_��J�P�#�1�x�kz�N3��_����z��i�x��cv<5����!��Z34es��QI�.HB�C�2�� ;w�Cp���#�����=�D\���o�LR�cM6X�o @]km������m�W<��#�4Dd)~��������\c32�h�;��}2A���yrfsN8.��tt?(�X�܍��2�In���2�1�)i�I	�v3c�l�m����lPl���&��zF������=����N�ׂ�ȝ����_�7���F�vg�9�:��υ
<u��`�V�X�13\_���+\�����oDWV}�,�L��b�1G��T�:�z��F���}p���<͎�#p����&/�7Ss��=W� X$<�8�Åv~8����a�Hogը�|���ꭖ4q�P˰|o���`��ʄ���,�Z?�x�b�E��C�h�#˔HrK�[6�N\�?�X���}��V�F����ŧ<`�I���U� 5�Ox^t�ı��o���fl�:�ÙT-���v�����B�d�U�������/8~��T,Y���Mp؊�X/���q5������l���o�i�ol��=��wT��G������i��wO��O�RS��H��}`撚[1{C?kl�϶�$��p��9~9k@��i9}�)knG�2���5�^��#������Uד��W��R㣵+��^��7i^X�58�Dg���V�MĮH%�y������L������R���Ӡch��Ǝ��j�F�^y��wu+wV�f�4V��2*�RSUzT�����)�YNLn�&X���mL�E�ͪ���8�P2<�����~" ���I��lI�&�#�Ӭ�N�N����\���oAL@���r�^��e����	���p; %��G��T5�%z��x���r9�L!	��<�������s�fގ����?�A���梍�:g����d��Bc'�%uu#}�Վrz�R������Ŕ��ifbE��kw5z��{�@x����v�/��*��l�.��r|���!)�dԒ<��(^��3��������y%J� �c��Ղ? _���в{&&2��~2���D�B�1)ag�b/R�c�uH�*����6wʥ:8⦜��Z:aNCi��k6��@"���&���H��*�l�{�ا�0q,��$�KLMUL�Q`�M�󂞪�,��s��� ��m�uj�%Y�:�x6�炦���E��6!v��>!t*Ó�C�2g i,JzMݷ�� �2d�T�M��F��!����w��@P�g9J�^�n��̤�� �D�&RhK���q�;�=����[�d��mdo�x��	���M�j�M�W1λTp�6��z<c����	#��v��4�C3/���������z{�Ͳl�~�֤�Я��Sa�D��Bߠ�S�-�S�6��g?C5)~��>�@D���'��"�1OU)H[��A���ї���.���g��o����F�4P+��]C���;͚ �{<�s��Tw�H#��c68�c�=�aBf�q��1��2oW?�'��ﮝ�GN!2�7Fa�>F�J��E܍��!�=1E[y;�u��O#4u��R�7b85(%�r_�]��@� �B`����������|	U�y.�Sli/�Fl��Y�#����&@
�U{	X"��؜�����0�V.���ѕ�o�
�L�<�� G��8�3�~l��@8�Y�� k/�.A�(.3�q��n��:�,�o�=йV�j3��:��Qi�^i�e2N���#
���堄ͩ�E�M m���8��E��D�#DK�]w�D�/��h��!צ~'o/(�9R`�	1s}C�jp�ة��i�{�umYh�p��)�jK$�7\p��B��!@i�y����ꊠ������Ii�H=���{ʪ�I`�O�\)�p$؅���H4t�V}؇���%��x2��2�p�Z�65��_��\c	*k>��z��a8?����ʖnC"��Z��.��3��<h|�h�r�r9�B˝��ށ�����>_���5ً�_��9 �s�XJ�c�fme4�Mc��65cԙ+o:6bA��Z���y[e�u���˯ejQހ���cڧ"�͜��Ƞ!Ij�2z!���W$2[���9�?T�Ud�8��#�X��k^���YT{�5W1xe���+r��o�l��zuL=�k܍�95�����|���a�-ӱ�X�1���[������<�'Yx<1�m)���$���gZ��v�'�8n#�?a$4���-�q�{G,**qfnj1�.(�>(�����Eć���>�����~ݲ�G�Up��#�e��!leD%9x���Q83���3����q�9MXG�s���1�ԭ8̀�M�J���5B�/#> ~�s��sOC�|�I�SO�I��FJ.u4?�GC2��n�=V�_�����{� �q��Q�2(Ҷ�\�l��2Ϭ��/�
���b��)q��������f�8����k�1�Y'�ɒ�xx�dseTѫt�6��Ԗ���3�DQ���ʕ_f�����3�����M�+��G�����*��.l�
�������h�*f�����ti.|�0Χ���ؙ�93���x�7oU�Z��d���AQN��p��\�=�=�f[�x��T��h�GT���q *�uACvi�}�ˇ�y�/�H7�A�b�"b,��X�7ǂ���}l��ŕ�Qa>^��h�)�,4�P4OR-�[@�d�[��L��]��"�O �R�պ<����g�#�N bI�Kf�'%��ѫKa�`z�b	d<�V�� D�MB�������N
���>���I��3�9��˹����T�qX'���$��J��b�l��3u�Y��;��[�4w|v���A�(�mQ�m�ߢ�^�(���R����2��pm�����-`�Ϋ9w<ٔc�z���v>(���Z�>��A���l���#��gqI��-/1Lf�8�p�mlL�M'����tg�4Cc�Ӕ����w�n�YH<|=����N;�lBҫF�;����h�s���$Yd�m� F��+�&��sBc�
����X�r{��;������ϰw�tW]J(ٕE�ڵ��� ��l$����l-��Ox������l.z�)��)�!�'�q>�t�"F�9���f w�Ӫ]�#/�V���ܖ8v��q�/�e���"�䛟3�?Srkv黛oG� �,9h�U�fb[+���f�׶�'j�L��/(�a7�C���6k��,�	@�x�PH;'�|@S����������:e�{��5ebEd˯����csFB��5�u�]�J�o�n�Z��t�l�(�����m^�k5٫�ʯ9i�Z�Ť�쓧2��So'��ZD�}���n6kg�Y{FƴS��(^�
�vK�b�Z��
p9��3D�a�wXY�9�9�2M�������Ȥ2J3M6�PU.6��w�_�z��!�PA�����20~��ً����/|��(�-C�p��1���{�0�u��Y��*B˙g:={����,9^���,4���Ʃ+��O�A�D9�Z� �"�{C��*�*�u8�Z��G."�<�q�0�(f�1X�֞l��Z3H\y�ٍ�>��Ѷ�8�DB��ȯk�P��Y�&n�3��$�}w.���%����hjCL��E�0b�b��pP����藋���T�� ��F���n�f��/����XY�!e�qs��t2躹�^Q�8`�&�@�H�t�f��Dp��sW8��
����B	�N��I���m�hE�Ld�]d�xW�W��Q�q��[��XI�/��mƺL��格fm`�7������ϭ�
Q}�ի@̾�����O6�D�u)3�4k���+v��l��D�7��t/d�G<*��^$��_���n9ǛH3�R���P�UW�bx��<qC���Ѭ�p!(bT�t&-(h'��Um��^�� 'Ě�X���Z�l'<��a~g�p��p�6���x3Z�,u���=Fٝ��������
��PV�L�H�=��U�/�߂�$e8e�=�>C+=}(�[���s�
c#���s0&V%���Cш�����M)��~p^�(�%VE[��\��͏�9�� 1�4uĨG��j��M�����S�C^*�42���é-S���v���3n�o��X���"5�9j,��&�C��S�*G/�r;l�����?~D/v^��v��e���~F�����։����9�RNKx�w����Ֆ�rh�YD�!����J��A��7)�J�G��
��̗�M	����|S��Ά$pыV��/ܯ[!���7�[��ۂ7N�G�MR鶶ۯ��j��+��I��e''\il�gS�'~���v^`�_�����ۡ��<�6\�r��sp�i���*��4k�c�)���T)8�ۤX���ב��Լ�>� �T��d1�ȒE������
Gc������u���썯'��gC�w�X(��b���\�����i�c�	����6;��'�w�r�X��0�fM>׉��z�Q����d_}��J�Q�m*�T�2�X�L�z!�d5��8~�[���y.
z�7Ax�VC�G���_�*�ΐ������b����sp3k���ow��i���|3��i���^�e��t���r �V�k�_���i�����k(��X�Y��;�'M"�(�va�Q
!	� U���s�+Ǽ���,��>��18�5��c��*Q\��)c��v�/���m'�u�����?!���m��CtT`�p�^Q\��y_l�j<�����55|�鞥�-@y�ް��v�v��M�?N	[﹉��ļ1EZ��
^8��+�j/.���)p������v�%�k��� � ����cm|���g�!h@ʈ��;��G��)t���Rt&b:DPx���1��1S���(��6u�	Uh[b?�#\7�K�����k�{�sꅾ�œ���9|��~�Q����~�u��
��腭 �o�rȇ։�ےY���!�X��<�ܰ��9z�
�ڱwG�Xi���Bэ�~:�����Ӌ���������G�4���C����^�Ǒ6W���'����=
 ��]��9�ם�J*&�����Z��c7ۅ��l�WGJ��%d�ry�x;O��F[}�r�JO�9�(`,�t�e��Ji��y4̸͢zӸ^���a;�����O��T!�
"^�'	q��~fX�`�t���5ҵ̢���F��*â��ц �l�z�_��47U{}��g���*( y��ӄ�;L@cu�R9�DN��$��83�
cj��6�	�e�rSw���u��ܽ���ʈ��A{�r�b��,��b+Smjn��%v��l��SS򝤳�`ʿ�/$���eK�\eG���iZ�N��6p�h<���V4qo���>V���m��GP���[������\�J�g3a7���p��鮄�%Ԡ�\�!���)_"��;��7}4�M��iJrG>8���%xr����k�M������U��Qh�`с���l{w�E�x��>0a��ylu��V��9�Ǖ="���]4Kd�r	��;�"\'d���&. �_Y��W�����*g�D���|-��ȗ�mD�{�eP��8qM�������#ڑ���ʏRi���ˆb���x-���Vty*^`�g�|պ������@{�F�3�b����_����.<��
��~���K�^]���g���c���lH�2�P4��R����e���av��bq��X��:�Fʝ�C6}�f-O��C��0q��P�ր�<��kX:��Y�ա%�5^�3���`����wNVW��ApX�HW�͜6n�w��g[<�W�x~Z�|�V��C@�x��}&X	O[0#�V�_�
L
��k������n������?�u�����$t�D��@�+�»�v<������j�59���Va���Q���Ѷky
|Ĭ�ZjPF}B;����E��17+���p��k���M$���ά�	�ўv�
OB��7J%]���$�@�Vl`v")3�Y2:�g��.�Q8h� �
���xǛP�h�ϥw��T��;��ܘ��j�Ə̉�w���z�$��P�r��ߝ#,�/�{fS;���1��x�v`����d������k�0�U[%>S�bYZ$�fX���?��	2tW����i�x;{^^�k��x)� z5����Fh;bl��߸*��l��9������	5��B������n�TZ������䀚<�y�:��&f�0��r%c\�H����4E�(f�'�>�����l�A�d��P;�m�&��}0��ZI�����Z��Vt�G�W�E��FU{�/��{y���ˆ���iP)>D^�Ef<ְ���q�Ol#��y���� ���l�8���N���:��	Ǜ֓O��_��/jlLW���tp�|�,��f��	1�i���O�Q������Ȼ�,�Y�C�O���y�b���?^YasRp�^<��
��EI9��3��C1�}	�U����qD�0�4c�P��ӏ�56�~dW�l��u�|T���d�o�4aV�*)Gn���3)����=��|`ܧs��ZG2��d�i�Bm4e�Z���$�8y=�B%��+cqQ�ѩ�*��C@EVjF3ꕪ�\=�"�R�Q�uU�S_&8��j���i����c���2�sK���UD1t�@	?���%!=�Z"�G~*}�Ts'�1�"]��2)0�f�M�-�zg'ͤPj���p���?��Փ�6��a�^-�%�tw=	w��,�1�a�*$��ω��d���M�	v$��~YBi�lE�����D�#��i�޺��r/��F}�5,ޔob��Jw��F��J(�f��1�(�R��:H%���&�����+Ē�/��}��k�P���+n��@�uUg���Ȕ�C`O�^�h�wg0�|2P�2�]n��IK����(8v�/������[������3Hږ���,�ׇ���T&�D3Ju�.�F~?�p���Ӷ��5��"TA��F��C�����bsFn0g���69�n�B�2S��7L+RS9�_����0�w/P�v�8m���E�V�8T�-fs��f.��i,�W�S��}�vty�s^�z�Yf>�x�дR�w<s�N�bmYf�u����:N\�=uF@�7�����F�px�׫�-uR��\�=�;ڜ)^�e�F���3�Ħ��o%�t��-��WLI����>E�f�Q���9�l�)��
�+�����T8�.@�Z3%�)�iY�ؚa�l�墰嗀a��0�)�?�N:�B	ALx$y��@��,�g �0��6>��D��R�������1kѺ���^p��&�������`���佳�<�˘u�玿5F��W�M�/���^�2��{!�?�54YJS���l�#s�Hf�	���w^��m�9�{� y�(�E{�� �����5~Q���%�K;'7LW�~�s.~^P� ͍�h/1gpO���J�q�B|".8j�,��+B�!R��������E f�����F���Р\����~}�@�ٓ�ͮ#wk'�솳R�)�����S�'W��b�u��6�`6t���Uۦ=QG�0�=T���*�0���f���;E�>Gn��8K���/zsQ4���L�
�5R]Dvm�a_㜡 ���o��mi������j��T�ܧ��N�6!$"2/�!����c�װ1+؁-�a��������{H���\���4��=[�DzSh2��wοC<��8��7���Z�'���^&NaH���}�b�,,��6�eypl�-�a?K�2�A�S�8��az,��W&��6]��fA��ߓ�B� ��CԷe����1�DF�N����H�ɹ�*T >�w�`�~4f��$o���zAz:�t>�~�8�c?������ׄ�0!��s�s"Stg�no���m�|'z�)�5�!�O��7�Z9�j9Lt�����9�1h2�eaIg���V">A�( G�0�I���,�i��r9Y�^�r��Y�ׄ��-ʳ4��ja�鲉�
�C�m<MC��n��S^�D!2mW=8�e�c�A��%�U����5`�DHA/Β��DP���%�c��ָ��r���Mv2�K���:��ץ5��������ˠ�+��fl�ۈN���81��o����E`�6�R���*���;�u���I)�J,����NT'�����S"���R�"Rs���D}�#���^k�.qx�9�i�����	$o��Aꅚ����6�մ[VlQ9�54o�*J�A�NgTƲ���:^H\f�����3~�J�s��"�?���mB��r��95n��˨nP!r/�YMZ1�<�B����4�/�6�Z���Jk�a�x�1��>�x��=�2W�����2�y�����9�ೞ�-��k�X-�ς�ز�}�5�묣�A�J�]&�&�-R9T[g ��~SGYi��~�E!II�qF�K'�_���jL}�_K���Jk��	���C�M������!H��h�w}z�Cl����r��q�����
\�)��y��	,o��#��R-�Q���(o��s���k@��� R��PZ]�l�p��F�����+q4����筞�%c?�-b�>B�h[sҲ����J?x�\������]�|�}��@��أ�?�ٴ~�*��/���M���j�op�fS�o�~U:�����[V���d���8{͐5�zĊ-Ò
5rZӤ�L3rl�P�j�E�L@Q���O�穃{��*-)��'Q.��Z�X��S�~����%��@��H0t��`E���Q��O��6c���_�����jrs���妻�m��3����
 ��K|=2����M�ısĸ��r�`_�T�*�cWȘZ�H�=�V ��#�)�QL����]kJ���?XShw�L�����q@��	s��v.���F���	G���s��HVX>��� X�Y�|$���&�GaVE&�u�Y���6�@c��M�i�U:�����������@mvGY����}�`��Z'%�@@i}n�l�A�/m��o�N��o7��a���V��y��P�[z��34������Ⱥ$�0�BI6�Ɲ�X���v�ȉ���sr5��!�'ajL�fzb������ǓIވ�0RmC�&}��d�u�f��1?��֯��[=� �S�	b��i��$�bZ��A�`;�S���d(C��۠x����a�nEAS�g"�ct@����p-H(��|�6$̧Qa������Ԭ�j1��}���	a���Z��bf�mԄ���	��s��S��Hfko�'Y�1����78�̔��zn����dj����I�V]�l�Qp/��˷}���O���	�Q�]Д�yl?��,N� �m{<鹥$��{���j����	�CP�y��k�\�J�1�"�����h����e�Y!�<6g����-J��〟�<e�Ff4cY[4:�� �@:����Z���C�
0jy�qč�7��s��>d��0�ɰ�繊��)��"����&\�ʦw$T�k�2�lɦ�a���V9��R�Rn��u��Ix�"����:�aШ���u�F1D�;�C�S+D���:fx��j����B0u�L��(��IJ����2x���~��z?Ӂt��D%sͪg��`��`�vի�[UD�*.����\5�;��D@2�wD9I97��EXZ�!�m��]	!%r�a�0]�F������E�ۻr"�Wm�%�,��O2����񴒳���,���Yt{rB�I�,*~A���Z[����`�1�����L�������҄�͉��܉�n�$z6��Nu��bC�P%rR�XeM�~0$�:�K��P%�A��''yk����E
��6[��e%��_;iw>r��J�h����ӓ�PbȺ��\B�@O1�2������@�zcY��P�FȐen��o`*�16L}��0����9�R480�s�j�:�gG��x���y8���Q� ~T�Rv1$&�y�_�^U1	�;fc-n�Ļȇ��P�gU~u��-�ƨL�𶋌8��O	j+8�����"�3�cq��W�����b�*�M�>����G���J���d��{��1�U��b �s�=���+�bR�pW�W5+:���\N�v����V�P�ќ�Έ��[h��$%57�bX����k�X[z�;c>�Z��u䀢D"�@0�NVa�PL�s^�
I9�wn�W
��.���hܔ�F|���L�����{ޏː�*o<GU9���[ǀ�mr��;�4�cލ�3���bp�ڒ�������g��꫽�aO<�)�sd���;R# �<�ɗ3m^(1�x���|��B�*���k�8�Kɻ�������x��)Mޖ��-G3���U)jʆL4xuJX"a�Z���FT"����I�TRⲹ�&��gVA��p_����ɳ��^���a�>w�;kONT�βU� (�K�Mv�aa�0^r�+��N7J����O�������{>�nS���8\���*�@&*(��_�A�[-4s���^�{�~gn������l`<� ���I�
P����oR����<�;����^T]).�D�u��s.�B��	h�zE>(j?ck�]����I����Z%zj�,/~���w��.�K�E��~$t��c��I����`�+j#v���w"^�O����\�ϼǃ~�l�+䊟V��˛��,���W2����� EJn%�:sn{��R�f�.R6s*��=׵�|�����Z�����MWF���rSBn����4�����רH��\�E�@���NBdG=w��8��YyL�`����]���831ѐ,������mP'l���r��|^��oqC�5��:� �y�xdA����fw���` �H��4�������64�<�r�����0��F}.D�@!��\�r���B�������>��3(3u�j͏T&'�0����.��P�x	�X��C��̩�x�����J�\��窙�5���H��|"�*��8ҙSe%�u�\ȷTFF�xE��\9U-`z�YH���݌y2����*bzH�������z�}ʭ*u�9!��k���f`�³��^�6�W�bh�Ѕ u/��o��C�9�J�YE����J����.S�A�Щ,ɼ�L�4�9��c��%֦���a��}au&���Lw��pe�|׵:�?}�n�����m��)�����m	��.Z����S�C����#��I��>e�Q��j:�;�rcwz�ŒF��N�-�,�$��h3ԏ�vL�����Tɩ2'�o
%��+@(��r}^O4�:q|WV���I�Ê2%�^���H� �A�CX#ѭ�}���a���$�lQ
�a����uz��Ĭ^���M����LK�E=n䑪���^Y�<��oA%�"�ƶjK�IH%9�.-������	�A��>gG��G���E�"Z2/T`�U#w�qQ���q���7`JA0sd�������=!KŚ���o���;=UX�G |3� ��Z>������#�t��u׬3���45�p�\[�@��ڂ翧�Z�l��țx~qJ�n��a�˲�i�7���5���w}`�ܳ�ն������p�PM�̞"������M-��|��
4�+���l��$�����nliR0T�k�H�ø&��;R0�-�{(�r	���*�(b�绫��B;(��;�gyO�%c��f��/=+ ك^UHeL���C\��Pnp�9`~hq�kcV�R�l8Z�:1M_���e��|�#�]sx��t�:�&6�9�$�I�:��;�ڋ��+��b�i^�h��N_�I /�Oҝ��p��¯�op5X�Kcr)��+�z�~\�P�W�l!+j^�%s?{���\��P3�FAEjXI4h��}�l�)Zϩm@�b/��4C�j(F-p��&$Ie[�9@��� \4��,~&�*��m̼r���f�����~r������(h�a�Y��F�e����yޣ���I������v�k����yil�K
(��/�j����ߺ(iW��!�p���I[�jc��J@PD��:�PDT(t�f@V����b��Y��Y�(Ts��H�2t��bd���[:��9�&�8���lx�uQ���d4i잪�4���[+/��{S
fQ�/Q������W^6�/�8H�����_m�ge����WI���o�y�T�֎��+cg�Ѱ^{�/�p!v�@�#oM����MptK�N������
є�u�%gv����Y�}/����݇�l��/���@�<��@����[�l9�/�ԧ�����ώ)��t��XƔC�;g���R�ⲯ>=���Œ�����`���[��mxC�q�zV_&�!��5�RA�2\1�Y�g�QU�r��&!��t��)P*ʐc�5L�`G�c�+W.�_S]Vw�\6����U��� �H1΅{�b�G7Z!�PI�S_j���� ����k�]	�l�E��w/h�8ޮftq�Xs����[�>5e��N��W�7)���fF��.�//�ъWl1�$ڮH
Z�����E����q؋�X����EG5_�X�GAѨ53��.�Kظ�2�l��cdON9����%��LqY��AI���5¯]O����Ѓ
����cT��>��&�?l�fC�|��YsC̞+�J�'+�<s���^����H7JJ֝��R66N�mm:��k�|�F�AT
M�\��1t���YW��_�1��r��d��v2���c/J��H���ɭ��_%�3��k��7���/;B�T:c�����L���^�x��[^����B(
�M��ms��9�W=p�eVX���~��E������ x>�=�I/�t��yyu�4ЃP�*h�����,��&ɏ��W�)�0NM\�Ynr���⡦�k	2!��oD �(�'�ˮ��ј?�<<�`����	E�ޖW�^@����P�,�a�%�l�� �Ɠw�8g_��aYq�!�䰑��=�u
�Q]T�� 
�띳�rD��颶�W�mѶ*4��c,���m�u%�y���]��Fo�>����t��v��;��$��p���nKI�o��x���;p����B���
����'����1�6y��/��a*��|���)Y���Z�.b�Ć*��t�K}��ɟڎ���N�����h�eT�L"m��� ӗ�(d�� i�9=C}!n�*y�o�Ю�U�)
�Pe5�>�Z���1�fjT=�S��c�[��Q�DD�m��
@�To�1�� �}\�2KEO��i���cp!��Sjq��7d�|f��ψ���{1�����qU04���?CL;v��ӗX�c���EBo(]�*O�y����D�k�����B�m��ת�R�*gǤe$ע����&�I�Dr�����&���;�"�ԗY�� ��p8��=�(R�܊c�'�#�����k��R���s
]��{)���8�Ԫc�E�[&�-ǒ���,e��P:��)��4�"���p]��_B˂Dn�k���6_c��ڋF/�ʟ���r_q�g_������äKx=8���	@�\�OSVeA��,��
 ��`%=B��at��&	���"��n>�T�u`��vA�_LԐ����%L����W�*k�S�Mj̬��Ӻ�x5�~�_a�C7'
�vV C��r@ߕ n�۰���>��q��[�J�~�3��|J�D�0�Mz��G�o=9�>ǽ��"���6ȯ���ddAOÔ���I����P{��]��i�z:�����`~G� h���-�J��@nN�ޭ��1�	-�3�`E��B��������9�?DS�E�+��gq�1�2�ه�.R��@���=��\�þ�������R�n뚓��S��Y�rΦs��)��9sﺽ�3+�	�+u�ķR�)�׀���\��p�dd�c��~��/2���[
�bp�#��W:���d��?H��������	���]Ӧ�"�c!R���#���BAa�m�{�)LV�N'@�M�}��"�E�E#�6xd��6����8
�a�#��̜!����m��"OU�vTȰU �@\�� &l}��7�1��V�8D� c�.M�KWn��?�S�O#�U�4PTC"�=g��`Ŋ�������	]]��GD(͢2qܛv��w'��. �=�"m�;L^Ժ���C`|3!��=uk�,+��&�$����z���W�6I9�<���Rr�����p�;�=��˱�)��ǧ�0�b<yG�$0?�	6�O;�IT��[SR�4�2t��VM�]�NOh;�pg�n����e��I�h��_6<3��Hq^�v�Y.ɓ����֚�]��X��;�٬�;i�)~!v�B�nzE�.�����vA�;�#�?끌e�u���O��]+��+�X���8����.h7x���n �����b$����'>�COe+A�!\fk����5�q���uy2���e�KSD���[OA���3'�7��&�p݀p!��T�C1ˌ�'2��h�mZ��S��1�C����?ˤ��\��K�m��yqO�ì3���?��W��a��\�v���h<�XD�2V3%���X��I�Q������p*�Ƒ�v�;�f5$+1�i�~��R:D~o�?4vX�Pi�v��M��>��?~*��I=�t��5��M缠��X~����[���>�í5tby�7*�i�����b��'����&��&��i<��rēO���]��(1v�m!G��K��2x�����].uݡCd�k��͠RԾPj�M�D�G�_��1T8	���S_��r�A=��o��"�9Ċa-_�Ƥ)�K(�ޚ�L��cT��9�b9��������N�gKP#���՗�N��c7F�qŪ��f�̟Q��Ѱ����D>��(!.h҆�Hh�H�w�@TY�cN�/d@���h9�����G��P�:�O����G0v�=�g��4�u��ićV*�\L^+o"���&=Տ�X��5�قw +ֲ�.���YO^������\*hsp4����5��G�^>N��s	���
��l'����
~�`�Ƌ��L�� ��t�2���	�0֜Y5�ʕE��m�{��m�	of�)��R�ōG�"�tunګN����q���Nj������-�a�ȍ�k8��(�=�W��H��x)� W��#^]c�~��ի���L�,�H����=���l5�tG�,�+ks�t7�]�je1�W%�\==�s��&�G�!�u3����_q�l��L����v�.q����|o�q��4>Y��\���79g(%�����a���MF�7`�4����&C���A5J���Vc���8�ĭ	�?��E�,irA�����ڻZ�o3�������jw�Kǝ�6#?�Ң�C
�c�$�ͨo{��i�K���-h/}�C��8�^֫R�z��
|��_���qM��+���o�y=�g�%�i�P��}�'Ϻ�wM����Y�[��I�0�\���2�?\�R�Ӱ�}��(��,�-����<"݊�5��6=J����k*e��-ºO,�=0�	=����R�j����*�*O�~����}�˼���FBD͖�$6��2���Sj�����OI��"��Yk���A+V���q�p�J�rr�P��gL�j��d �':�u����ɉV����8BP�7�o|`�$�62�vN��\���騀R�=�p ���Q�d�6�� ?W5cn��~����%P���k@7�xv9��+3NY���N����$���|l�[�:�|�8l��n�����!��OW$��
��>YB����"�0a�0\Ł�@B�W�ı��G�TweG����%�F�ok�J
	��ɔ��1;^�e�O�1vNˉc���o��~uW|t�-������O��.0�>�!��X�$��V����B�|ۉ����6r����~K�|c1Q�ԃ��`��j�+GA�~�|�nr��{C�].s�հʭKQR0wvK��o���\�����Py��\�[
7Q�X'�=ً1�Y������ٹ���R@)-^����Q�<�0��7�fO�l�L�������]��E.W�s{Ư�+�)�H�X�(�B=6x�Vp���W�����o�ɱ;��x�&<�"���Z=���*�{��a�����@�ݷr,�H"������/��x}Q:GJ������Z��УW�e������^V�ɤ��1P)��|,;P\� � ���r<��*1�JpF��)��[� ���_�a�H������T�����6e�*9��3���HM62)����k�������HΟ%�zU�Fj;���,y1I�My�1�kVܲO���7������T �I�(S\��M����|I���z��>������u�u*�@J��ts[A0ߴ$��Uf���<9�m�;��k ����J�w���&~_�	��sذ��������~��`���鯴���ᎋa6��(��0��_E��_�:������o��� �!��or��
w޶o`)X����D ���7Nj?�� m`�(�.�/�!���r�j��W8������)Y��P^�d��-�r�E��� ����a��q�M�j���+X�r���H�'��;���)��f���� �JȤ|@�)E���\5��Y�R�ѭ7��T�T��m!�TD-��{+[y����ju~�D�.u�3����2Q+$(��eJ����H�Ms�	4:�Fݨ�����R|��G%�{�-�	J�e9�+k90����l>�i i@�1ǁ&��E��N0oM�Apud�_�o��������V��	�:�����v���U�
k��xT��.a�@���9�(�����6F�®E w?��髙XP*�i�u�3�����mˎ���72��{tY��d���\��=u���q�R���H���k- ijݘv�_^4م�ZF,J���Ѩ��6!n��zdK�2tl��p�фEKD�[��B��L�u�fr��$�4�]�(���c�xȔgs��ZU-t'݈挲�vP�I��'pȍ�Vݰ7� �1/��u �������;���x;��"O���^�P����Ou��*n)���G8�V��DjU̪�E\�$i�/��[����R�u���hWc�fݳ�E���ϴ�������K�T�"��d������0DV�4��!ՈCYٜtnz��h���"��`.]<j$����ׂq���3�X����8x�%���ԤG� ��&�y�mT.;	r��c��bC����ЉR��Yv��n�Ӧ^@%Ot���Kr~ߌ���{�$�����[ȗ��y�aN��^�@(���xג�h:�0^�xp��R�W���>�b��� ��T����A������gteGRݣ��ׯx�]�
uK�1.Ɇ���1^{�;3��.H�#>�2.��d��c�u

��pG��[���h�ktP�J�on��'����H�MI�$�O��������=C{���׫X��$'��
�4m�(�ds����JM⚳p_Gu[<��wĥg��D�͐ѱq[��u�c�.�}UJ	��C86P���#<$�k�=�tfdƱ�nG�h�X�W�����%�z��vn*_���a_���i ��t �5�	�QK�u��8PZ����}U:���i����V!r_p�:�U���X��
�D��r�!��h��Jd�:����d�U �^'1ѐwk�(�J��`��a�R	_��A;&��e�0���{9tI�,����N ��z;�x�yv�����I��ĕ���\�$�u�@�"�)�����ekýs��D�Z�p�}G3���>c[��)r�����;�!�kaf�F��.�2�I.?�f��C�n�;��q��-�]�3y�uƊ������Z�)�(��WQ8R��騧\O8T`_�ʛ�1���D&4��)���Ǹ[�a��2j�N���j�)*�4�_���2��+�G�B+����+�ʪ�Sę=���>�<���տ%}ޠw;ݶ�gp�3M�B� q�Altj
�͏}�����.n9�zva8�z�V9D�����'�?���=z����5����b��s.z8,����@Ɍs��~T��!?�1bn��;��� <��L��ٺ"f����@g�.3澞v�qAm��5�]�U;IF*�h!ӅOUc�m�����?�V�q1J�	M��z:����k��I�;����^��R�3����޻:��$a،&���^�?�04_{�*z�7F	չ���ZAmv�B�9��b�Hw����"� �!��k'�aX�a]��ܞM���Ra!C�s���2�uO�����;{��<���>�8�6�Sb1;k[V�:���C�>\�շ%��B��H�^�gA��7(��F�
�|s&��$���q|�q��:�W�f�F�uZ�]� ֟�̘�����ԧ�h����ɡ;j�G�Fм���KT�%�N1��l�s��ĳo6~.(LG�X�7����Ƅyv,�;�$h,�
�7V�n�:��;NF,�M`��h;`�զ�I+g�ɋ|��_�h�Zy�u��8�0����������~�N��o���- ��{^��=�;T�2͕�|��ͽ�n�2�&��R3�f-�>D��������%� }��
�]�ŷ�]�x��*κ�עzQ�'��z�Cj1�����5�x^~�	D*s�@͹�l0꙯;�j�"�����q��í���f3�R���J%2l`1�hGD�O�ݘ8�}E�fbc�n�[�$û���^�o3�>u�kX�5��f)���ݝ�2_�f�)z�aG�-�T��	�b+��9��'ڐ`/<�7���13ă�B@����@.cJ��}.�Q'_j�B�*�]0���1ǝ�ūԎ�eIꫥ��
&ގ�����ߢ$� L"���n���E�3�^R�M㬠��CU��O�[�5Ah3Ű�t����ۡ�����-�pd!ܼ9��.�h*�~�m�Nb@�@���\RB쫴���+����v!/\��S\�0���É!2�V$��l����޵V�Lh|�;Z��L��t�?�&6��]�VV\�U�OF�gq*���˛hޙK͜S2^S�8���6�D�kg\���y�k�*--�R��[�����^����c��j���m�A�%�+���L|הGL�"۫-6��Q|�`"��s�Zs�?��Q9R%���[t��:���(��Y�?H��&��2�pd�mFץ�Y��N���Z�ى�̨v�sF�M�x�4]����x��j����;E����G8��ȑT^��BQwr�4"Ö�ν�?�.]�����-�z� /�[TR�Q�W��!�Ț$�;{�}3�Wa�t��F��P�x��s8�ɢĸ��`:���P��]�ؒ�@�6�l$�Ƈ�E��V_��e���G��j���*��L7�/�E#�L�!-��	������4��#���$�橳e�y(&�o�฾�MȕK�M��s0���O��y��o�{n57��8��2���V��NZj�����@IMw7�k�`͂aI�	�mL%WU�ｺ"�U�i���gs���"_�����.
��X��M�"Ñ���'�l}�utR�\�I�ݿ���/��1���d�r��Կs�t����Yd��d6�g���>�[=ew�m�t�"0��u���|dYsU��*w��.����@Ao�4�=����p�oI�=�
ŗ:5�4C�+@�as1<R/'t�_z�@,����'rW죈WY>����l���X���`M1sS{�5dqÊ�	��Pl\�6i`�~e�����A�e���Ơ^��9KP���M	�C�!&����y���7������mq��c��yL�D�y�i��,/��t�w�D��}���T�8�Ĕ0����'�[
�T��nB�Vg�2�Ώ-�>�fc,�+X��!9�r��mc�Jk9tZ�C�k�>�5�b�,�ß'5��c��R΍�ֆ#19_���n2����������*�9뫳����J
h�e�/�/}�C �^������5�x��+�>��RD��&��d���gH��+�<�։V���*!u���r�q1j�e�ڭX�'*�T$��g}Y�*��b}�u�C�D�1�DI���d(�1獔,�+�/ބ���v�m�j���;��X�h� J|^��[ �U�G�#�mrǂ�i<?�C	(\0@�"��yH 0�I�ǷGm�1�<��ձ�)���@)��A3�&i&_��<�(�d�,�X�s�Z�U[4�צ0�{�M�7��̏CO���g-7&C����ǂnt}^r��ϱ<Gt��"J��Au^#�Ceu�w��w�p�S\7��ْ�ȜnJ����������F|�$g�T�iGQ�MK�-� Cf�ߢ�5��{J��1ʊ�n�i���9o���k����ױ�3�oI�J3c�%��x6����Ŕ5����I��%�@���u�Ⱨx��gw1졫D/޿P�)K��|?@#W#.�G��B��h?������`��9<^90��F���s����C[�O�8� -(,Ia���C?����,��(�aYNpJW�_���iY>�^H!�P0�#iO�j��s(�����+�J���n��$��%��R�E�"|��l�O����+����UggEGx�LE�JF��ˊ��K�^�&��G�'Y�F��Ô2�P�i���%p��5W��t��O.s�H'���j��|u2d){z6��@������m��Io�9`	�@�1�I@�MLq_/�U��
G�� bLPL�v����h^K\�������
ӓ�w���z$g$�vg��hK��nM-�Di|��-8��p�?�CuSZ���9��7TEp�����?" tp�mi�-�[[@��YyCn��q���e*� ^:��U�����ٶi5�,�Rr׌��ww��9��5���2}��OS�(����)Y�d���1��\7781�h�41^	�D_d}��X��Kf��+�u�;`~��v�t�OW�?�W� �%��,�x��<E������O���t�Cۙ����*^ o��%�*}���Ka��T��N����R�j���H�b��A6��W=Bh0�R�	�g�R߮[t���qo�!�#��$N-d�%ٖ۬�4?W��K�gK���˙�w
)vy���L:�ɦOx�0!�/���s�)}'w0<5�p�:m����Bx4/�T
�+n�.�����;
VCòF�$��hͽ�ڮiM��S�����{1�3D���?\D�����@��7z���t5����"��p�U�GMK���|��9��#�İx�eƢ�1�ކ!�/$�p��w�Ac�I6����'���8^4,�%�Q��gN�R\V��'A�\j]w!��{�٪���r/s�
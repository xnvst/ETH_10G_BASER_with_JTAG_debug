// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:24 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fDq+4oIf9SthGbrDl/jxLXqrBANEwB7llQVDCRwVunPBi26dkQ2VY5Ct2f8Hzi/u
eZcnfUz9HTiSIwGVyXsNJiWszxVBOaB/2BUt//BOMbTb7EfbRc7Dc2CbIR+7dTvM
eZHbnMCoGHllEN5zmsSavu6RqVD8cynquj/1kUdXsEA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35520)
dO7a4edv3wfILtm00nOodyrumnnS2dJa9jjiOCWAu+FjIOb4to/9e1KLFZ+w9WYG
Fz7+Xyf5PSfwx2nHJIYxKab+fIdDxQc62IMRziTOKFnEEmHFqJ7Ks89X1cXgOd2h
6o/ESQFONAnLuHjCSbp6cJ7N6VpGze16UKs+QLQb1BUWcCEcwiV9Lovv6hUW2lMA
xGdCO5x+snr64SyFEaZZZzhwQ26vzAWD2fwmdtWEROuT2uy5cfiUsYeHQ5xbTc7A
yCY77YdA67H63NrzcPhti2jNSQJllGgGcM5Xd0jSF2LyLZJk07ub7Z/CU/ajw52x
91UkDpSEWHVI42PlUkpyVqdOf3jxjOjaSbrpwB46ZZ2f+XgFp2RojV2I7/g8tm9E
P9qihNzmrJMdP5m5aQ6B/Hedgm8REOO0lenaapWj1S59tI4sSAmsc07eJoEPlJwo
gkaYp3rG6nIquaESdn3nDC0e54gkXQsczJCOhjYA+aWbmRzfsMh/c3+6aSGCXGhf
Mh/vbjJxHC7rQvXjbikTiuDwDQZL0QdRgY4NDbSeD0SgHWwlW6syIfboJcCHzIG3
7q6X0PDloBY6huLA746yZ8ztlC48dHNzz0HXPV+lR49dPGaHQtEHHlzcj7+aKulJ
dZJ2OizbMYp0XK8QKxAARNzAmcNkU6HbE3wFybLrfPifUkfWoXjJhC8/WMJ59h02
9ehBTElGN7Iv+CZot8dk1PthVEBkVg801D4AYroud9TO5d9dGzK8WQ9Fc1RYV4fR
nr9Clav0/oo7JzCnzU6WZ0Me7tQUo265lKj0gmNCh/BZYxMHFTUKW4fm2kzNQr8v
l8iWmXU37W/e6leK7o/RnaFp98GYQ9eXWqRaaFVWEN9weyUZdZqj8VO7e5rRBI8+
ZnjmoMPGOw84XIYd9SQJKAqf4ANLblVn2qZtJVgu+y0X8LeYyOaUxmeNMzEhuMCO
oACZk3ELlnKCS7HCOvbITTCFtMAohWRL83jVgkz1WwTR5JKxQRo8Beh8WGZBh8L9
tV8tb4KLeE7pu1ekgwEaKuwZodsr7dDtpW+V9QPcaFctq2CDI3cl/ZQym9g7xekY
WpLXL/464P8B5ODmhkkWrtIn3I/9kKJzWjpHxHNclRaoMdPv8NdpZ4a32H8a9wWw
CyDV8tczwAU4OWxBrUt72PVlWFIGk2ZwIUFtdhx1QkBZxMjapQBxs2qAYwOt9PB2
QxurLr8OcNiMF3rbuzykp1SZ88XuG9XfYwBWlCfxVgYrnYnwGEpyTmUR+GMYODM0
mH/m6xcvxIN1ywF6ahKL1JIlgHviE7YyzhOneXF7QHbRQlqBFb/IQe3riSSujnSg
lknSqQ4zJgas8g3gbkSkDLmYHHLHTjXFYz+mM4NtS6x3iwdWyw42w7lEOmD3CdQx
ljEoqpx/CduNNVA0rO8joOydKhXxqC1XIL3iku2Nb7K5pdlnVP+x4RtPWXNXpHXY
D+HURoAQxoOaE3Ly/yoxt+UoniZu2MipaIyli6Y7MbKunUsAyhEgOeVW0rhr/ESy
SzqreFRZU8fLKJLIFIvXo5AhxobaXRqAscooUeJmTD1WuwgtPxWsV19Ub9lDrY6a
0wXhZ5lEL+1r39OSinkLssmcZYi4KFcXVwxRAIUMyAxjYcXr8fXK1MTkNw7bWJCr
ItEHdGapJIwQwxtH+ZCq3EjpC+7v1OdfCwNulnBdy2kC4Sbsx+blTi4D37x5kJiJ
OSRnSrRQfFgB1CM/vEHo9VFWwmU1zAi83vYMdXeRXwjnr3h7LlcbrZa3vWviksRL
1RuyOe22VqOO8xGSxJHoFwTECmmtoo+dd5RkquzQ8RK2pmIMIbzSByKUDBAJSVLX
YhdPPJD6jY2Pihwr0LSkXTbyzXPTdhiXAzeGt4v71Rti1ZEn8RA6P04HXsu6VVEk
dkvyzh5S7vKhbeJNMFULbK704MyT2WFhJWRHZO4rWEaQfdxcLrfEyz2r61Rb4PLi
LBZwaGVUL7ewBNgE9kxPxk/qv1N9Zug/6YIzDn/mN5TAOqnhrfyqI05eo5aPs6lg
6eMdflL8GWk+Az9DePFHFcDJjIhyS4VEAeio+8/zQpWVzqEdZudccqjV24BIi3Wy
WjaCZoOqR9DI72hdZWd1dVSx6i2oqT+GvMKhxwnwUrQwT843YopVmKOLfVqa93Kx
o25jYwd28ZLA79nm5Z7ZhfKE35nEDqpLdhf5vm/i2wZSJEs9x7fSmd6KE5dtBnq6
wr1o6z0ECp0yTAbPMj7uZwypeaXgxgXkFezVJhuunnbUzF39mzn8JiWu3kILpPBs
Z6J4UmqqOB1O1wFSCEG4RROziM0u4CtDV+BjHvsHdosys+9GkyDWztMzxK6Wz3P9
PzKxPvrKO6JkSPBQXDHc49M+/V6S/4qBQhGxcOKyQDmen/eFXnrTz2ZR43W37WZw
SFyBErCF8d5W07up14TBpL9zTj/51XfFPW8YVBD2JH4Icc2YAwpmBYex2KeZsroi
xeSz7nSi0vrVr3HyHNmGTYkY+1eAGpVcGTVVlD+uiYrWNjDaStMgWvtwMlzpjyWt
1Cv4rPbU03Z6rWHIekA/5/ug7Fml0iD7/qTQJ16+amdAct/FQssGi2BR+bqj6zVv
FdwiK/j5vr6OzO5XsM56FaKwRohELNykw0vWC7YkOyux3XQVJVe4Uad0aCtPQEVG
eEye3tGdCwY2KvbzFMNS+wtx8Saw7YrE4doOdr/PGn/dYnAIk0QV/7tr6QEeGnfi
kZGdfIzQVzLTbsymb115T62ponYEXUmwiwG0nAYUVIfybZ0S91qHpe2PFG66+Es0
/qPWHfjpARwVbPafvlY5ka9DhnPE5EBgV1bII/E+kajddJMXc9ivfCyCKR+JbPX8
VZ1izlQTIdxmsvpdtI1BeLibEDbNjPVev0sotuCcfjbCB2UIK4NLmUH7gi2Ez5ZK
rB84Je6Q+sLKiNmWNlHsnH8uv8iqlu9l0xvRjr6ZSQ0rjRgd1nQcKHuCkQo8/y6b
nSke2ndrmCg4YU7+MGIZHJIwgEmDgBNtGatniVMqgCnfHCorVSYQdi2y677mDPWb
FDH3C43dqESXXNCVBYl35WcMVfSPnr7wbyuSau/7gBDsqw+03zqnTr38KajcIVAm
u0BUKNaYjvdtf2YTFisanjsVa+o11ahbiSAYZYYH7DwI+slWKLY5VDAJfliwMf4f
SXFLrjBonmknAnd45Ys+ak3HNBRBvHUqhvE76nC9EZmmzYykMysbP8PDNoOPUoKq
EtptzcM5FknLZ8DtSNJxgtFky8AgETs17t6RTuYWxbKmANFsZtyL5WNLkHyU+bCM
/8WITy6xKzOlYBwbAst3Efp72ngb913UiZNUiqL1nAUo/kJ7YHQcG6kfLjx+hBE6
KQezcm+mg4uVR4sw07BnZnWjK0wqpBJU4DxJmF4q3z0q+Q/mBUk70vMvEX8MUtLx
lMAMvAlApDirJf3snA1d2HwTyVNbagC1TpUoAkJ8HcnpV8LWgZOlgfJMMOQeppj7
elvlX4/6GoxPaD/WPCaPzin51i9Pv/aZMOyGf+fr5HOaLwluEXx1rLr0szon+lcr
iVo1ML4iL069Rk9fz1M/LyRgmFMv2Ehz1REYD8YOICMwauVrD32J/4TvmFXBHe4C
mRE34ZjDrg9FjjSmCWOpYV+/lmqaE/G/pej01XK63tkg5VFVZUUOJOzgzj2o+bK3
zDwLGsxy8KUPwyfEZofhr8ksELo+alrLbBHHbjKihIZZO3z77HbpwS/H0mVMGxEB
3EZwj0SLYjgS/GO41CTcIFFTi0NOM1oF7RObOq4rb5uH9oFUVtNobkLH5uOHrIF7
Rma52vztPdMwqc57JaTn2zDdaixB+64O/CiYdFn1BN1jj+u8oQTm3zZiurm833Dj
hglDaoh+mwWfgnfSmkFG/QLvVbpZXNoC0WoqAhU6h5J94N0hT6pSTO93NJ673Dqd
pQjgfFafkvuC8lyDoiNs8nw7pD9iy5e8Nklen7F6JSwzhVGWQf1WBpXIaBfM45/X
+OI+XMslOI6525iM42vBK/MyIOwZN5q72U1ydH4LQ8gw2pvMYg5VEsqrDHetRutC
QGEMROzq1ZXEZQNP3FxOWX/Pse0FtWn2SQiyMM4nFuoZiwkBDqd6mAmTt0wvdb1W
1qRGtmTw703wKrGnkYh7tt8hfUXghv+jSkq21eZSw+6Vq3OjH0H/jIpLK9QCmzyp
UO5piaUfSrLMaKlEcLrPqaq9KS3oP1+xrB8yIM0C7NHwoYLZk++FjL8yHizJWOcc
4+6bFCN6Znosu9TlKjccNYoNMsQ3r7Vze21E7ZACNseOVeEOKStUDqAGx9nKOTcg
IH9Ki0jwAsFqJ1cd+zlDk3ZOqthKVZsCBVk3UL2gQ3gM2FDWnJZpA/ZFTK6hDfFv
iSV1x9AGVHu0UDXUpIfuK3R984PwVi2ReTWcIPT+shXrnJIkNRhxKE+Nec9tSBp5
rHvldLS+4gR093xuNLruou4w2WVQ0pSXdSr90x+I4ehatrydIacSqwcTCNf2Tzx3
wTSBjKQW8ebhvm/XgEjC/VzER+L1ZEfbfa/Z90KxCz+m+BTx9hFlwS3K8p52oIRw
HTDxI0IfA1Wbour9F1KSSo4qc3DT9Rg6AJPIi2KtrkGZ9F/iSRKxLiSSlsld9JZo
ylBJdVUbfaw0u8rJHRLLAzFTSWylvayu6OlR73U8KKiN76V+dHl4hVlq0QrJWFpc
Aa13+1S6sXrRfCLWK/yK3oumI24evrH/2dDMR7JdN7GxDdU+z5rE65pzf2ER2O5u
pRtWnPdtm4ePuFdOrZiVmetz0WjjieZDV2Clx9FpeB6q+yiwHwW/uaJhMnEZbHIa
RutaAq8ZysQ7PfD3FXEI6NdUpN3crFKaAlVBnt9EXFl3boqHpUiFeJHZnUhCtJmP
ufaR7Dthe6Rnb1wk0XDjXa1MQYx0L+a/yhi684cVSQh6Tnq/8DKpATERZP7JoZ3h
LhkTRyOnrDUtoO8wEoEmFGDuMTpRa1HSbXv5unBzwhWbneGN9QQULF4+DZhBN4Rn
58n/DlyC0cL0ON/kIaYa5yIDerAIIszVfgjqJT9RUpJEtDkVwg0D0nVBEW5iNJLb
xwH+QEOwEVXSOIvoH+yVBxF1WYA7xQo0bk2HzSrfdMh7l5i+GjZfzIibwaBv7Dy+
T6RFJbM2k9camTS/M38rLdJn1GlnpwA54UYq5zh/8jooqxac1cTr5axZqc/Vco5B
Ve22fxXzMrNpLLxhCq1tRg0Ud9oibVHrDtC6oYkqHOkA+LpMmleCC0ahkkvcKynL
ZIIqLUtkoAuzVPOhm0RWeNk/LRf9QfWApI7cH7kpp918jWGtwRFsLq7+MdqA7HVL
7/Ec9a095lmB5mZSpZztGyjZ2VUboIeUB5QjGjOgIoBR4NOnJS6Vd3lai063+8e/
BPEDSMTQzjH1eEeFODujckBzaGLffAhaal7FVBDVkN7ehq1unWCdTK5oGeY7YfTE
Z6IFhLbpSL02r+zU9Nl8ZPnFgN9ZaehCClYeEd4fGshH8EMN/MlsXwHRtSEe/lxJ
2hzegTidXYPdcmKRApM3JcHSjGnAKTC7vHpn8z+Yc2i/iTWUw5bWCrHmfrQUkvFU
dP4/M3vBvmyNa04N0RYQm1PbEZ0ecq02/CixkaJmGkLxmUoy+kaAdHOFV32VNP3u
gcUNF4MxW1afu7tCjEQBEv1mXv909wdF+kPbGht+9VYh/2BCwSicXXwwv6tcDy4o
CPOkxvlXsZo9Fhz8Th02dRODEtW39ErD+jIguFKVlqGtlRXC+VIhUpoNLD+A1WBz
AEeS56OAWlyhXvBkKvyPwjqPgDwy4Bw6741kNjUW/wZR9hmZMFH9r4fHE+RlsH3X
RA81iL2sXsl2+xTIBXXWTnU338YXP1YhlJ55ZJ9trUJDsWKieyXV+IOGKUTWzzT+
sUOsGSEsRbJdta1sjJDfl1El+ayKFvQsi7D2Phn3BsZrMIOfWLTBHbNmVt3lCei/
Mx9pdZCkuelELFn0Cnq9oxPzCUjH7NYR/Qq2Jj51I3i0Nbsqji0a7nlFXahEPSGQ
GASPRHZtzny0lTvLnYHCnha0Z9exd9RmgYGY3uHRMiTZBaBqteq7puTSMYwmufoN
ySiCTapX02Fs49r+ilTiGmJ9Ytvv3xConNgRpkCPoEtGaTBjhnafeb5shQEewYHs
FUQHSRQLC8PhJD64RLKE20jyYDLAimNSs2IQ8gEfi7Q/14wKwFug/wqWzkeSHS6b
tR1gsGXgXMW4kv4l7V+VQtluejTf+D07OGfLPg2oeba84pbY7c6X6/i6Za2EnOll
t9UHUawt8hGQC5+xDwZ7YPdHlWrua3QIQV6bQhGwcvbhj+DV8COfurIh3zsdqcsg
BvO28t0sUdb1mpi0MYxeqzWZIVf6KsCDY1AxL6YjFu5R1zlmQzT8X1SwdKURvC2Z
k2jB5S78HU7r8Dbqhw893LkeDybSTs9Q/YRn3D1KX4ll4Vfe7/ZSvZpbfvXykEim
ssfS4j9NUKB+DdUP5+HBmJaymOIGZNevdZYZIBYkAtQpSvE++6ByCPsGQjQuD9ks
PJ+DM16FvjmyPO9D3PJiTGwPGprssYzv8FHqjxYjGyP4KQtYqElPBC+i9O2lueYY
ahnCNCDPNB7Yf7E5vL0T+Y8K25rwi52bZwJo1O0CBZcuULvlcAMn+S5VhK9OMuND
DRIwgWpHeRRJ7yXENEt4LoQeipgGr41UxsHjbMTwuq16pLsA/EdAUy/xot0dRTwt
5gC6svUYdc06onMKRRS++L/4yeTeQVQ7aVrPgXOxYP6/adgCBog32qH4mAowfTWW
jehlkH6IDcTDVhHSUsxy8JVRnt5kNd+xxFbRrw+N26JqYvMwe9JBthCyP6qQsWke
NVfmzbKrFY9JT/Jpl0MMpklY+x09mjRpDhZ9Ql9KOB/BarQCpT/1djro70mB8Uej
b1WyiC/1hbKXvJMUrCutrB0OYXGoqKY6rNjSGAVXsQCmUGDQbE+jBiemBmN+/+HB
VVWdKa3NDef915vQRPsr8vskn9PI0dyc92zwaHV8erKb9awBtvRLvAjr3y2wwRL/
UpTFYtxxpGr6jnNp2AxDgUjXZVRG+1UP9kbSECDGbfCoqEtqkh5S1YrrKFI0Va+S
IfKdiB/rA55ttSKBQ9QadJxZx+4YGrxflqqws+3Gu6J/M5mKI7JGyT7gzDh98bKj
6/M//eGE19Z+AYWYRYo3HQzYYy0v087z6ewZAfLcJqZBc3J3ul3y4e+Hv8HxQc0J
deqsVDP30VqZ2VQM3nJD9h4D9UmxM4fgfaqmikMI8Hd9zYGkzMpt10VoEj6NXHAD
oTjjsAaIu04DH01Vp85hfrmW8Gmeh7v7Aij2BhGB0s4B/l5eWmh3ho2G4DeQNnV3
O/60W8qMFXW1g8kOpR/dqm3xt4YMGEz0GqMfGel/wuxbZAvDE/4oo4joWuRUJo9M
MjKic/Mzr3c29cHUVjVuQzCUAIg7c+oAKrX10csCzZH8WWRP9qtwLx45H4LO+T2L
wKe43YM6DaM/9Wh3QKe65pJ5920oZwiQBkaHs6qBOjxbpjrNrE2B3bpJ+61kKIlQ
09FmQdrdHV/WaFMuxS5g44JciSAe5wB/a4/LLqPn6b3I3yU7EYSYETwBo7UlTyCy
2YUTNqvm+51gon7zIS8WiQO0bqeoZv2EWP63r/i86BA8EW7Q+XJygtwBz3POjln7
+XubzOzEvKMZLHatjFSUl1WvR/1Fx9/G7Af6RM33bDGVQGioCGkV1c2eku0ID6i0
DQhO6Fo1COEO1bc+kaliK3I0OrpvkjnAdky4gZ2wq4hbXtY9XWMVDajn+tVwPyrA
WSZDZBKf2hwsh7VnD7U/5MBR1CLlQDjxIaDDx070EmEaF4xlPKz2TyKmzPOlcdGH
S/+e7/OBGfKFlnq4nvwmTqeocOTyOgxyrOPcMGxeVrbLWWGPMbAiIpQjy+J6ACO1
PxZzZlrOG3CrK4NMcluXrIwtr3GSny/NpmOUA4Vx/ZnPGwiVjRm62JRjhzc3QkIQ
K2ZAVjOI6+c/zecd/s0LDpGOh0slbZIF2HneK/BhFv6laj80TsAu68XyMYh/FFnS
0dSdn/oSPBbgab8w8Qg9F9onNkeTU9di9sX6EBQgVIImAkDn0vq9Lx4NlAZjwOAH
rWBY3KY9SOcd444BIO77f+YjyOQObkWdwO9xUqXoHaAfs+cWoDWB955Lu0VeYAkt
KP1Kfdh5HDqcUACHDhUecV3IErBlN3ec1pZDzpb8rLPym1BKwE7rcfRqJLhCKsln
KhUkE/hoAW+CG609lCl771x0//rpcugY+dCX/rpQDnxypIXaPKuYDj2NWMAVS8mu
8B4iHBejiQwdZt0kYsMzv9lfqSACuBMS8NT8xfkEi7UJBfgnIMkan9hP1/uF+0eU
t/AmNewoiH4uzJEzp24JO+a6HTOcX4g4HdmUXemIwhI/AxVgCQL6ak/XKQ1YO145
vsCyf4fOi/U8XWrSmFxkxjLHc9zU6lp/sLq63BsDfyXaq4+uzZUbnj0bg8Q1IL3P
jLwHe92DyT4incYNFkgTZTBDNEad3orLJ06+utA8lEMrf8Bhqt8GZRGfVL/hax95
HmVn3zlbmaW3wCzzTkdpXBuzwxAj/ZeB8JYQP3H8zfbckKmSvWR2nqJx0lmbM4+L
qurxIo9IVrom9jeJ6aqkvdVzAOgLFp2IqRaykcVKKngVdJV/yUoYOK6sVg36XBIR
47CbqPwkUn8hPCDItfcu314y6wmyxpsDGgZ09hjL6Is2CSZONfbHvqnvS8ZLMmj7
scv/HmQK7BDIuMu4cuwSB5LhH8k+1WKhoYfdWZ3WPmnWTziGfvFrh0WpidQAmPuz
XQOoqz0VMO5rCKGE9f6ZYQEh5JMSEnniYpi74RrCd/ukz1sLFvNqnVaE/EWZRDoq
HK+y0HLVcLQqJv0RB0rsZ0qEmVOXv6/AiiTzsQOdWc38mVUxnOBTN5slxwjHDeQx
qZ92KpXNXGqcnHqmAiY0bta78Cu/ykFKvYtjhMnr4lPIuwbVY7gSlZEuU+lJR0Wy
5HV1DmJ/Il1ep0SWAUiDMMIp5JL34SEWwzVs84WV8Mbw8PL62gB6KXvZixch7xBg
T18Be32YtS9V3vkL98CJSbX6kWdP3Z07myAwzEYvVeVKFmZ55Lz3YD8PcXl5xb+a
s+Wa1PJAuF9R5EEQKllcXtZzj2zs8/6MjkaJn0sLGGL+4e+om6+5aEMKzz6JXp3p
hrqK9ETuNTaAL6S8ukoGDWxA973OXGFdpBrbU2XQME81WqqXktV0f91qcNxy/oqW
Ma0JKCIs/U8KBMDJhq2chMCEr/4HgNB3egOT4clRmTBFeyLCtstUZ1qs/uFW9IrW
rwEnC0WSuzXXTOf6Xf/h3XFKFghMiS5Ygvvt1uO9rKSD38g8my0oaAWibRc6e1H5
tHdR/ZGLwS3R3BvCvHmLny0zjSa0WwPPZDyh9HuSAUigcDmBYxnZFhByysWwPse8
COC6zRFnrjD716hHJru9PGw9v29y81+Qy8QzNyVqgFhWpDnT14ysmccRH4qnpnW0
itVe9o9h9wsJ8T5Em8cmCq4UA2Lioscds41oBw+OuY59gn2JyHHM0pTMr/qRgTJ8
YRvIT6CGE2/Wx80GkiNZMfjFIljMr/B7Lqt03aGLfarvMEyLw011lbO4wIReuhSs
mN4Ixzmrbwm1FC97dhCttCtiWtOLmAjNktXaXX+Bl+JHu0rRZNDt1rjyZkpn9Pql
kk8+q07j0UgLYGrSETlNGx2R2BoXBAogdIPkopuCoTB2ihBXex+N7UWtUInY6dpJ
cPx46pVA4ujVUO7M1Q82fW4ESN2r0RUjcjdL0oOC0qWPezeAYejLt15lOY1/DazD
qTsaVmoQbwZQJ+P4SMZhniErzIaTtQH040h0bXXirDz63q828utJFiXOT5788EUi
ID866W/7llqFfCVoc3Y4YvYNSPI7eooeKUtqqWQdieRGT5GnYAowODRX0wp63tWd
J7OtjaCqAXFuQoGuIOT3r0UTo5NODAotFCdwjnv6JfrPPidypt8TPZIL/QZvSUV1
TudNBo6YI2Fn/5pALdkXPMexse+jwUCqpWscjNdt2o93lbe4thPR3z6d7psfzdeD
21AvJu1x1Mmg4fMFhDA4kVdm0RQPEpLllu77LP+nTRsp293go265ZiG3EA5Pf9r/
eg5tw/KgXgz42zeyuNSOoCgvhxKllfk7l1PuPIIYfmdX9Gkm+MD5dLxqogdlGbOg
sxxd0L0vhaKXazS24nZpvfOXcexPM2K43oZ6zuOZUo5Ddwgnh5ViMT3RzLIo+I9z
KJbJprbJhCT0b2Gxv0iqmeOAr+fNIe0Di3ygLuZBH9DP1ee/NG4iovbbUn1ksuaO
0h0YH6y/r3NXTD9EJd/g+wPq1Y+nu+nBH4L41B8m+17tSNlHhX5fx8cP91ExnKyA
WJ4Qzv6raGcNxrqpeBhENaMVssr928ypG/4iLQuq1we9SgdXsC6IY/dCEqnQr8eT
s91e047yCdjzCH9ltfoMW7O05wHlE2jFBPG0fJER40I6L5AeOEstopFyQXPgZT1g
Co0s/9unt02F6UQwGUQGtS9yCYYNkaz+D0T6errcDxrkQUbpIrIxBB2Vlg1wky4L
TmL07DYBe292cbsrabRcAZUOX6ceZ7dzZj0xQJ9CVtk4DYjRffU7GdJunwlnWb9I
JK3GAaO8/vOoNLuvhP49Hq03ecsCtFToJzVnfXfKCVHiEau5kKmYbss4kUsfOPkn
znKsNJOETc6vGIluiyVUbcCRa8XHDjblfBiG7fkbIBuBAibm1Rlox9BngSRGH+OE
x0o4eS/1/Y4jyNdO1mpktv6VntYfSs3UIsgM+gFce0jenfM0Sdux1n20HD0/+9gY
uv7mDlo/gDbRkT8A+VxDaeAA/TkNgNJdFD42jbWtgvcvORwtniERZ/Sz6GY4QNAd
CJ87W8Lxuyon65Dh9e5mvvaFiZb/i3DDgsjpSAcrdOzH+3omKC5qR39pXUxnV6ww
pRZZlNybHNLpZ4bg3Kw9Z3aNt4rkYpmSvYebx19t9umYWVqN/UuykSbnvA2jAWMB
nzP5Df+E0Tt1eHd8LyUIKjYWm9gcDrvZiSQdRralPZm6uotwjObVY9OY4+Dejzws
LzeWC/NWvoYs7zrQY3RuPVaZTHuIcux4Sgu8fwsirEmVDonPI7M8S0vB0qphkXzr
1rcc43fR9NgYQgsPtRLRoB42tKkeRL0vTzp0TCKRR/yIooH1XAGkiMZs9+oSBGuY
mSpBC07TBFpIu9KYJRKruCQFYGqudFbBjH4b347uC1zrb5pNZjz+e1LpM54hehVU
vM0iT5Tx1/HeM7tn/ycAHWm3vHrnePy8P+D5NAmFIc22e2fZIJgXgkNVwEDO62ds
NfRGlPiAfjNKi5icvrdfSHzXItkBTd9J9ElhdrOEU9lZC+P/l1JUKht1LEhsurVm
YNdwIKCSP1TDThJSSiJD0oOHUgHF/n7HkYsg+h69lxuFv4BH58oZcR9HJQOZlgIx
j68Lh2fpKdlyuAyk55Zq0Lqfq0lXr7AbaM/l9PJaIUKpytSRIdWYEle3RaKdWnr3
ztQHCSK4howVnwE1AYrHKP1tecRR7UeCajVwNmOpc7rmJ9DU0EhbozwQ6g8vHY6i
XtYh8CAUdhiXbpauLKwqQ9ONqOlNjOnHwgwIlsCIikdlVods2kalW3xxsR8/zXq4
DPNIYgjqp/xpa4OHi7IJ+t21IaWZI+MaRhw1dNlhfK3FEp7vH0FdCJ5hqbRqf3/5
zTU6evFT8+ffTC/yfHxMiLrurZuAhzgg6tveHUVxpyFy0fy8+jK/2FqhY51j/zr3
1YhMw1DkLQ/Vl7QNgWg/t7ZohMSuKIQyT+OUa+Sb597HfKs6C7jWJ5D01FY8qR+S
0sXQR/X0ZaiI/dfcXpDNpFjp8lgtXem/bjzEXO+CBVz2Ih09cu6jB0Ucc7JmOOBl
d2+gbq0LNNa7E2RIOr51bqlhL8l1s5Wk9Gan/6QW/N0Ob7bSNiYhzfKekBJfvfzP
mOuwU/o8jzI05vkfnQt8JLDJzYWYIWfPqI1vM5ffutnTfEtZubNazRHRDXZ4pYS+
2nZL2bgMl7pnYXBCng2fpWI7iaQqYePxxDizylxhWB3p7WNSaICB7PNkWIcPdyqb
gH7H5PR/h6jw4DdfRWbH+d64EDYqsOp0satm1tMqhbAoeZJw+/TSHJ55ofg2WQt6
vHKZJNDksC5YIqVm0U/TIzYEr2xWIDdtAJQ2ZAxRrEl/mHe1HLWiLfT4Q8SQFq9x
ZnNshvgjM85/fPubCLnn7lwe5Ter29SmzwbeHmYSjsuDEjfgxiAQxrHTdV8ZAjND
z4aNMZzYFhCYspsqhxOwqeS8HJZcWo0hbyZ3dHssmtE3sdmbxWDsK67l05kWkXb2
ShDgjE1o7dReb0lj+BALVY73w6uKZdp+mtNvS19iToRH79uswn3eEQ721m6VXgFA
nF8K9EPdOssVaiX6/kzd85bdanYBmWdh/ntG+M/zCvhPAHMppImCZuFI9ajhAMET
yr41IOBEKk3QOAKJB2uK/ssqDMVTL+zlGAklbXeHbT98+cFIN8w1w5iixLRrTUk2
Q0xQOnATdbYpQKBxrSbVIOHV82Rrd55fR+48Dot3aFUcjGkibiT7SWMMGJBYSJjv
3Woco23sJgv4EUdi6G3yhJJ7eQM4H3nsb8PGRuGjXo96zjOma+rdUeAejRs/UwL8
V0JPA81nT7EbT27V1V0k274gNvX9xjkaoCeG2H1qxxLTKCbwV4wSI2O+sbcATBUH
c/k1tPXQy4ZMpd9hBwKdGE9MgrL9WV2ZWO1EKK0VKLMpm8M7Fs+nu8Pu6ogrDpPL
QrHFZaDDGjfx1lghc7gcTwG3ia6EwEH6LcV21OGCjwhML1aWhNHRbKItQZuFRGL6
lJRaE3Z6E9vQN0O2A2SqtlYflYEGSnHN3twHe8KbWQgipc7oLpW7mqyWjyApb+9z
XSm89tanzNdU0XByjJuJ3/e5iSGPkc7AQKW0udbhLAY6jCzOEPCT7Gn/+sZT+v/K
EaOwo2eOx87YqPs2uIBtpLfHx0ggkSukFigNc1tkd89vSQP0PiRpuEA//iEvoswD
DADpZA6uw/Wp/zcbj9LioRph9ZLD1M23WF7C7ibQN0E6iTLmiSWk+QvGJzYh4JxW
h7gBwQ3GLE8YAshFU0yGLNk8yv9bolys+wpdCKOOintdseVjoFtTvLgjnceb3Ur8
d6OD9NNTQaPT8CsPS8wepmrj3p3slkcSEUntU3RBLJgrRAuLSRZl29gjaZiAhp6N
lTTADBUdxvlm6eTESvykQtxyp2vQ+esRgvnIV6VbQRlJ1lzUVeHzXz2LowAcDGFX
jZAqcQ90P1WqtPv60bt1Y0gymcLg0rF/f6mb0U5kbtehvuQycenPlPdkQy7Hn9IT
wm09o8JfaOFPDEuuW3T8woig2HYpnkncp6yrNjPAAhl5uRF1kuvPbJzc5MmF/zZz
vA1Q+8t4nOt/L3AOttfaLEYZMDAw+pY15/Wc/hcP2Pin4B8Dcm3qXWzTZ+qDXtRZ
34QDrZc3n4gt/X8Gkq0FhBMOaQWehYJZg635dDdQKGRKkHzQBLzDr7xCrjuc4+0O
yogvFVzymnZbQoRdgEjSZrnHb4KGNyBY4zn2ML/WTxNcJX2L4gfn8TFb99W1jsCF
0ZpmavHOWVwtJjA3TqAV1hfRcpXXqM9UfvAaHDdd+V/yJddPnr8+H/buUB/Qk2JS
jaQ5p6oysBJ5T+EsPfMxHlTOwyuA7uYFvShG70zAQ37Pj8vanTmQjQ03AJbMVhyj
jbrUlrXxF3GYNV5i+WFp+cxbDMMIw9LsDuuKL7l+p9I2j9yfxCm4AKXhHx0fxvEj
WpPALHAJIdlsLYsLhLhV/FjECQ74agu82Q6cdwUv/jzPhPm7HpusEPAkGd96MNPK
G9AxCxOaSPm/zunzY/xt0Mj03ZOZ2p4Q5N0za5jw44xIqzcIB4Nvxo9hcJ6TjxI7
QYwvCQFoYzXfLDaZCFhXihgQ6LvayZ0FMUGjzlVNzPfOxNYr4LdtlDZAURaiFsbk
VDDkL8ENvzEi00FWdYNtOoJG1DF985287aHHLolcb4Ws/NUCL+Kd9W7sLHZF/3ow
FvFyFQzl1bLDfMMsm+G77N9g7LBCQPAbeMiE3iz8Zni+kX4OlpDd3bLkGErkPVeh
59dSu/NiU/l8K/MPMCCIiSc3saz1Cj6dpJcZG0bLFempISwFlWy4BFjbl0Bzs2mn
FQ3SXN97W7WTIghA0qifbY1fFSoKOtnWbnFXB8vle5Co+eMCuCkmAPqtu19Rir98
ZAgVBECsIIh5D8nCfpmgONvVBYqG+Qk78cNOs1wLSrvNGXEZH8FmwsY6GB6J00Fy
QXifNV5gXuziNDPktzM6ZovEgvGTBrgJcJXhqZhbwxAvEBeF7ZW4MplVzaWJKqpe
L3+3a0x8AHyQxmaYStoKMy8Osg0ATRpCL/lHo6vqCXMr1VgNaYy4R9rNVIELrEDG
fwVG4tvYvl9//7dVJiLtFRt8Rac5WAtOqW/aYriISovbQRrZDOngNTPgi6XrM/hX
bG2mFh4E2SFIsTEEnkkBvW6sqwstV5rtEs3ty71xSy/AXnMNv4NxFS2UUt4EE9nW
T/Kj6C0VGaCgi/SQRMegzlpJ/C1PiBhbt/IVj5NqbQVftztW8C4vmHteW++FSo+r
JNa9nj7LS8jYCo0ExVoyfv5YEXlfTjoNUjfG3ZO+T5atrTMAlr0wfAYuYQMmj4mJ
qin/XtTdi2Z5QycfqwQMyZ+PDENmEYBGpNXzHqOQpeI/B3m5j/NxiU1wNGXMi8Xc
J3a+V0CNM3C9M1+EVksjkxG2/HB6jCgsBUefLaZ0dayhYNU58aCjNwsU5yEZM948
+JFcZRu2TOX2w55SfH15bLoE+nYNB1UPOAGRwwRm9G/Vy+oSp4ZAXZoNAlOy6xY9
6a7iKLeqHhCSrjwJ73uO2Eq9sQtsrAdaa+D0yqo12qOYEDU2NMoXzqcuz6DCYYY6
ydnuAyHMmnpmiC8m5ExkefB3l4LL7cPb4l7GfTbWJxOInylXVXypW9/QpPu06wXS
xQKtpf1+anGFcf5XtBkdGr1eJt0zE/vNi+d84/wqtpfQhEHgN2Osicu9bTPlar5S
l0idDghv9tvXZG16iLINaaYuPHbm53muZgiuwmnXhqqipfI4weWuCx155ESl3ZA3
QkD61hAruOdA5MoTHRxQH03P5oVviJgJH+Vlcw/b55pRbronxlvPvpX680/RUVyd
ZbYhgy/y2kbxAWThFTBZGKUwAWYm+GHzuAHUMIHXi0LI4JVmWzwIJEPg6Fju7+CO
LLLFONGnJbcVb62+U0MBgimVuFxr63yG55D8m2DYDb0Wb9x8G8JHJLXXV+DTjXP1
Fk2JI6nlAys6Yeo4w9r3arfJLFltVZIqk6ylmhJ06hV6jorhL71PKml8crn2XRhF
5D6n8cA+V9avW1pRSGVuPW0my2lbTYNnO4ybjTDumYvR0GrOPSfrO+N468XOLDwO
z5MWEmCWyiFZOAXiKWeTEPuXxT+3UcmFAPH40cnDmTMioYOebGl2qpGc1MeyEoQH
UxzYUO2Ksmt9mkFgq3TybiLusXil+kN1sa3fecaTM1Ic36von1wW6sPoIDzSq+sh
gnALwPsw/YSw8goXVE6QfmBlFq/6aqooKHoGWRvuq3GnxFj1nXVWbfrYegJ0w+nw
HunwT9X0VTmZczNYfIgCGqTk2UhSVB8kl8Qr00jscyXSRm79kFWXIpIxHP/tA9dS
l6zoF+RhlkbMJ5ZexleGWYtBux7+j5VjERy/YvqrsNM2Qdiw7thwnuvtMpn/zUTu
qZ9VBJSH+4G/PeOAOs3ytXwWuH6Bil0kaP9GhXlbAAHaLQq1E+jltIAXAWsDoS+t
p00aOqKbnWm1D2wUapiRq3DepeOgFANeNR4/q0zwf7OsRIHiljvIFv3GhEpMgWzV
7G/+0Ed0dxxLtLOaLXWwGbhRzoNodDrc2lASY0yGuEXO0bPgRCjFbo+up+Mt9Cxu
cm/rvIoNToSVE8602SVQyB3zRn3NY2xxy9DPDrGw9G3csnqCFQIOUpPhr8kK8Xik
1JoAAEJPrkOnAp5Hk8zIwsPzUjmw/0CG+7x49kqak6w1lILmOOAL/wDg4+ZqwsCW
32Xr7tDEBO278s3jn/yeYrsaHvVfVCs/BU76MSgpX8imURz20pigxQg/wLfGo2/a
Gng8VCVcqKZ+pe+dp3GE57j1eUIEf2LyHDndeAitCqGNj8EYZgb+i4EVjLeTbVt1
DVksntc1cAeiAqMnncC9QeRNca8NS5zenKBcMhnIrgdxuyoO80SJ/yEma4odMDQB
ZUWoo1ADl3Dwi5oHp2FF2Jt5sY7eevx9T4wan0Izw2MzGp/oBee6m7nQQp+F/wrD
A/tAkzW6qhF/iwmHrC2mQxqrHQ1QCGSm4b1ybo2Bfoie9JPkuUT7qwKiR4PrFu7W
Y8HiAJGy2RHdrnyUpK7EazmvhoZo6+tQH8/5qVG7Ox6zakOK0c08hks3BzY7e2xD
exiELaQtS0Hu0fTmxm5MDWp33K63t5TLm1b/BYS2NCn+C8/OxegaCjrtKzxdaoOj
GKP2y/bO7I0IzV680o+TvjXSV93Ap2E3XZOHdHYHQS3v5wOfxaE9XvzbyGFJGcFs
DhfDm1bzhA4OI0Twl1ex44uUo3l9+7hGcOboAA+carrBHSkviqEQ8u5CU8rmhbWk
QQsGFRk708+Joun0Zz+R/MrCcL8+DncVNJD6Wwg/bcOKZz8kWVHTohQ4vWa20lLw
qZXXIWy0ylSfS+87uwca0OtDEnd/Q9HfxN516HLCcovYUMEq7eSXYCl4Tde0uMF4
BBdqSzVa3hqdRcWmpmRwTsIe3VqyQ72tacNLDxwTk8xSuK8395d+Kuj3k/jXfzA2
iLQj74Vk9qhMEmfif/0Bza5dNLMO4ELsAakq3NISqa0DYIapUX2j1uKa5BRwgIK6
l51HEUWrd9Wt7eP3jgZ+nxAM1ssJs2s/hS56A76gMg7WC1fq6A3gkOnyOijDDUeJ
Hdfq+aVWPB1ckj5Fw5x2PTnbxf8I/Oej8l1RPpZeRL4oxYCgFCRbFvb7uZVqa8U/
ufdMokAVZnK0MOFi9HlCi+RY/0Maibx42caF+J3asrupO2RoPgasLwvmes0uHriG
s7Bt/FJGoXUMw0B6KrL3NQOlRHHFSaO6YJwaqmavt18Jkz4Y2nERO84+Qu7bYNXt
QRgzrssXJbpGdIrFBFsl85QBZMLMzBKu8TOL5K6mlzs6JQ9xtKklLKtVgup8pUpP
hUN/mQCwGPDjt3BWYmz3H8H52lhoZtQdBCb0kwHWcAwtlW5jgCKN7Vg5O4AXFeKM
hG3sVr2LcpW+pSdjIOQEADaEEDqysZlhKa8tQF6JJLCpi+5FxugQvjKkvmUKWGkT
DlCdRWjjAwcgSOXHoceBNZQqAxc3RrzBMfXsBurR4WwcNhtVQGYorZufGX+kYJeo
KjdMI1TCdHuEvHG6shFB+wUEU7rxYSunXCsP1knXYffPZk2Ub6j0eX0yDUDjFoVv
EUrDgMp/VhEnXtyiA1UfTLq9+ZpldHbtHqyb21VmdihOBf3JboJDkNQVhxUzIXnC
ieIK68HG3hII8hkAJTDSRvR5uSMZQZXJtZQRaiZIyku/PbP6JdxZ3mnIiP/U+x90
wT2Zfj6veyT0zrAfl74LPZw7+0Q69823N0pTVTWtV+irXAc07XqBV/4yk3ifhcN+
snZvrx4o812+U2hsJx/SpDvAIzXH9J5UsnfDJngqB5K7NsyUvhw3rrY+AafSoGLn
V0onKw1En4OWqluMjsexnj7zFVtYiRZXEf4YIC3rv5XUjdyGAgxWu8R6osMBpRaD
lnfJSQ/8z0fYV/+g0RpNIGacvGHuxdb7L+0Mki88PwRUGA+HYBDZSPjL/vHxczHD
OPp36ctGbfcPStgcP7iPd3qNCW+XzS00yIQBjVSKUp/vsi8i8MZe18rZc0bEbdcq
/sbeL1o0GM+Y6R9YGhHNXxUHs8niCT+vitEwCWUEiItHJAp6NHqDIm6xMUMpyJYH
Vx3Qum3k0MBL/4T5jez0FlkNFyL8zeC5USz1gonvsR1NU0TcqDaU/LzqYvH8d3o5
fZQlHSmLVaCsV9IEwArujPL/hY4yZmShdeT0grt+n0dxfFRH7xCnYSD9nYwqA/C4
cR+AN0/FBFPNCzeABbo9T7IaOaf7Tr/Re9tkugO1QuozwnqijFGMbSIbuHxCrdRz
Y2SECMlxJ+W7S8xgOfleC7+gawv1U0ZiLICC4MjUnwRbS7589QwnD2sutEVIqf4o
nV4zLalJN+Isbj/LLZbUUH7YqubEmonTMEchmBhxwkNSSHCAw/97bEZfmZHJOjLa
ZWcMVR7rGtqxV/dBZiMpENnh5ogPPPQsy8P0FqzRy5vrtPFkMfX/d26gfZLYnT18
2yUXj0U7T6f7NBvD+7zoq12bbo6+nLpqMTI1/I6AEiPb9QiTp5bZjg7SvIoh1suZ
LWWHfCgjBsN3NbkwoWssUtj3yOhc1l+APsSWqKL5a2nIdhy4+yFz+qy5LU9DVdRY
7A33c4TWamaSmsZabmBcOPAgHwIlSruXmRMkdYl04O1jc8KEEIcnXfPa6gyqCGOx
1C2FuHAjx0zl6mOli1q5baOzPvBzdiSfogppJbAAYgH/rFXQt/Ufo+SDaaJ+xMEE
3sgjQ0NZwX1UTt+z63zwl+sMcaZi5wvRuz9JYgHmm5qOfCPRoglFRnBccjkZDuZB
SJtFnvBZELneLymg8xeF+HgbZe3xqZJQjuLsodFe2rIgkBp9Q6XPQg9XsLaVKbhI
guT8vT50brlIT6+jEkV4e1S1KvJpZsKaj/MuK0tz/ux6XNIpqQL/FOnL4c6bmZUA
TZ9LihslLynIhcxSbznmEkISeAwHy73tvMyfK+gVhRLpOMNVg6AUiAZsvm77gXIK
JVtnCuTaJSvnIN40d3j2OANIY3bzJOiYKzO8qE9HRdtmh2pAAqOXsFEH2B1ymSKj
ZBwuw2mvJ68gFDzyZVRjPPHqocWs27CWQpG3c4dM5fm7GtNb/3iRwQsqBQAFjMoy
EH8FLaqbM//HtOIX0kfXVF4RggGcDftKyxriBn2WKL9wNM4nro9TClLbdjp6+loz
dKPNgnm3p4wjgd5u3Vo+Q+rjnomxsIyaQydkbOPx+EFKkJT9GRQTGE4halmrdwOp
HQqcLhyHy3qWBzg/cJOSm0S2qKbAM+FPUm4EswNrcCM4x/xnsCj3DLcVVxAvJ9rW
R2BDMCmt9rxK/BXFYbQx2AoeFkqnGnt3kx2vvI6DFMrjJiXxN4O/UDFJPAaxdFRT
Z4DjfVWRKncOCU5uoG8Fd7PM1T8/ay3Yz5hNb2D1AyvbZ0wenT3mlIXEnXhAHwWX
Q2QDoRWJTz124OG/he4NxeeLU8/Vo+/APKRP0nzjRHIHziZxtfTmP302vbaqAA1v
p11UAZXJnVZ9U/jHS5Cl2l60acEU6lP6H2z9i5YtU0Ors+pMAK/JvbL5h9Fzjh+m
14qOR2T9NpGQeEmh4tBzSzNuFaOPZVmX2HGn9mm+khI7a2MTZyvGRVRWDPV+oo3e
NywanNFVOJtiyClKSgH6mN5D2wv+U4pQjt8Q0MkfLGWZBiE6y6OahsFlLaL6m3Qq
uVfoSvULt5N2FTztD5hS93V1eyo9g+hNK1fIqXhDmaIaApQ/BA7koNnTIY0tbFBo
zgiutriXlFcfIeV+rOUolD2AJNp9RLazSK+PUCx2XPo3fG4GT2ZiHU28LodYAfUR
PQ138P69T3fYRPiC1HRIn1k3Jj+rPkhKP6eIklR+5Fg1KXg7IjMb0gVBq7ifnMoa
lvESnTHs2qYJ6RP3YuNXofRDTopmC8lsfIbortVihsKHcCDRjtHiSSW8NXYVve9s
063DY3an2J/zy83zcAjpK4D/FiGnADfg6PFK7VfjK1i0frj+pLXxH6TYc++5uh+7
K44tiLqrEXYwbJs0DapUrzbaySjUoeaS1KKM1dM+fr5PmcPzumiLGzN35uLWWBP5
RQutxwof9Qj5yVRqu0ismhTU3Z1BWkkg20bengYJF5FI7QtZDKOQKq9atrDWR+zv
JROOP1Rn6uLX6QkSXJIPdPMKkMtG+/xWVK5eJNK9Q3QOJAQ/VueVnv/tAmGp1Ncr
ndDnpq21CRsFDnm0wGcVEcgaO41kJFsaFZ+Q9PM4QBnO4DS3F6IDzul1zcf0QMui
8r28tB5tliz4KbhziQNu5QNNsdJvO/dT9osu9ZCwR8oD8QnfFRFRU6536lonGKp/
P8W8+Hs42wRvFH4F4oIbwQ7h7P+Ax74IL6Uo7jmzZPbSQov7Xmr9lsaMidNI/io9
ZqlQeReQcYDHNeml1UaKmA9w3fQkp3nKShFqkNKXe2snT1hWI8zbMTgrS7OcJrFH
A9U4VWqsJSu3oNPxktbjPR3nYKktyiIh1LUsFGLV4MDCLNjcIu0k1hB7nU8pXyRK
BTu2NAgY9sgUojsNzqJ1WJzUWLdiuWJdA0OFDB6P+vxStXZg7Oalr8R/J7c7ksg1
OSVhLYWnFLSvOoUWU80FmWn7k8VI5tkPa/2X0ekkBnQq0alTACwLM5SY4SkxfgYK
y1IxSx7SdVC7Xmw6TV1VXkRfCYVpKh68zK21Nuz4J17FW6Rj817yco/2lYyR4Ptg
LX3JtL8CULLkYSxYY7S+dsv4VDQIuU4bhuPpN9rwwsyT2REeS+mlDaHlnbfdHqZt
OJ47vgk4qHHIBN9cKxYemONtRcil73x0Z5MomHE+ngNmh02ya+7+VDYxNlC9f6Jb
ZCIKFTgMXxZT573gJe/nL2yEP9v37AYdkrxfkfdYFGzOxim20TCs8arc/o7iafKf
QbMM/lyMmy/19ZhX8uG/shjWcXzZFETUNqHPzYoutc+4hyviPIZ63l1Bhyfgkj0O
ktwooXAT2w26vajRaCc4EeTAuEBAZxZBJ2zMeA6iizl4Iot63AB+MYLMu1EoIS/3
aJUotVZawJAymNDnPD2yYrdhvawpKw05kNEv3jL/n/MZbIigLsmgmd7p4uJ3pwoq
fC98B7Q4/2TDeFNE2BtRjKYgP6lWMFaOTQl5cCj7vhuCG2NIDuxaibecGqw2FQ09
yj+fi0TvGP8HdrtIebh3fuN6GbzxhQe7pQuid26TdMttEccTuYmpIPjxUBJL6rLL
mJtTexz2TykYelqU2PeYMa4GJCMQxMVoBYAWXUT53k/7pWYUyeAtEKf9xkfumwcL
5S1eBqSUQ9j1mnxP3XRvG2JTss1h41seQCvAOEeDaEFYb5cCcWd1HLr4ggGWS5Lu
TJCbmVO/3oUCTHV0t/7yYCkW6S5CEn5yQ4ZLmnaWUFz6D/RUoe3J3E6s5yYmoHDu
9YKk16fRP+WUPVEeZz+tF9JmC6UYJwetkKJtsu60njKGlclxcErOWSwEfs/PgpEZ
aB+YNhB4rXcxr13aLJ4+cXCaHSJmJThfWRPNQMxdfJynjEvKov94N5YCvy5bwZwe
S6BAq+Mrzk1wg4u/OfRPmFd7+Fdg9FS5Or8sf34ctWTLBLsKqBpE1UodBS0Mp+wO
yQK57a61q79uCDVqb5r0fSUb9iCXvxcEV9pLeu6RaDAyZVMk/bxtk7v+/obHakPW
tGgzq8YNhDWK3PFU0Pok79cKZUKob/DxseejxUZL3NnzVTe+fSxR4JvJ91IfsL9S
AyfbebeZbsfE1B0n5l7CpGQFzLYJym5BniZBc3dXZ24h2sd678dOOXxYr1eMMTz9
G6kTog2DXWJSNRqJ7RnKqebZCFJ0PNB0kg4GRq2OZOuO8eUPWtx/QSrJvHgC4CDJ
sdGIR31u5j7VEu6eO1Jdw1N4bmO3i8XTIxHuZJE5sJo/sLmNoOLVJQP6fNDuHVGI
sAy6kPTl1V6vjkhiEecCJ8KZNxsCOGCsU31Fj9gjBlCBZYXNYiVTWOam29EKvcwP
Q4w9hsfjt62bMl5nzlMcdgr7Z0jstygdZU4pSkztSxY9Tj46R3P93aJImhBfLLJg
J12oIcJO7VslCheKooUyhbs61aupFhaGvpIhwqsYKgkM8B70jw9db/jot36QDhc2
UFqsQv/ely+3XTSa4AjKK+LjoFJ7/Ca1ArT41DcqlCXh0Jcv0OLji8yRME4T29/6
yAOeqQ4w+kGVxN7uHM31BnP2v63CuxBHDa0mbMLVeD7UsZ6nYGx9qoQKkfHwRyLo
oGagJZM3OMcv2v4w78MCC7k58h5q6xVHxSGdEqYqz3dgWHDckkNmOlv7DIfZFO6c
L6Sha04z+oqymW5FZm7vTkw+98gpnVdOoj59+VKLmO0URyc5hxdqU/YnKjDs8fWe
mbyO90s0IcinrqQBC97hsmQsJ9cehmOUMao4ekgd0KsRDAZEqDez3AAjkcLsEPwe
DVOTw5N37+vD92NOAmCWJXqbiy7cDLDL6sROIdaMu1KVQvm5oAQJW58OpW/7YtXX
3lwW7pw9w5s76UExGMptOD8x3pzDRr0TbMb5dD2C5EpICug/D+UX4/cCZFD7BjcN
Q92Rfw04CpuNlOI56nVgOx+D244b78KnyABabjqQ+yqKVhE9aJ+M2DDFZYltqdon
v+gglSvBjf8vNSb4zNyZK2BVV49LDcY+67lVF57nU9Vy8ATG608SFEy3VMI3K5Ad
tEmWFiEP0YLMYjJB6jOQ0jKEt3JY1yLWOOPukJ1W2S67v7i6jMeup+4JwnA8RISx
uw9z3/HF4ZEvdlhMoK2uHX0haMO6Ck8YT8IijaNUClsJfEr0VmuFj068Hf21wNOl
kSml0boU6HSOmjFh/Q4vPKdAm3vprtoMHryl3m7Zh41RWcBZGAAmMenSGwXGFnHZ
Rprbf7O13/MeDKl+VHS/+KpiSx1bdYBE+w9+IpVj2CWUQRj7lg9ECd3AP9/JkMbr
6CosQ1U/ZALzUEaEV0cmWhnBRYJIvuCiXq8OwLH5N7LSY7xO56GosVZa4/1UKwqI
uR34zlQxh0JbIoyW6X7CkD6g27GYZ8sKlm6NpbjZX4HHts0vQuKFdS1up4cZ2bJw
cYaBfGcdBTTTeYeY+kpLLaui2NbBkTOBm170IJMPxv4odVx7I1PS7YzlS6eWjAiW
+NfqYEABAz/fEq2m2VJ5HxkhVwOIbuMdX+j1NdCVP1NNLwsVK1ATLmAPAa/Go5CL
jsNXGZYRpdURL2JcjiFrtCdNRc80r9NI5dIsorydFx+V63niAmlTb1hbrA7uowuN
wKnKjLql/qLSnPQ/MJpRySe+bK23sSVVrDfsZA0jd4vAgvcvB2HKws2amEOu8gZ1
O1xpnYgeCAVOWq8n8k1yhvvh+VJic4jXQpi25/lBiG455QQrl0lAwg3piLjM3GjD
lws9ngx+gui7raECXO9Tle/VnVKXAaHWemaCaAOD6Kco49D2+WWLEZWAPhckG7QO
J95nDtzmd+N5swha2nuq9Wexy7EzvyyC2Us+arYE05mcDhIuJipgd3KWUNYKZpFH
78CfytMG//IP5NWCmJBWO8TpsE75T7bjIunrjK9UGtYTf1kRbuhYJFs6vqj05hxx
pirGOGfNNtE/9IEtyyGq8HqTZ1NlkMpjEXhUyyjIBmqrmjA1FLm9HvD8S+HK1Vgg
A8ppvcUVovylOfvMz6s7GIDhUrWWep4wPvadwic1Za0Ptg6C5BTjE+P/vqDNTRfh
ldhcFPg6X3SzAOruCoGDpGp1pIH/WIn/U0nLNiDV7SyB/KwRmewtdO16JTwtOxpT
7/QExj3iy7DtdqafkD28dBpqpJPfANWK+bu0mHMhhWVEY9gEUslmoEZWkBUq3K72
ntX3A7scLjCXe5xW05BIcJWIKXX284ENYhQqevAOdMG87lP4t6w5VN+vMxMs78IR
XsummeeQdIt3MvtnWLomENIr9ZhwUBG5vaibU219xdNUhbGhCVurcdrNhzSNZSx5
z/JpXoZ7gsTnAgEt/7yCeZ12HIQ948N8Q13JWh0ObJc2Vl+mFa5s9q1/Hq1e5kZl
Qmi6NwQUqG4U21SxsfBAYeMPZ0+BU0QLJ/xmPt25Wil6K5aXMSm5HgudNVAZoQ1S
aywdPRG9jCJUw2MoY6VTlik51tbBpdtteU0q+HcnXZ6zFA1stLcxqUh+YhalGQSF
iCQY8dxnDL86iN4qR9ASBoRZLuVyL+aNmRIj31vlg8obdrtb9UMqS1zgcjgedLvA
4LS+nLF05jI/AGh8QYZ3N0qiyfyDvt76k2X5T8kx3uvr/sCvnktCHhvHe2D+A+iS
KsUDcBWIfik304dL74BfgM9GGJd6/YekU5p4MnWKzz2bZM02mZAfrhUIKTK60bcc
+/sIls8/7IMYWBRvGvG6pxn5ogsUAgOQp0cV2fUnZr+dcFhhU1C4ondxtCccvfuM
GPnsIsUJlghfWeWxg1rNn4gZ6MRXqY0Tz1hdlYeSVVovAMX5MdvocdlMIL5FiWim
5UMuNW+w4qQziGz5H3+fnnUfWAC/PB+yRz4VRRKwL7n+jUNDuwmj1kgyzt8+Iwvf
Ja3kzaHHX0YOyb36aFtTeSjtQXHZyDfZFDKGmQc0opI4p3ojl+fNAicoblh4sXzS
p3KU8CSNrmcm/U9mLQicXA4JVJXFti8h0TOFN2R60VJCKVq+gkCtER24CR+nsExe
s3070dUI82TIzrbHjNLy/tAWpsnimsySHPFGiDQiiri1l9kIrtCT55rtQlK2kYX9
whQIBgaQKorfTBGBkj2Nr9LSK1eSH0GChjutxP7VB3EmbQX8eVUOGsf3A80da1bu
AigSvcwb4GWai5eVbxkECo4KyJHOTXJEG6KQ/sYOBwlVaoERZKqQj+wfImNyn6iS
ROnQd6PSRd9PmUVbmaYD5EDK7uzsjj0AGZ3C/3fHYcst3bh9hdXjtPQz5FvQ7JNu
ZKe+YvLFsHy5j4P1W5tm9/FwM6NtEYZCxgufPK6mVUQB2Hi6BKTPfh1RnVxR84em
Zuccz0VhrxfUdyrGt0LEDKk84Y8bWKY3nLHf0hWjOUjiOqLzgultkHkn0JHWdt+i
a3c+ocgwdO1uc2sDZnSL9hW/MdyGWYriKp2iufRJeFcsUturaRkBa2aW8q0AmREH
4Hf45q5LgIK6867I4sXVOp3Z214a6FMq3xN/M1V40Vp9v1mqRwrQbinMBLlHb3S8
Fv9QU9rQ4K5hEA4YERBFpomLdStSMaYKSFtucqHJKtkFIxmdIJGg367gKjVdm7XZ
lRfpcjTP8M1jup9LWJUEsf2hWs7lN19xKLYgsdv6iIIhTwcf5c2m8XzoGq+luqS/
xZXhteSl966ImQeHUz1dbiP8z+vSMvkcnap1LBmV4LIe7K6VbglBDMwbBon6MQhy
Vo0HZ/+bs0WhGUh+i365s92GtPx+nhZov/UJlRBOpciabgQIpnmdUwsT9hSgaKdW
3nf+C+uPYKLYsyl7Axb+CC1/HWnXGvzKYETM6kT2BA+igZZlvuFf3Sm1YXmY2nSV
bfuvtlQ6FEKT9OJ649EwYzvaUmis9pNC33r897UckaYtlQitP7+skJbyYs0N0QCX
B6y/9b8hiGXMSWWRbKJbqqkCqdSZe5jZljVQj5g+W6f64xrGcFU8nstWXTouo68E
hR0z6n1nQKz+BHY6/Y9foh2sa5AbqPALHfCDlUBA99WBNSdv3sef98owMm2GOHiO
dJKr0m+yeIW5iF9vFhfL5k7no7aVajHaGg/P2xPekQKhf+6lne/Dab4qm5RzFwHL
Jv6/rmLYV01TZsMebfl0wBaIe1PAronuZAPceZ7KF4z/v0+PpwBno5NNW4GK1RD/
xEXz3ltuK+NfxGMlv6cls6o5t5NoyMmni80iVrjBdc95SH/iAi7qcNIyGm8lengG
tOUrAk4Bwzm9iO//7fYaEFP0cNakDTrUJT15dPbv5uPMc5adNTRtx9z0nU8EU4D/
MoKfCN856MN5RIELWlZ5A19j1+gz/13pvjgDIcnWtbmqjWCDa/icr8gvbwioXRTj
gi9VqQMZ8x5u7QN60mm+2ZWPi21BWJnTmJvLUUzQ3oHuJWkE/CVW4Pyg6cS4xiDr
I6L5Rmb+jIxp/p0QKLr8r4PxBx4i3hXlxCmb4nvEpGMkWv5MZ1bcd/LwmFAhLRiz
ZHL/WWcP6U1OewuGoJR/GvHMDQoOWlkPZ9kVi5J1S0Lkh+DJj034wLJ/kOSu5z2K
9KfW48oeap8pjr/Oi77+Y+Txvm7KWYn8HG7/kd/PtOEntLxsGewfntEKMi4gfQRP
DfYiTcVwgubNC+X/Q0UkAU6gjsJ9LKWCnE4DGHJQQm2Bd27jI/NvsOKsbISwgJEQ
GvHG+bXXptAZFXlRRTb2YSgjItIABORLXgcRsHEfQ6JxMDAkl56Vq8LU4UDuyCcV
PYv0Y9ngkgPlCHSTvS7YBaaB2S2jAxSOUILD0LE/Cde8A2JpuEZ2IKK8KKo8mVm3
PvnlluCJ0aA4R/089cZD67EczlgzOzEu1VnpOEm11P+PlC/N37PYNGCqrTjtkBLa
weWnr5oPv9maffeXSA9jXu8HuX5NdDWszXr7hJ7Ma/xjKVBDhXY30ShnGgW0wlv3
bowjYahH4BY8BaS7G6AY2Je8P1vWtoRb0fU+xLpNOTkVbX91St3f383OS/t+HgJ8
gcnnLBNbHW3b6j7uVah3F3R8bIk3+FnVT+LmxvCFySBl0yzg7pbUv+QaV33eTc2a
dRkiD1D7B+PzAKgWi+HOuDMNuzGrqUr6/tjgiqerbawQkwiptCfIbA7o+yazmIBD
8PNlazxhNVbnLb8FYQGzSjBZmx70QNP8UN2iMv3HuZUR/uzcx4fFksARZbw2SMeO
AfJbm2cjY6lIInbUTJkShqNAxk1KMzuvN1ZgunB+A6PLYxMcGaZ9ZRWq0vfNv++X
P1M5s7OX+frVKRTQ+09EvfW34xX74r7bxTLVVmT3EVPyE7FsIuCQRmk0pJJT9t1C
cT/BSUNEoe4ogkQShLAd1zcv5TyF2XRrtsb/0xo/pFd+C86EuezGS621rs64H2Pt
+n+4DYQR2wdzJgCEvlGmojaMSl/vviDTAE2xz5G6zgetqRl+g3ILVF/RPI1xUfg6
FDo/R3cEtWCUoeTiIwPqj56Nr/xYqlqCMBoGQpK8rGkvDvBN0Aeys/yYNem/Jdaf
JmACiDR6JKuchS4EbfdzwvuctSYETLQZSa1V0wFN2QC8pQzo8dDRRkUhT4TurFJJ
aMUrcIjOOqy9sX8F2WS8P0/GcB6SHUM7H8AvbNsfncWdeghvHYnj3XgwJFXk4wmk
43/NvVXJWUSHsEMW3hEE6GltaBh0Qxgwlo03LIHL8R4HDVWngg0fS1xUcbTia5fB
Sh3sg4bo2gmNy2J/UbYR66TFNzC9RXfny/DQ/2V9REtZ9R/dnlDBNpD62YFWDSCP
tCV+NnCVnll8OVqhHgOnEulE6FeHiOYihsajDP4qJN8pUErcEyttODib6Stscxoe
BuaBTu52Itt3lqTrewT/xUIVe2aiPVjmAv6XV9vznPxbk6O0d8oFSqKTYktDWm2w
onGhYb6oYBcefSHXOosVo6P8j3LTN+bzNoJ8CyOU35jd0InmSceQEFBAS3f+nbeK
6wKUUkKXckUQAtv8XEU107dLV8WOahj2NPgITBKXYSM9T10QeKRzE6g+FD1ZIMLr
dfE0xCk46I1ejl78A+X3kK63xav1CU9oLdb0RInD3W+IxYu3sx3uoP+awEimdGoP
Yy5CtEFzRsP2ZI14N03xNv/+ZhC0MxpHQhmGHPyH/5wsucI6DBK7b/CXUWgTbaMN
6hPT1/EzoOb8iXiVLi2UIHWcT+YmafnPpz8F2wcl7ghQ3SsOcknxObdqsH0VJd/d
cltS00V3C06Cp/JpnMeMXLwjdIPLS1pudGqzHo8tlw5FoyGs6YMGTBB+mND0rj+s
f9nsn2G6kKXCdpnuc/H0PoZbjsN4Qzs7m0PuK2ItbnH5+eESDr//yX9puozYOzzS
8VU68+dI3f3uspXXn4E+CYaGb8We+pXUdrG8jlr2AKZcK9CO1t5s4SMw8lpRN96c
ijQTdQgqrZch9tqe2gc9Vj/WM+JRETrTudCrI0BK9pW7Flhk8wKaA6dQX9f4FMuI
cz9gyRV6pXBMBW2Ry+wzrcHUd17zHSa/Aau6H0OM8p9A8lHRjXSH/OoZ0rd9xvhl
KRhaqKR9SbLly55Zc5xfjzncL8DfgrOqMqV9tIj2o1AxxtSjyQeS0/wLp+D0x/Wd
MO/iI3dp32Ojuc2g+YsDzcFPlvwyZfX4xsAbAOPHTgdfoNQXwFzCfQxqCtr3ztbe
oME0zVWsuZKGHsuyuOWRFkzq9r/0wqZ6wP4V0p0Ak6snp9/fZUDVJH7D4pJOswdo
MyQ8Gd/B+zCu3e0ilApquLwGGTplAuzdD3NIb+wYpou47UC/htB2sRcS8Bls0AV9
EvKzNvi9c/0PyZowEUDonLNLrTiPoMcDbFYA+ZdvwKJoizEjLUBgQvta1556K6vO
3ORmhdw3NwnpqtQozudqsvwGAJXLtwrojTZuAdAer6cn0Qo8bla29i8RY8xHeAb0
9TOPJfbkK0KzhkIkFsuxcP8jr8ywUU3/Byc2SzLkI/5L5UaSiBVUpO+W7H/kPb7w
Oda6O6QK6FpOBXTZsp15bVD3OJdAh9wF0rWtCDTiY6vr0/EjDnO3DoLtTE2flHCX
R+zl87M7aCQzTbNrRDOBofDJtiFCczJfEN83CXm84kzefaumjHNi75w8O227VF/f
JAAfSya3GPezhQTD7n0bwp5lpRk7XKgUmT1gNsb/ABLVNsqRh9uqvwIZ4DxjsJw9
0t5vytDfcOHkqJpwe+vZbAEfP488CxH2MJoPQZVCJB/AAxK19Ou6Ea7m3xDVxTjY
f5CEmLkbxt/n4bk9Jr0WRK8fAaeoegpR7SjDrCTbIryt9yvqF3n8hLpNUrK24njz
nUr2XF/aQJawDOcYvG77G1VrmP7OsyobEElHuCbKfIhzxGqYh9TuOLxyZAw1yA4y
97S+UmtmThAl9V13avrna3iqJRFRy/9/JOdaiTInBWBfXerlywjjuXDbg16tJMzf
Fzv5RqEgMLxnYezmzJsE016Bxr/XfQwnhMmSkyl08GukWyLqpGdgrfjC8HErUvoe
6LkvP8Cu95PT22geWFL5r+YxEpXnDddNd1SUNgEjfhyEbTn4bD6GLJrIWxz04VB7
sHzfB/QyCqeC/GjHIlLDbDkUQsqrK+IA1DLGIablTbEwVOgGyNqjKAG307gZJM5e
dvwMpDli3YuI07oKpk5JzUUdp4Aqcr0shPm/0fLHeZPDh4LO3RIe0YweCQ0Cu6kx
AMJDR9ZZC1Q302HWgCs15GWqjAm0B5YLVoecfeS640/5odjE7u0UMe0xXBrZeciW
xqJr5xMK7FIXUj8yYgx3PL74Nuah/mzwvzm8zKZw+2TaT3xDt5VoSTM7vkYPb8hx
o6//l6siIqOo0UFm31ZfKO7BmG6JcWeV7ltIfrQ6sZC9X8eHNEsEYOBOj64wH4sp
FDeEhijMGa+7Tsmsrwugx4aek33wDWVVpvB0bKhitEldYeQD8nql81a8fjEaC2y3
/3aVVjIEGpibN1hhBFSvnyO2UCKbjljHJuJB8zvkzsMxdMoGrFur3mZ2TDqYVd9O
pg7CHA/DF97HUvVyfusr1tTracNYms7EHMqOby56ko3/NeiECfJZ3aX4PvoWYM/y
CEQtyl4tDgOvNWR6CGmkptMGvdCPPqAIzck+65ni+iX0OFRCFRS25j/96M7WzFOP
TBToR+Bjtp5ZhdAMTUO0P2xL+xJE3oGp0frI6C6vysYKrJKVTmvnANUlkpPYpeDL
//lUD91cZM1hYPSt20mxbDQSs/8SV0y7px+ucZ2efgCJdDETKVqPrSPhiKjnB68y
votpuIec1cfYy806j4C5JKnMxPK8ejfX+UIq0PZJw/FeMiz7nd63kVesFiTVNzrI
TXLjfUGKc739DeSzXrpd1/SnmtQDVljsQ+a02m+c3qC6gCih4D068QaC5l7sT4oN
rpk1gWwn1supHQ6+v9BFrjF9WR+rigPmCuKBh6JyYynm7ZJSuhD4gWQ5mCMNhhi0
xRY9YeCTG7PKcSMGML8vGL/BJFHbGl++gY9vvXy7G7qcfMaao5Hge5BD8cT2fa+3
MJJQaUxtXYZbknBTGTJM5uoa6j4GNmKEJNF0Mj6n3vofzJ310KDalpVKPPbtub4S
qVQFEVjvnctDZDNG9Y1Kg+weATgtQ3WHFtuEmL4o9kZA84zejQ9rtkaAOpQKj9xX
yvkor/6UGAVoTNLUaDvWsNezuUaPdp2MDV2S6B5qU0grqoSJYptH4oVReKjhDfRM
LuE6EYnVXFx76rxM76/ErWUzBJq2HQsLp28457j6bGBt6nLPei8M85zBhJ7kz5D6
2Cic8MHFsJTIkylMQklRCPw2pvYXiOsxdTF0mhmzGEkcZFv/LPyPBsffMDxNI3eo
OjzROO1XyeYtZpQ7yQR+qCTOI5/YxoVU5QJ/I5CWLcceitUFNZALGTk/MINdkgX1
J78Vd3VNNn3dMA3tJkcRTJDLDe5ytw3ySnoBEN9UxBYGRKTxuF0mQdyixjx/ijiw
ErtdavIUzcfM54tQnRj3ymuXAYjh2rAAjrg7HCm2xJRKViQRH2DhMm61hddiSbtV
dX8lIQzev4UoigTf2n6DnppHZoYOVobdZ38Qog27GmIPWXoedwMolhD2xc1rCb6b
UzieXmJz7vidqmfBjXQEASL4IyMSKPMvTptwppxqxUlAOxNtvd4qskZU0SuaH1sv
y/5QvDyJ7WxTKbEdGClIsYFN13AXpkptFHfDDRxiZta8regeTdPxaD3BTPVymkkd
V4ntpO50q4BivZrlit1/XhBAzdO3qv0XZmdKg+rIx5tO5jTFFV/bS7vXAbpn8Htw
Bn+8DsfPN28Hp4i8j25ve4ZIi5y0bMDELrVnDAu6wNAd5FjC4MdD2u7EAS3J6Y52
QcJKx3zccpmKMggw96sTQHzJFvt9CZMO0pb5aTGoOt1yTsa6PoQxxtqxvwV1EsB7
8YkhRXt67ztrhZEm46duM8364YRZneVAgx573zkWHY6nzsTlcGIBTGw3N+b8xaG0
z0cF5eTCtnyYibDAYPt9lkweA5yy8FI2df4kfljqVEPamLEyaz5J/cU/yYgWEefW
WqpjNeYFA3QzLuQeDz1TriR5tZUKA+WGCIbxX7Uv+5ZPHWGrqa0vEMEuEeLWe4SH
kpIxW74cYGVcMGwO3/DQdbgoVzHP/Nz+cNlxBtoiG7YqCTiXVgi8Gk6E6YwIFP4p
QeLqANvRM2Rj4Srji8ZysEjLRz3D3zA9B5Z4KRwm+xmH85qMjDUmHf3rhYz9Iqvu
v9L3Bwnt5VUQMwoEgdHcoTU1nXtOgFx0+jzOQFl/eVa+kOcFPc/0nlH4SMN9LTJO
jkryjsEAnPpQ9aw+E+HfF3aDWiGwBIuYUV6A3I+aWfvBCNM0iJ17jce/95MkjCpF
lpOLljupYQh1GJkSiPB2CCrBLUzMuY9qn96UCMQB7i1j2NUxGMjzx1W3HrTKprRe
sOJt01LHonB89O+7Yp/11rVRERHWOs4neiTrfYv2ZGbJaYWh3htX91T+TL1iQNxT
eR+m3u1kGVmvMv5ako5t94aUM9bFgZ3Is8pY3oNzfexITADwnnVfKopDSgDG4Jb3
6imbgz3+T4l+EsbyLdIbenoZZsIS8KHaPjIjO7PWobVv3+PvYjVSTwTf5NRxo6j0
sZNUTlLRYdU8VN2xNCzXuJW0ZQxARTrMhKC4IU82xh957vnuZ06xOl0WUTwYmcWe
qsCpucxYeBee5EDYiamdN0Uydz4ItE7RrRZEIXq2kCHECOXhA9Pg34tFA8HLYOT/
xaW0FL3n9kejjstIvng2zHJ78yPQ258QnW2VNNdX42/7d0UN69W9Dmpih0/FGHuI
C97zssQZyxoDSqxEKSGAWGd8sVIFpmKSSUwwKMnNDTTJ2k09O37cr9nkr8lGKfON
aG0a/Fqb6qyXe7nTutmGTblRw6Jwrel/CE6Z6vJUN2S3VEfp0rrChSmA6DASXp34
0e1zwF3DG0Qs7SG7uPlsfuw2OS/VsrKxXIyUT/MzQuVt1tjLw78UAg/3EeVFc3YT
SRPQihMXzqGURYYOQfwfdsBB4sXAPjiS/ZkgnFYitimQUoReWG00PQrBnFa8/qvK
MuLLmkSa2q8hrPiQiKXZS02HAhrdgNKs4Qd5gNN6fxFh2vJt58ZXUG+sN9KTOWlS
SfK4LHTyqxtkLsWOwBmxV3m1s3bYnxqxRnJxvGbcwrONRdhNmLwr+wisGxnXbxcC
dhwsLipw3yX6cNQEr+BjBf4PwLzcce1rtfqg0ME4ZhrDp54uvfhvuOskqlqMecyb
C9BdezW3chS6hiAVCpSEhMjo8Yi4poJnpDs/ZnPLpqXwoSNsrrIgbczJj97oD2gs
hT8NFg9YCCX+kb0BFJqCa4GxbZBwirAxRAykol3FbAuZ/W1hDdSJ+sI3cGDEHB+J
HwNHn57i/gOwPKtOroiaQjiYG9gRGUduhFN0xMJpIpn8vz75+IpC3BOYdnf4eDEe
027qQrvapzCloP86XC1nt62meH90UaCVlNaBS72SamypRJU/pvJ5/FD9KpzByvLH
WQ4BUmtBzCy6MATHvmz6kDREMDA5wG1cdCIIz7P2Q+KVSMUXroVyAbDX2wTZXC7R
eQ8pLACIE783jSwGUrl5m4KbFphhXCtKGYz+zstuJRsQvO9eJG18Vt1DdoZoKRW2
jE1TndASJdyw3jGUACYHKlOjlJIYaz6fRiSDNNi5/k6BGOFUSrD5Lx1NRTJlzYCB
DEjTwGmdRAYldTAhiTMIEoLrc2LP6j/8SbsFGn7zi0qJfJxDSHq0hXyWaozvgDcd
zhKE+NwaIqKsTdtZ1lryp15zexvdQsqkg5K4E7sliu6u0azFBLx8VWFbwU2Ka/dH
tAI0qjx3k1XMvS1ws7FItTUs1jxOd0NfP5n2oSTZed6dFLi4m10jWdqhdHb2FJxc
MmZuOFnd+6iO0CXgCzfGL/7RYXMveS0hMet8QoPJfdILaJaj99ED5YJTucEF/+6w
vXqiBdZVszR1mGKdhRlzymeoUKaAJAGcSNvTQvFCCHtuq8BzzworNmwtod0QNSC3
+MeVDP7IMrYH07Xs3LYDhqAyXTeOTwc+rpgG2cyjQGoWyPZ8FVZ7qBLBCrjmOVd2
hbChrrI4BhafK++/lKh3MEcM64wz6NxJib1uxA8NVbZx0IQ3fxaez6bvKkaCcHwz
18hUOVzzOQRcug4tWUAEBEn04Mthv37bFIBVceEikIAC+nvRM67P6O1inD9waRGu
t7hTq9ucplHtAFq+E9bxpVJ13fSY8BN0q9JRrbT05xE8k8ATaWcjrg3sE+mVxfXC
FUIsPAQdvf5/0nCZ9Vqf9UJHYXMTjNzu1hAZQ+t6sP7KAJm37seLuAD9cT7C2R73
HZVK4zXgReU6573msnN4JtSZ9hK0P5v19DTq6Wz9vZAVxhJZcc6K9QEU8I0Ppcjq
UOU/8VuQ2GHNmU8/+mv939TRYiLRxdUk9rxxXUCcFsVnJQQRB10YyUsCUTaSu2ZP
5rkrF7lTlRUi9XH6KiioKflAMvvGom5JDF7Lz28Ylh/i6WZG8V4ioMWH3rJMW1Zh
JRJOt80RNJVoNR/oRN6uZE/OMbtdGChnlHMiBWI0RIyU/bYEr7OcjrekPSYCcgic
D1wZ1okrsz4YoZLJhkOpibxB/bHezu6UtDidG0gaJNCzeBQ0aM+6CJ4yfmYk2nTe
Hgf2zvq0pbGImhP0Fqu9ZsgnGDqERGPyhxC+qjIFpAbNrUNh7gwopr83nNbV9T5E
AiMSN0JWaoi9yU9lknC5xzKaDsZMImhiyiqsWvEbmj6JFc/0v53jo+w9Xq30KZAZ
L1wd/sBkEu3GqagqnEnj1advMiAbHdgU0LYRmpNyhBVye3GFaL36HDCuv0bwi5nV
YOecfW0WaBLz5X/5iC0SI2v8KwDOw+KTGaYOSFebWWBGCedRJjic6IlB1IOhaXJI
vNACZJbs9BPRsLuiVSgYXXGX94WKYHf8LiqN+B6kXOj3CFQdU8M4K/wr+8cKtQH7
16tIDaPpNnrrhK5fCGN/QxxkX8pfxhE888DFFwE2TuXytSrbscoSYkKOAaWBDPAS
pB57ryiryfbc/p+paQ1zEhsbfoc1NYk/odDU505rgH6VPiBkjpcSYQpG3+HlwEXu
X9OtjmiUfszB0jQzzacIJ2ZcpesIFNmEUSjjG7da+6PPrOI7hlNAxqAnVfePmihb
oFzAeRt9vV+krRV8Io33UWymk8rJbqKwZx6HDWx2Vo1vSrqnyDNgywUbhumd9UKE
iNzoKBYfmkO2npnbn/5opEj7yTxZcO9j8+eKHAO7TDWTiLhfzsHpnew/ExsozHPL
KnmRYIN32aoeLpGEk6fu6OgznpLv7oK+LQPh2TuvX7gwWGqBCycnKrdgOcvQOzsz
Zst7MHYlD/ITydj/j7DkicW/qoo3iIoc2s5WatnWknnCrpZtAgc/yfjvRM1DYzC7
tecS8Qvjr77S8UPg5Ko/4AffJ87ScRaimGobmRzz9/gu4B1Xn4QLMYCHMEUq/qL9
NqK3H8QzGuYJ8aQgPuj9mhyzkVzxS9pmBFvdnweLlBpc9eBSijZaaimJOqOf4pE0
BG5yrgUMgUHnOBOlXWk0Ba+QJyDt+i6oib7ua/znv5uQUmPzAeIXiN7dRhvzTkBo
+/agzGPqCzq3AJNs0jByH5qfXtqs9jfaJ2uoXZONIpYceGMEUTR/4JU7LWBtVgJi
xpJsBjjjPZjREzwG+gjU9Y62T5rctHrQoCAe4ZS9JOdyiyvi6uAv7+OBglUd5Iw7
sJE/s3IcEBLn+x3lBWAR+Gv2KaIxmuTDYsXTCD8SAxx245eKYKKWQvrVP7R+udEH
S+JoiFwoJfNlwVjkh7BWcaD3gCCw1rPoziWas/oKXn1ft3pMuMjyJ3GoaTULju2R
xPoBS+tUJAs7kDVPVAyGfATZISswA/2KdWmHD5Yn0CwOT0p1tWf8L88jg8Gsjyb7
OoImjK80rpby2S0HEhCgAQPrqps/hc5ufpLrYDn5XSNJVbDY3LoO23gjBxL6w4KS
TSFp7ALF/6Yu/SRI6s2r2PIIl4J9p7laoaa42clgS/z+2a5TplPO+yX1ndUGuYEf
ytQGlWg5v3ro0W58uL+atFCekN6TMFO/E0sIsgKiLl+gUx+z1m5C3xv5meVl2lNg
jqaadgv0jie8cep6i6A09KsjJqupgUtYkPkUPGCywGs62BpKernFXcWjMpWUvuqt
XO9cEnpQgU20v6sMOCPNIXjZffKx5ulzdsa42XFlpB7IDW+hWEQW26FXAyUlEm6F
nrid2v+to4zMR3+qnqAv0oTatXFS/z4GFs4jsopPag4OvDueHVDCvaZKlKBYip0j
CrdHkgy0N9kDaaotqcOC1xKCeCMLbxg2O24W2LxwbpGWrubGj/9GcJfibfBJuom8
l+EufSuhMB86VA5imkkGRuwCNu2LJe+2Oqt6YJCRp8VShymvMCl48MfL/RNDuSHh
XTpYDkY8usZG1yqQbmpidkSIcBZNyRfE9Cv7fJa2Y4C/m0oXemN7wpiKyNRBZkEX
SygLriVf21aDo4BXp0g4Kub4vhoCiELIwbHWq9Wy6kuJcUBqhYrwV8pbohFOZpnE
FKl0WW1VmAhaSqoFUEz+hD0aseg5KKFIgRxFoGhflzvywheeHvL/XGqgp5HzULw/
HHu4v+lRXFUoH4UIz0acFR+5z5Jlew5BlanB5YCLUvmTELJaojCQcNmO7rxHhDlp
I8RpoWMrDCHyZhcKtvhqLomqcEPFXe4EoOk+NZa25yT0tti8hgPbGnyUQfNuFeG7
LjhaVQ0QusFGZacdko4+nsfR/fZQULeMrMkOBce01Ov2pe5GpW0FDMNaLHvMWVbP
jRklEp46yxn30cILZY+yNdHCaOp3uctVRvgDcy70t4ZjkD9rU24LUGtTO6dEtjwu
qZwbYrm0XQ6ecG54EvmTkWJRZo1rMmmZMQ0gGTzkkH3Pzc92GQ9HG0c0XVn2TMsu
srwTxEvm0FIe6f08JrGFw+anuudxTnGticAhLeQsrCZoiFc8iskhcIkfJHfMyt/2
Ou1E73ns4nHEb6olXHyJCbSYTAHxKOzxxuowL7J+sfg+aBx4MzDxWPChFbAaCjAn
4CoqBGqvizAcL8+sertMvn9QuSH4ZwryDyOT8tzCOB+IoVGN3AVV6ZUIibkkxdTI
36oJlXsJBHJUibHNMlTxEZRaGRMdQaKuWvTy7ZIPgRHZrFHv+dejKHpsT4eSn4U9
asl6kzhbAtC+ozPo2xdE7PuK5PiPm3V/4OczLNlq3r4XcqklUt5h/K1pQb40VM2C
yhB7DfRz6HcFbFdDEfDTUme6Yh3Mk3hrwYTwbYGFai+S73uE+bWCA0Gx8SZnIPIU
eVGLmvm2rGOz8lp4q+5SbYJ4arGnnREzDa6ZgFn/4S1SR38K/tXq4Ptcw+B8Yi6O
562vRJFqJ0ghp77iBK2berLq5Y+FaF2pXaMDDsgciNzx32ppaeEdHWYGBQzWHQ3c
ws1uqUL0IxtyKtgtuzhf3Xx1J/QcaGtaroGbpZPXUzWxp6m1oXKnUWBcEGxn7xZ2
thIu3oE0He1sE9flgwFBt3MwppHhOsGOrdgCjVnl5qg3DoOKDfQOOdUtS/3NOTaz
640wEGtmYTfhyOgD6nDeBCC9hiRVJVjZOOW3rBBwvjZ7/5zBQ0sgFgQjxkDdjbYI
c0QtnJ8FQ7eMrKkRlJKbja3vQwem3X26uM0qLc/4yuLr8tU4SmOw1GUH7vczun/e
La6ZW3QcU1nIjawVMLmltaBQ14RnQEGV5ShXS/rmKl99ZcYtU51xsg3U4Zk3KkhJ
m6c+DwiWTr8ZQv1WsU3q7q+n2ZYKJ92GkH+EtcVWA+WnjLMtrkxFacNPqqcNehES
ilRQ+JX3yuQWUK44/azrrHfgQ9osyGeWwrpZQmQtL5IOE8NbL9R9RPBsz1aDeXXZ
62Hlo0Wp6yiYjot7zjMeNWaNtFYLP414yRrZaWIhO6T9XX38Z4ZTyke8fMK/52kU
yQ4ndspKxtVwcDuLZkyTqsFnWOYTbEQw+Q2sSMbiRc05QoySw9TUzGVs++5J32WQ
Q1LYQZic6FOj4LWcRGa5Neh1/cKjNRBEzlmVpSMsv9KmOuoWh+XQfM9+BklYghk6
CKnWoizVGo89kWNHvmZh69ir+OpS+IoRRs/1NbcM2u5L9Rcm4uLr28DSvr6nrA/x
wNwJHqt/9NR/xX/8/Bel2Z9J0RpkYm97zy7IZxqfdNzPGDFRsNf4NjD/i/ccAS86
k+9BA3tdlDSI6bwkzvygVPg6T2OCgGGdl1X6t/Y9HEiopQHnVqUdb1MK3mMkizKs
xRZgRnM9aFL4qMuwNmzAxUFhOPBGjbRscIVc13CYCGm3BFLin5HJ1+BHQzp8ImYE
EC71M+x2rSgX3XV6A6yHFLDXQx4/ie68MxUuwcYPupNU/JgZYr143G7lXCJ+K1tx
tT6H9nqxX9CH9IAljzRDjRn9YXU6kIggI5pGKlf6R3lw45P3rYC7gv8M9MVyhuHs
DH+utrgwY7wPDigLT+qpEiei2WKxxx+zohoMrVeVD7CZbWMUwnSBHPkMLiQgp2Tl
9YfYTzIPPkcSLc5pySOZeFuUt1JTl7Gx5pR21DCdzLRGCM7ubHmZoCf6dPnz1AlP
kvlOHg8o30Vh4I09JucKXhP+9EvAAcCM/bdlpNeZM2XEatg8Rhaw9nvmbbCDPlVo
+k4Wl3gEuNGApmS4BHiV9ShGQr8wSaheD7b1q7ZMNQyexxl+0b7muLJIw/ZKTMHg
7NsdsoTOInGTFQxDPn3M8K727OUDEYT0h44EJqfs7BPfUpUVEuumAR0PeOaPfM+j
6ez5jv5KYxSBTtn6YsDdxv0TK02l3hwJW90KVYxH87tPhkp8c4Y8XusGezgLR3K0
dY9BT6LEyRUADiQbSPVR1yVJKRxWLPLa83JhtT6aJRQJgHe1ZJzVKZpdkvhemUgS
pTxRaBMyWIhofHiWKx6YJ9UQbuADxqQkNQ3WwwJ8Y5Qu3hWZbaMArp63L3+WypHI
xUHYvg3NdEG49XNuV9pwyzo1nUnuQYv97b2C8PyVWnDIe+zHMJ142aHGonHc8l4h
b/bEOalyZDaz8JEXbPBs1CrR2I7sWJIPEkTN0TVkX6cF28pqJgAm2qEvShUnyYoz
UuiO8BH6wI3c5H6FapYOsqfcwGF3PrXIVp2Wr2KQbz8FepFALARp7WU3cLho9OjK
hIo3ZO0KOSNLbNcFwRXeOsGt5APuToJAngpL9N336Eq7wM+uGLmXvYZpE/GXyB2z
AVTS1PkRiALIHnwnHrCjP44VjnBYLaFDgGuwbPatXETTb2oLIkMPseUdIklxn25h
knukZp9vtyXSl/iJWDOMioTbqve0uQWNOUBHz8mRvhIh50PuhF5OUM4gD439F6Jc
poft3XkGHDhnlo5tAEtowyU8CcuQkcHbDQs9lyJqK8h0PiUrK9Dr/giLCGyJP4e3
hHvIrY18Dl9DHWYHJU3mJzbHFiNLDJPJKEMmRpr2CPnU3kFMEXmSUpcjNPUZBiZR
0glWHgoSPtBmI5jsGjjXDwlQlLTeOjD8aIA14g2ECjvzgdyoFIFKNpt0nas8cKfY
ZDVZWAlk6eEqFsrzNtUFlcHO9khy5fmNvih4iBAtdc+SrwcIUarrVWidfHi2hnb/
ZZESWlrzzaRFwsGx33fiodWi3An9TFDfLYX4u/y+nDlyUYo4ek6LRZEv3P5zJNIo
bEATTp0uD1sD13KOPsmeAGZbhzYhp4Esnvfhlx/xk8nUjlp5hQD1bPeVqY3LeebG
RsR+0Ele3wsyyOM2KanxcysAQrIC+3mrRX/nYUqez6k9T+nhEAOwzBgkYmq4efpx
+eAdR+5FKboIF2gLpNKmIFGrmLBIrubqAkXlc85r+DB4BEHVWb+T+2z1IjyPSG2I
zjiiHqGJRH+Ovww9mKcjR204GGCSi9jCi1W+VJ3oHnXURvP90nySJl3S/xgCK0OE
VfU3YVP0ZBCEZ5gth4Zb9M+4N8jUvZjc0rckuzgy9SEf8z5vl9lfCGlC0XATAHvo
vscl61rzKUvk3x+RCsNaM+kUqm++ma62ynu2jdAT3mseKzhv2iyw+s93EBkiu1o2
M3y//Dy1JJYG2H7z+ppJoyI7c4ogMLBkn9Z9S74WTDKIfBp8y15tt3F0IENNcyTQ
PqML8ifMpnzk8UqFGIT0QXKEHfNWbbNR0jvmODD4LqsoCFOYygR2FldH2LKqlNkX
V8XOgmqZvI9wXkZdRqALVNh6ggMa4ahv3XT7mct1xx4cW8TQ/qzxrH3OLlJHXyzc
v2zv5U80bV1EmCTxt/W3T+9pXRIdxmC6//mxeiGfc75u49hEoVDC80BQNqOp094x
0o26Rtc6iAMLHGlf5ILZnU7rIFxIEJtsq0q+YvYiYq2g4ojuVaveHpxB7vCX2GvC
4otXfjcCtqU4ZxZwoZlsL9J/KucRYodPcQMPVHb1jkUYGcu0E3A0rzCMRtm/KLYd
D2GCEsvMMchvduxS05PXTl4jiEyVAfETUXyfrUZ7V4K1GYGs8ESDzFiOeTsh27Bu
zdk6SIym1ut7JYOOoN6vBDvQErdKwD5jWnQYajN5JvdxMpjo2j6p+3pcRrCWrm/b
xhKkiN40693pQIlRmL7CIcHJDZg/0U0WPk8hghSLOoeAsLsWE5KsVC68oumItpr3
pPNlZ7i0ipv5udswkR9YxHIwQwOg9GdECV6jlWL6NeUwagmBK+MpKXOH5YyGxGyG
wwWS5xif4Y4NDFMdH9Y0q0Xz+qFcCNF7p2Tr3aQqxuMPd7R8y2F5vkpuJ3tPwHbv
Lwx3M/e61T4mcbkr7DORDMsurCa11xApF6pF96rmwTSzV5fZI7UQXgLSKdmR4kmr
CuGx+7Tcl/KsXJ5pd0JQ9R8urqgdFt317wzzGGwIMV2Eo7wvMRwTEl11i4K9ah7w
DO7iIZYWc/ktJ+lelArh1Fk/lLdCcv00kd0yWDF37FAAueXYXa1c1UVH2OQYFEAG
lBzg+pO0gBe4u+clAlSAgUuzYFJ7FwEKOC+J25YD60LPdqS7UDTiT+Lo1UyR3BLN
UA+7eYA3I1JfHmXWbGpYPorH4PAWRLUhakDXXrYAqBYaN2mjny1FrKbI5XI3M0AM
Qt0UhWZZ5BCI2C/5r5N8B7vzGC04msAOxw3InebEQ3S4E13VuASQVz8wRZ6aDcF2
JCvmWXPWg0ZnUX7xzxUjVeRE7J6Ur3qJgShl6RLzkiuDlqMI7RXY/krBFN/as69r
/1x/UWIN6v1TsXVr3wF0995Yf8ZTENExunwi96klOt2hFKjQkB86ljEpyXfSXPDS
VqqqojvmYQkUg5v1xCAO+uMLzrwvmHfmC9hG/BLzKQp2EXfe02anVcF2W9t9mHMb
dcIj7pna16G9TLAO7MshWbLbVEOwYbP3yhgzKL68abzA2BqlenyAe6ameHmAR/ee
JslpBL2OXblRlq8hLzKrCyeJIWDfH5ZrGtFzZKPtQNTXGbv6nwSVoDJKHhh65rFM
KaN9qtMJBgK3dO3vq96T/cIBP3GAOcoICDKzfGoYfWXrogkKVIQlmLoBPLfX4dw9
6CMXCO2FSOetERQfzY0jrPcaQmQaEe/hQqCywUGCkHRwI/yz0RU76Eurmd7wK58e
XrWzDyyZOFQICPqQwGQNQHUkqOIwQKBXgOgdAYa/Gp0/EJa/NI9ir6KiR6/TSYRS
oYIKsapMn666vwHgf12AI7MJpWqMQrW1NhI5N2zKrgwK7Nf2xHSDud9u4mOVXnDQ
0fuOgWSgwx0W2gjOyCbNZDNmNvC13GO7F0x/Ulh5ShYVhQhGx5Ka1x2sL+igVXkU
RaEAX2NZ1uaXlXkoU7cxD2YPbGCGU99g1qNF9phVWvTPtFL5Ien6N4j8q/slqFKg
cif8lGk1bwNRuTdzKUOz5tkTT0QUpOhrxFXwFdBFuuF17P7QaCuOpOAm4KvuGP8T
2YWh5YikerRzBG4T4VUVrD0L8xq8OgUGYfnPv+7rYzsZ0NVgE55xlqnin3iFNclv
l+xWzOg/INCfb070WWniGNx/5Z0v3mDaKFHQuwMhGZI8BHI59Dj9xTYbL8inxxni
Ni5lCcYJPEf+S0tQbVlQKmatWzbN0+bm7MVoKHVtGwOGlNbvf15C0ZctvhCkvYsG
twPOIgFgxK66/K6BPO1g69IYW5d887tHoSDwbJmHhILUmfBRqWOk/QlS94F7SFam
iiwb8pxLdPb1mQ+FCggA9hYMg9PgQjEW8oKv9qWWhWpQvF0umFpnV43NKfkj7/JB
F1zhjYzKeDAhoPU2XJbT4q1bNqIXrm2/2WctMRkXUarpaxHDRz3aN3vCM5olagFf
qVcRDCOVRsJv63PJ/j88PWQOLxfOlubPLNAzT61VfClEycMCD1C41/zVdAxHBN8N
0nfkXVPxFkaul0UIL4pO1Kun8Oaotv3bKp+nOsZ018owdgzGljBshnjgYAHwkNxF
pA4pJemUog1E9mPODCV5WOv0LNKVuPJhLxNary9tpkP9l/0eipKru/Y5bnrux1Bi
p8AqId6cQZZtyR9ZlQ43P01Bslwv97fKa6ITyTH+Bum/plYeKLZZVKkDcgmt2m3q
36Eg196Icfmtq+L7PDZWxJIUtzEk8skpIq7bYdUyYnYfkJqWUNyKr7cuJIY8wlHx
RS/ldp+dbI8wC7RGelvYqB8lGB3m/P9gvw0ZMwqvGvIuOTxzUnXpPZk3ZH4zAljJ
YwN541yAxdIl7KllJENDH8rRBE8JHL7ISTGi8fyNt6IG2Jjkxl/ahRZhBO7Hrgfr
ZeYq8f5UNrJU54oQmt6tRDXrRrU1LlRmO66WnWpYqWi3uA0eK0Ban0yR/1pzG30G
6zZJFPpe7pEAywh8AL50QBizn+vnSJ0YyjnbLFej1O6bKLCU9JFnIlLU9ADddKkL
d+AVYCJ2nHES49FNG9HVfc7Mgw9qqIYMe46GAJ0l6TwPjGGyIXnkAn34ur3f1vhq
MiOJwRrVnDnicvC2rbNfDUWx/9Y9BN1PHgrmZNimwXCHbP4ZiUNS8wqF8fbhR3A3
2sy4JI5ON/mkGnmyoFjsjxwSwi9jr3MQy64lLNAe9fWkUOiX3dqL7q2esZVsYmqy
icKH9hId00ukcwP/olfXHM0NtTofR/N9yGHrVuYSKETQLABcUaihYjK/3UVGDpI3
me1xC3VKwYXWa5H3dCCoH//rb71uEJtp1Kw0R3Umk2KDuyFgG2fWSb4IMX7k0Dud
kVbbyaJuSdWOXTO5jMMVN8Mr0QTV8GHoBQwmGdKgKBgEonCUJAYAi3vFb42d2JQ6
ekuQ/afSC5b0/Uhi5yzeqJjghucwkcWzpZ7vxaISX3CQk2L2IEv66WfpW+9JzHlR
ae6ViRKgtF3KZQ9scxAerHtHlosw97+sOupLogyVVKgm5C1ZxdnpqvGcs1U5AA85
shICxoaypkRX8KHK3pydnlq6k1m130QqJo+SHq+1hBpCDj1Ei525LOSuS0g5M5fP
vEHRJ+18AiG2R+9kNT3fLAuIyCcVzRjtS8uOwJS59xxGQkLHrJ4yByLLnFKWq6kn
nn4WiDmiyAb3PF5hzdTC/5oZzjEpvJuoyRkdzU+MMLQngWG2+E+8mpH7vUrGv7Om
Npkrvb+1rx/wcutC1X9tgFtoULe3R0mblFgW0vl8HYhCo7k9jrWxD9/s34qVF/j8
oqeM5res3z7Q0sVqc87Y/A0/an5TwUbNgIY5+Y6KsNhDdF+oGJtQ1u809ai7G8BI
x5d2DNmS+2yPoYkUR9V4SdGrmjLQ3KxbEr4FVLn1nqBusaphx+Tgtspe+3rqibMN
nb/RqroR1F6wXS7FnEGeMtWy5JhRxNAX55A373KxUO63DZ5LTSqEGhX33kMUwcD6
DomkJjLRrI2lV4aJZwGsNiD1B5Gg5+n6HMhD7kdOWA0BlZvk7oNmXaPyj7ImKVZ4
/Oy+TssrBIOLz3SpNnPZ9Bs2/W5Pc3ORxVNei5x6MNrdZm++IHMORqfxhz04uu6g
/6qDawrf1Jo0r+c7JiR06WWPXZu5ilzAw91egkseYvqDLK35apCFNOcGwPrM+cXB
6dysqmldT+mZ9ml4WUSKo0rtlCT5BQr9Z8ustJpk3gUv2fzDh5s+dlRlnneJfeLS
JejvLRgBNzUZM88VqwRaIK6itPmO9rhOIWcHjTXocDl7VUjYsSa5JoKjuW2F5U4x
5l6tEoa3E2uM8LPWy77AYG3UYmlg0jmKHcQ1PJoJB1Cllnilxtbd6QBkLZTxRgac
+1EEYTCIUYGpZtK2wq1IiPj6ipRY5vniEsgzqVm3mkMLBY4xla16RuQ3JbqG4rwI
v/+FCS/kgpt51h6z7BbcHIPw9Oh3dsxSBILsodl9rbQJ1r6L7qe5wxXbVIONG7ON
1rBQDq4jPmeySxsemLIMQSmEj7YituedYP1isvZbq4yVuYI/u95QQQx6hnmB2z0c
ohSu0pzo5FNZz5d78BrPwesTgH44EuReV7y5e3ISNMrnBX/oCba4IeaUVb2pjsWq
Q1DZPQez170uaO5bX3h+HwU7zgU4aIBQxsX1FcOzfeEcM+Q+L+zgieBZBWGmh3Tw
7VDxdojvUzZSg9pYpbrSGXeqR1ExwWZtwonh/CwV5CT71z/4KbXqETHh/T3LInMZ
jDZcrT+F0+ozVejyus2Nn9f5jfQNABPzEGvBGjliOBCVl5hgR+5mR7nJ6JpKEwa0
ujaQ+NomD/vVKtrps9EbP9uFM8E1+GLcnw9ETJlfPk9IKtSVpIPkFxOc0p9KDROb
05KOfqXIJH77TnqDwPQrw+xgGjojUrL7Pn/aOFEuRvDAX5IJ53zUQrSBGtuWh60c
DDCp8BTaHZbRx2MD1ouk5FJESvTyS7ap5StobAz7+yyVugfZUNOBS6X8oRLp8/SB
ParoAAVd6l5yTbnyh3UxA8Etuao1d2agseNRjQbb3qE9K6mt58qx42v5g2vlbiqW
idrIMLTT2yh5a0RASb9rgT8r/FRLefk9QBkI5xyF2ZnSVIUz6epUTQHxGwnr67fQ
iccaw1fRHl7L7yBVG9kyy2lLesc4h5WyP39vYcDmyKSMpHfysUSeNMiCIH+BUFGu
hgBkPzMRi799ZnSpxBg/z4B4cBEY9o+uimv8wrTdbi4bG9mdMo14kqrR1Um2vC+R
rLF/5CFOxqGUgDJ0etuKM2H/JHSECyiJjMZ81zxh+nPMrRwn7eJXI1mtjKAhyLi9
Wq6mxMu1Zurr8h2m4fEaFjW7Fw7CHThRxRtxNeHckT1zgkZNOX/FvK/D/PcWnOaj
F6NjpY+USfpHDH3fsgrvBjSV9v/XPn+0KpUcTHu9mSap5AT4+tg+qyXiLFDexGJd
RTd6VKX1MJoaAq6yoXdKbzFCle+9d+5WKj6DaG+e6h2/nYgjWPfA7QTE2rY7aVlx
9zd9O9Y7VFx7lnJmHrHlUMh1ZZnovik8GvYNeA6q/JmBlQpDRusYXj0znShsR1EX
+nJ5VuiPC7iPLq4Y+RDdCsk0aW/CkRG2L96jFhV1yeqk//Prw/6BUkmAix5oG6F3
rS/CR2tMjSoBrZKhPUhsLczI9u69mV8Sh25/G4vkSLJU7yEEi9bYBiAy+vwipwyq
+eMitg3e+RKPiJ7knlqIMO2MgK5P1ONBdYgusMPeGg26DVTfvvcT5BjyTq4TTnOE
NSCYJPXvVaOHrJd/HqZvVhdULCDAYwl+rXpnez3DPXtaouOrp91/8PFhCUHi49e/
VMGx0hOqgfaauT6us6HVu2cTMCXtZX03ZSg6P1weIsQ5dC0jA6T9P5v/Tul0X/uy
ab5SUvCyAa/UFzm2xxWl8jjIr43X6UluxSLSCrNoB0DK0h3HUeZ9g3HAtvfBNMfM
pL20VU78dRTUbJXdpLZSgd0qeZdWV4F9+1RorqRJvdQMr0/5X+ci67Wp57ftTIek
7p4yRJcEVFJNBcZ5W1TsbpLk0rrVrpBAwTXpYxwqHqHD7vJFLoRCLf2WPjcdf3BF
7ext5F5bOlr0ekKHQh6MwggykJ3rPsoS7uXjAk4BrE+sZJKR4ec3mK1wLiG1g+yH
xXUNgU7/9/lQ1RSxDFY+eItVXnSz1P/7fXfUuQBCWnxufZC2UgYJ51UBjnVc4Caz
vzYoX2L9ms5vFrxN2e54+dhcYhgTCNlOfMRaV2N0oWGVZs7EKJthwEvASeiLALhz
M4+SVNvzg3Hu6CQfuw9/46KtCJmEdQ19XJwPOhd6cg6hZmYziQYYTxeCFvcncsC6
/1Px9dNTLxkx32GpxbqcKQxU/lgjpyTZ/quUH2KXg9TlWqpLAG57IHnaMPEnpmiX
Z63t93Rp0J1AmCWHslKi0aNGlfPFEmuZUt/HfpAz2x3paFyQehabZ0pLN5Ul7HNf
wTMdiqYTltHE3LdFsX0AshifymW37lf6azojZZJ9qTcY6K4iQ/7E8ZeZSjc49Kb3
MCuY9WlfHkzF21PE1fp1D/ErePO4JlBoRD5MDBU5zwZwIW82J8g5zkzN9iad0UDu
sP/Nxb3GP1hvcDNJdcx3rTGbRogX52xqU11meMENPo0rI1vBue5xu2CYJ05rUv55
yLqYx2MOm8mqbHsSJzsB0jjafKZMaPkiFHY1bOc4y4yMplVukyuDXAnQywugyKBK
KHnuByM/w9+kpFTS7k9dL4kRGWNiGDEmLRKz+8Xqk6Eq2cax4U5DUySkClf1kfBu
pmo8/Mk4/OOcVPGvZ7zFxemj7sIAOqlsXHJcvgt8tPumJ530EpqwFD63MaMRtmLY
YcAlYbNGQ6++WtkGRilyAT9AOVVNrBRmQW6hD+PYpvyr4dNlXZJAynWeZIYclQAF
8paIZp5BQPzPg4nNn43LLdnYKvhCleA4o5Of9So8Hwih0L34n7/FzQBgNNhRS5S5
jmqeai2Bmr4+5rnR4tgL0T/l5F9yDy4zWJHezOVGJp97wkY1WOSs9P3HgwaeWRRR
AmQ3WtBfzg7Ih4ZYqMM9/BTBJUzldjMHOo5nnFZe+OQOnmB6so1CG7uMImNiN4GZ
pQAUgw5+ok4h+CI9gjQ4UQZllf+Ghce03ov5mHylbJDO8C/1qnYP8kciIQeJUOxP
Mu9SY0b8T8LoAXM1rMCikj+ONOQHGqVEF/co7UxcHgCvkgx/dvuA5K8DgR9Uhjh+
xmYxO04dS5wdFV4qgzf+ExP+wCQaRyTAij/sPghXDT76VZVVaL9W1PD79yq967DV
Z8gDoPE5qoCCoCugzfEOej3f7b71+W7PtSQ7mg3krA891PaQdiw16+xfisGFgGxw
mhglgkd8DEU4m3nsLZnq1Tlyacm/206+maih2UFDfdJvWpo3kMb/Je4tNSKSKbmm
pC5t+Cd61GddccWFElZy8QnhSag8H8txc8QWCWUek/bnMe7kk0ODjAyPkrO6yhxD
j6aaGABfmEAFbIseCdnsadBKgBfADzSssM0O1UGweHEHEWiZrO01RRUkK5C9yomG
QsO0MFZHLUAQp0/Sj+PdTz0D2XPxStf40ALk21S9608RJy8zPFWMGQ6TqgWEnNjT
zZv553YRiR9RXBlL2vGG8wpD+F4vfJq7LQWGaElttvNe297uMw9R/GhjTmLA7hyB
MejjzKj7UzzgvpLH4zoz9ekDHwQGBQyjQGn6M/rMV0LN8/JzCOuyP1HbdjwRa/Dn
wbubTVvlw4EWNc0920qCDZznDQ8cdLJiAUBqfnBXEkbLFW7xvOn4HRgj/yOQJVmi
F7qVqj1cm04BSDaprLCOm7ZWydULw0K7GYpAECIQVkLOTtbf/HoguvWkCvF5ml4g
zj0yeC5TG+vdiTDdZl9XjcqeAuEYIz/5d88T6zw1ojN9lClC7jLxTOx4ziEQotOR
sen1eJlPIVlbMf9cutbrmzVPCnN0+kmPt8Xc5qZzlyrk5Do8f7sLru/54YBG8+lV
e4mpDUn4Dv5C2hb7k4R2kfESGvD0tVrK8aNiLZRugZjJGWOmL8jgaMyrKOex8Hb8
pJIjly7uiLl54HkOr5VZh8UPI6Y4ppU0oC2gRQ84Y8hTSoX4VYkiu3XFlFtcX2wV
fkm2eZ+Ufxrxq5N0xydsHHEd9vLTl2Ok1NCDrdOI22P9JwkTe7wrIN+cQtNS8qpj
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F/S+uOJSAA2wCb5l+I4B+nC4LSK9ERXhzu+c5tznoOyaimKnXI48BZ/XKV/wvdSS
KoWI/3JKo1OhzbyNPXu/WznEffGRGMItdYTUesnAQ8hn0hNK4TD+vBLKZQ9cZLQ7
Byt+/dkDfbCRvnVtl08wL6HWWO9X/dwscCdOKIoOon0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22208)
vafvDSMKHt09ZmapRJs37XBe2MsqSLjS6VOKYVAlAUq7EesAU91MRoE7cZ1bZ7Oo
BtXMYiDpD3gHw/jvIr/cVdge4S6BmbvRVlyts/o9th97oHbWneeDsZXMRxFTjJSH
yOfO0X8cg2pzGdKqiaXXQhso3/OyEuBdXCJUd/Ljz0vfsx+1I2vBNfqQD5sL1Sds
PuwYo8pJpyaBizSJKDpMIgVyctZU9/wianGrMeIKuMywvgrvoKA+ZPk152QhUO+6
bLNytsXvbjkhz3L6VOoT5DXZOW/lbMe4EHDCLjjAZTCtXUguwB5XjRUFLZAfY9V8
pMyk2vcZdwKXPWiNlHldvbGP5WNBQVSaBW49Kv7XznbH+fHG7X6R3cA/y1vTAWb2
tHqeg+S36hzPWdPnsx37gd9d9xArtid6Z+Od275dQvdhIuRGtwo8hEEDUvcwNwN+
KU07TcWkFohS+jqcqSOuobkeLIRxJzdO0jLL6T+U/ifuHV5zo/zJ6yGYh0zOwr1g
e5sZJIqY3hIMzjXa7LMD7b0oRrPiAltbpzU2jM80aUXGCGZY+k7mgR9kC+gdmKdX
Wu9qqagP8kCJ8aFCMMCBo+7es5/hiM3b4fy2eGS8aGkJ2qXd9phEX7JTU2z0W9tl
3uIiuTXY7bMmJ4GCL+HBn92IjohoP0w2cOguoUwbGUM4vbF2V1nr4L6GYnzxCaMy
vOGofYyElvXUD66VnZX0kvD5Ca2qUUVpeMlyonTf0psqNxBnxPmG7UzKMcxMECse
4a4BXCooCMPamL2bIz9rMciafwbKAFpPW603Ci3Kmn9ZoatAVO7iRPZy8o1wJGA1
3gH4jfUCf429zX7zXBlYHCDCFmW/Z0+ygAwQx9hTkRYvDQjXiRUr+PgpGCscdrsI
e7PKyRyYeEod11ZBHjcp391UE41YBRemxqk5zQEyP1/1y2tPcdRszWT9pznmS4gm
wOYgdRgFP1Deh8uz12VucOlyZTh+5rfd10wEoQjHrSy6dl0v2cI46lKsPotQQNR0
jOwFRiuSe7hW6TURbhzzsymEhNt+3NpbHFnwI8+jQXW4X3sSLK9byHXn2x9QLqSb
MCWEyeRLhdqlrmWmf28gpLb9Wn1PEbFF2pnltRspPgFXSJoYOqrOx0eHl3w6IaM2
ogOiXqpdQskTal3wVeJo1ZOoUWYLpUuBuP2oCaBgDVhMZ3k45jHFMEaWwWtiAw8O
fdcLiDvujCC3q+naPTmsjSwtOqbR12qMmOojpFGcL+EG4mqcicHzXAA7EGs5xNPS
8rU6Yx5nMCnMlhLwsu5Xw1LRcgD0lEMKs58FKMvhz9Pe5vO0B5mfR3b7E+GK4Lyr
6QdQI7pml5cStxUH9BXARDgliDtDdRZlX7UlmNdHI9fA9NznBwUR5pUIWilgfi+y
U9L/nX2k28+NVUsrKKesHoLDC5quwkKeoz4/wHmJGO7Lq5hloS2TKe0sHvuhjx5Z
QL8YawbqRlApKOM8G5c0bbFFY8gbdIjfdEGJoyRL1GHCyeNK7I5wZFCZCQeQDzFB
0PT3tEcPHUfRZI6g0gHWDbREJOWLnuRcrQWM4XCXZFBPWKqR5bjvWOmGv9WQMzCv
ehpQR05aLQqboJqz0tAnC+Z9wC9djWXC57ttKbTVe1kFB5gcwc2iFwKgzXICj8rc
tIztSNPyibznYqdv8kqTRfhKXVXlR61XiP2R6sAgz3Neby1uRUriSA6GezfIh4I7
AruLEWpk4Fg3f8z+HIuPnOfeJnJfSvhznEuo+KER1smN7f+STH3Eov4t/uHl3W6m
RQnT8p4by7n4W27evUL2QsEs9sdw+uho2LOoA8Jy5MQyikZmLpRZveCttf0U0gz6
9F9jU/wVZct2oDMlu28i6nYSlizwup2LYWF3DnzKDxScKX1vWeW5gs0jd059IGx/
XmXKskk0wQCWTnJ9JHoV4h1M4wEFz+bZ6wl+BSoN5o/T0FMrkU2XV9LC6uEa34By
R0pTR07ZGQdujXQIubv3TJidXdx5Y1zpO2B+3D7vm7dl+M/cFTguMeOC/0OfnUMJ
WH5jfjXb0jUE62yafAJbuemXCuZLNT7n9+csZY2nEtIsX0LRIneEDLVUO0eIaaUH
/c4TffWfzqbtuZSlfa9/m0JKNw9PwBK5KLXUtWDLjslQuGkxVs58X+gSnJGB7VEW
CA25BPdhZfyxA4BX5L5z9i/5L1HCOYbmThon5EjT4FtUDLB9+RikNYmcRg1sqI79
gRqkvV428HbbHInLLpAeWP4L8VwpPRMi2YfgKWwBykzn2hrxCqZ8i9xLgE/4Crv7
obZPseXbDOqxKsUEp9va0mAGNnfQBPlYpRyYuRo30UgrpniuXaGnorD0r1ghY9N8
hN9iPFgRoQ7/TfcLyFcMl3qqOQ8d2IwNltMnykgfGGmTKMdw6eskjC+RaNDz8o85
yptVlRqHaLWKf6AFGZzaT2/+DTm5E523lrYdQ4kWSFZlH4eD6wAuISL7feD/oBhx
JSN1hgRWFD4mr5NExTFVFqa/WZCnaI/cDpAEv+6fYcGTB5hZIjaU1JqfZMQoPmMO
9JP71rDq2yFynqtBFp0DzvMyEjKI+onhTwUF6iklnxldNgHPRhbsL0AizNHn3HdS
Phm1H14jMr4ycP8gTK714v1Dypj9qDDc5iPii8x4U0CDEottg53wcv3xdg/ZnD33
5v0Ewoy+DVytN5WO8t/0tdzBZ0rDH//iEEthlJhmRK0H/NpsvsYDUFD19M29qYCS
nLpsb1AR4PUgA0+XEMHGY0/MNvyJl6xv8ChKk5I0x0OB6Fjsu5roBFQ6qImfXjDA
Rm6FbvHLLi7rnyWsw6JcoxgTMzZE6I53p5WaLergbPQcSk5P+gNvXpQMc+MfROLo
+YBqAN4iq45vODRpm9e/9RLfPkg1o+AHS4PVOvYEz/7T+b58BEvKiEhZ/fh5518m
n630Kmo408SIUeYej9MT6PtbGkq30mzyGyOoBdLHR+AU/iB/v1jicriSL6n2F4dj
ZcpCnJWAS+lEaPYQo0l6hL3KmGUJil/PykaNf+K6Ep9iEijAEj2GoH8b+K1Qn6iI
FRm6fb4hnLpdNgZ0eoe2Hb6MDk2I3unm0uKJtit8NJfjm4gEYmtsgJ3nnsF1bQBk
jga76o/WIJTG+BaJctvyB5PxiFqCCJvBSiVj86Um1J6AHO3YCIT+FnNaCboqfy8f
p2drFV/fKJOUu1f5eWODghmLQEQKBjoC4s82UcaN+jBNkddrukKgIl3GplNg0/F9
syHnMPIkJuo7oj+7Z2ExrTWmZWfpZDP8xXqWWEfatncheLHJO2gsWcb0qLUZbuhx
+vAIv/y1MKG+DXSVuq6pk/lpokFPMGMTJhwbDWylUdYHDQnbN1+0FRtH5rktxnyT
vrK67BHx0tsioIs5aItl6VCj4AHTzzgHQya2vXEfyeXJuEwAg7oQLKQV2M0yZTKt
NpLMpChRFm5rTgV+kQOJY4H0zRG/uaHivmnPUSY0r+mxSzfTiIvbV94R9c+R/DAg
invAhAE2FQbhT/N1DNltN6IXYYJsLYXTyZhlYqu5xFzCsDF26kvkhcXn0xiBT/Xp
C2JlOUyT7MfJWZu0tAO6w9eH02mqdWODYe6cnhccyO+0kffSQdU30z1wx0DtSOCu
hD/6zOSvVFrg+GXHQ+M5rE76OqxC6Osycd4MbEpTBGBEyJGXmnjjYU9xZxcl4Hq6
6V9LdCQjwVZlJsHxaNlTVypEYHtnduBsaD2cfY3IbB93oPFOtfPZQnIKK1GaZvDS
qxAE0cKLqOMNu+QrxlB+yPe20SKpQYMXR/zcHMc0w6mJOLYSNl5w+Ww7pM6Z6GCa
dk6OstCJs2WvYk+y0o7KVO1y4Qm6AHeyCs1S7Li2ueFKKQFIf/79MX8B0l7HZ9Ag
DeS2pYvM7ocC8IPWlH+bd7NsteSJvgprl/WTbI6GXlG50WqkYWcnr701AHeDExXF
kT2Fweq9pKMWQeQRC/BuPNixVhOpyGfJQF6rlGq/br/YaZ1Om5413++4xpXXj2cy
YD+nIQkZfUW9UYMfQkYZOYWvdJDpXiaLeBZ16v00Iorhu7SDCdTdiCkzNS0mxwqW
ae4cxeZcKYgb3nskOffrA2DYRbQf3pqrS/xrzA9Sc8686GqsuByMf6aGV+UvonG7
5zGqph023zOw+cGySTlqUrMVkJn0NisRcRzQ9ll0itq1vK24Ay7ln4pCYY1nf0mb
zh3zbbzXf+ov4nF2hRwGLlCQozSxhMAUnX0h3hIWdV7X5IqaTAE9RN9yP3i5glf2
U6jZSHxsoO+5aVKF9zZ1APUMQl7X6CAvT0FStm+F4R7lRorNs/2UmHKHOUJl9lvi
RULGZqiKTc4ZFB41npR+88ONLy/pBlX0MFHinHV277QaIMgIHyIW1kMOBFF17kqi
uQSsWa5SwNsj7x61nQ/HoonkRfayk1NSQodlsNGQqOKHYgTugCXFQFBpl3PKJFib
W42R5O0drYwdU54KUiwzhxF7qEfTkmAjoAPV3giruLAZDXFVVoTvNZmsOiaLDjiW
NwVLmDqKMpPngX8FAAnRDlrfFSZQwGblKs+B3kKaF0SJSBKhlHG7AUG1rYXAyKNF
t6DvX5TYZcr+hny0PvnnY4MKm1WJSJ8exVfS28Rmc+dFnjueS8CWohWEPeC449j1
opNqWuLipnGLm+L2lOoNLhRoqXFl3dNimTxO64CoyV7ihIIgna6ObEDsA3R2ElQA
3Fu4xTWQOdRuUAJ3s2Mk1ikMVZzFG1Muhr/0RXhUAcmtElLFe8mZHgJCxRxaYfz1
EOamtYFacE+P/RM1wLC8Sosn5wxEJgdUCc2GmrAlPNEWKsPHWaRIlDxc4yvpWbUR
5DiIrbodZemLD3nZVKt460gnRk3xW9MwQG+u2nTK51/2YzgOsk8z8YDNaPt/CUZl
MHSf33e+TXLgxW+3NVygogq5cwCcsnMtxn7VYFybYR4rOCi6+Ik3rrARD4ua8mer
cYoOlrH1xnJdvEpS00cykNkHfBTwXOFFu/8n1buWlcqwEUGoTke40+G+XHSQLjvI
qHI31QVLAHVys9ZVxX2AY60+Zr6+S5xHzvWI8mwuvVK18R/5oMhAJx8RurCWD9AE
LW+VtR2DfP4vSF3nXkAOikMlUvByZg6oLE+hbEQDEWYSLdm+sDShGOzumZKbTecI
Zdqpz71RK/5WyHKfPB1Oj7ifKZHqAFaq6EolEFTei80ye9HAl3dsI5G3I8gqxRsw
AIKwCGN/SKFE2WNkKpCe/pVMq3aX2gtG3DsY58GcdnxxFCHzTDWJKMwDWY/evyda
oLgq/1sGI0QXbbapTfT+dj/OG7Hc7OpBeNoXV7prEfx8GBIwxt7OR2HhQILBO8z2
QcUE9NL9P/ZPk/3hID1z/nO/RpU2at3JzqGt+b8wD9Ls/ZsxkJfUpnEsyypOOSXa
AUaCOeQRQwo2+LpZ/c4TWN7+bfLhM0bfnWpWFOR3h449h22gJcACOjg4rtpJmzFj
oVjJn4sA/7WKZkqwrHjrxYD1aQCmhLyQKv5EXtpwlTeXWKTzxvBDcUkNt6pygxh8
KhgBQkb5Ayitis5fOqQ1aDdFTigJAGlY/tRSrkJX1ZX1qmf0qg2YcmHGcYRM/taE
J73+QUuYy22OuLYmm5b0Lcgll5A0WJRHlGGjCskzxTlW3UBZMpL+knzepkCxv6kb
9we7AFDpe4AuaLmNgR56qdOouGMQ8L9C4EwzLsrI1Czgq7bMVIBKscR13DiQydi6
QVsiKDnHcChAJTj5aDM4rqZEBMqFQ0ZeJBOfwKzN7a1tch7ZGqMDCPwnF7YzdPhs
kw4sobSe1LLEPOYNDwrncpG9hhnDINUDWipCY518CS92UDlXyxvBX8NnvH78pReU
5LhNxPsZGatDSymGBa+VxRs4I25XX2OqyC23J2r26pNoxf3UJpNCmt3zdkfwZghx
9dWu9jobMJwjVlScbBj5zwMoyUpFTsBDLB7kxlxd3PVQ9stK/8TvHRaL/76HG6/F
jTAiSAZsU8ZcEnq45WFTCsyeixzpvXf6wZv1S9GJNivFk5P5TTq/P9w/MZnjJdL0
u2a6FGswJN+v12jqP6A7uEzaIVzf3gqND+KDFTl4u79VlwtvXhu25YfIr/1x4EK+
oRRdcT+qGnsQdJ3OiL/Tnucx8Dmb5jQ8p/vlrbaAQMvdsoOWn7yPSy5QNM1kIsgt
a+1A6OEopLVrV8YhbZij0blnvR/in/Ie4XB1DVMlU/LmJEbgTKnxIAUcDWYv2MFk
o+ypXAvg+j0rRSKzAbgpFXvuYO/eEVOdMBO1aw9Gf7HvAwHhI5lGnnX7WhxCQBLg
dR1ELEVwAvuO9pqqSoVvhgTNe0UINaYHC+rXPmfRJHqyJ2+L8APu2/+qoelOxWac
5prerSC1SQVp99ndoAKs7xa2JLHbftK+uOcpsrOYNPD3JmvXre/IMshidWoP+va6
COgRCIghFtj2S7As/fmCUhF/iwFgsDMybNUh45xgXq2yIYFQxGj6P4XAjoAgFrSA
Iwb4pEQBSMkuY1RAD6NsPbnm7dUq2O2Ayhnf1zhJgtj2/LQrtnkleg7t5TBmkXAb
Lu8jou7JCaZs7zoORpziC4V+d5sF3bTW4SYCE6ZqOBqh/qNPbxsE7q02T0riliUb
cDif3t9PxKPB9ybwsVYmbIjERdwL9AZ7L5WtwQs5M212HG0RSrxyDjULNBc9MHS5
pY1d6D3uWEBVcm8VbJ7rQ1eC+ECdAxxP8jltlby4Kbh5yBzih9O1kNUU667FqlW3
yUO64ddJrh3089v19VupbqMuHigRTmkUTzm7Sa+jxsSi0YjCPGDKVydMZTOVvHi2
TXtkTPAZMBfyXLYTI/31oTXfKomMM5wRWgDWd72FrEjxzhUqo5AubAT3pPkHSURS
iDVYHLgdePTiKHwmRjqn8Xd3JydsL4hFF0l8ajVkV1p1fRBUwfJTZmoULF7JF9DU
j/79myiOQoF5h+EFXjZnobdk1L+wuhONcxQJmWrjiR79ZTHcm8wol4u4mROuMwSc
OBKdLXNCQc3B6Y+OaD9bbt9TVK3RBeA77rgOJUyhiVkSt7lbz0v6MEbw3afVjioq
nb9h/u0Te6hb9nHFTTfhlOJEchOGUkrtikzfIQy5OdHs+VmfEi0JZsQuk3QSZTUV
IjNdeYWsFc3vaXBYxT1mfxELgPttI1P3Wda7XC0MdIwLfDu0cQK8Ah/4pQj0re3H
jbup9yqPRDNbHn1RBRra3fXTzgo2oztGnLElGMEBMPVqIqCTyeJW2kTlXBigJNHi
7B0/nvujn6ZkScpHSQnkbbmHnRGzUs1LVTAEnQzns0ihtmXLjcVo/a2R2znPKP58
bTGcHwf6gQyNW1mbMFPMQSC3tN4ZA++k+OgQByi8w8eYvvKVdWMZmDr+tw5VIaNm
kHF/gBt15pCyhOEGYHsScQeKsgGGr1lHgrleQM9fvA1gob+lK8acubSNRkccZbDW
EBUJm4owIILM6LBkYttUddjWAqxcj4Eq6t4YLOQreOpnnNhsN59/sb7+CGeuHatq
rs8eh5y3XuheMdZRPcZmw037GwvjE7dbRAdEe6+hafdrY2SHmKIxJAEz99EaMEkx
14vn2MnSbH7TwGeG4biMVkc3YZYWgTYuJCqJgChmcWZAKd8WT/GCa56yIq1lTpov
TMuguOliISfQpBbSMMvozGRZ8rzo+zwNi5bjzIhWXxBZoxBf4uH7kS2C/TQvNuCJ
kn/6HtliVeYUSXN6Mw65t6y6i80Yn7Oe6BuNi2K7K3qgsfpQlgh5PFd237/+XZJd
QD7XJvgJq97XbKVIl65ffaTQUC7nu+7wN6lwNQqqvwbRdzvYhH8xerf+8ul36bEl
Hc/JXZPlPpqcLX0qabxer7sIOT8dwsV3XQNmI++e8uLQ7s0IPJYW+Xvm/zqj5iTj
hDAIP38+xn4G2boNPhyTk6HUUC3+RvU59Ux5MMa1s5IzfKS1XHI055gRAn2xze8M
0gTSF9V9FXrWLCuvP81gI0JLe+R2DIMbJcsBVo47+cilgl1gwq6hV529o2oJf31B
4xBzjCudFkkflty2RAQpklp7ne3F92HWw0Yi/CjLLdTZmitQAv+7o6qgR5vpO5Ww
/34RmS5DsK5u7miNopFYdWkmmNyokPMROVCqLEbNG/EM7Ua5dizIv8VduylCnsIx
ONfjvoRuSLBKhrpaiilm17E1B2CcVH9EjgsSJfxGAiSy6LpsEJbIgexL1xEF0hir
KjcEPQDNcl6Jc4vxIHlPuWXukBajpwsia+S2a+JCttBtAs45H1VORrQu3iw2K4xK
iJsYtpiBOIcnKRvU++NTe7mkxR+VpNlvTuBDnqOvPQPSbOgf0rX6wR4lLgPAUQuZ
ahkmNN5dwuZl9t55IiNUqTdUwwhGmzRIoVS5gdjHUfEX/Pwq+6IDMlI3gXoj9x9K
1dqQMdiXtktNOYjsCHOB+0X0O9wHONHnguExdcA7EHvgRURDr/pd3ZLSUhBtZIPm
iSc1MO+MOoQQ/C/xdd2lhVOYy7Z3PEIdSi8C89d/zEBS3PuBH4CrA6/P/rCYxS9f
6i9DcaeKDZgjNL3Epqrd+jzi5JA4Bg0j9cNvg76jf+bvmyfL5JtMXqErMthLf/eK
rqpMW1nqVWlnB8pvbn4ThZ9F7Qa0uMzCRPX6AknOj+RvxnDoyZdoSuKuwD1/3SZO
71Vk5IQ/xOpjOafGF2N+/uArR2fiW+KCAWGeYzkkGMeglNerE18D+lDrP+65jPeE
ZTizVTLXjqjZgw5SifyUhTNt8OOjeHYUVz2jjKTpsQ+nztY7Eh1RVm1C2Q+xenT2
SfwcgqS+7ztWGzQnIs1A6VllivAoCf9ECKKu5T1oHIXECa07pkE9ZIskXXEXZ5NC
tAbj1yHIMn65J7k3kZYOD1TAMFVfOmw7eyXpBDTOcTWZ5VKJcacnWQqaD5Xf9kvN
VpLk9OxtAf4xhQZ5JYmHOHAS/ZqKgmWT4LM9ELYVK0Cr8ZHzAKXZ8QB7w/7VQVmT
yaCqsjC5xevUcbwzqhWF+U5s1dulki0w1X5QslFgIUG5oU7vIllMC+vHMyaGMtbI
uUtypN6+aZ06mH0IsEMn8M59WL3v+WB5hvojjnH/dWElccVV2D5RdsRT6bfwgkgd
RJ46dBsPN/JFBbSKLQu9tV8M9wqDzTTD9TW4k+2yxh4FZKi0Dm9KIrFgskIQNDyf
rV9OSDYH0OSx8knxAK0d9XkE/7t9cumxgbuf1w9+Vvksp0eQSVshUsbtoNc314S0
yROG1hX5t9NMxZJtiEz/1Cgzh9mdfYPNp4/0/BUrm++Qlnx8Vz2x7aHm9YRk4/Jy
ibJOp+++LyOjW0jCVxeXQENSDJEK4KSPyoWJfx9XjUO8X/lxMm6Oeb6/Qg95Ntlo
DZN+XvqhQE+l7JxYPzDuqETv65mzA4a1G8/xyJbdStpqSsHygaHRue40O0iHwj/r
AJAp+aCkKLedW9k8VT5MNiMAA7XrGCL4OdmY57xLA+VSZ5MnHzYXldv897u6ct9b
v8e7X3VYII77tQ1ILH6KUTH3CQk0avx1NdnXOOHt21RRCNUo7tiBIS56gq1pSdA7
0EWDWkMH1+U3aO+VPcrm8nDgEwMXPerAcuSWs6YDzL1mKQh1gfX9/uPf4iHHVrNw
anpUPIxc9c2Gr/Pj8ERPDekwS44BkJz+Z1ts7XTMdEtYNFZP2OPR+ffkPus5cWvm
BBd0jtrZaxjqKPOm9S1kX8kDLsh5PjPT5wr8SRUcbUaGeQdWqfYSdqgRlXCYioLx
Dwh184JDtQ/Qi6vsOJZd8q0MdQ66X5N0tb/E7PtFEO75ssbO4YGX8lHIp69lVfGR
IqF972rb7qkHQoeXeyPj9PBN5/bBvGizlSr/eBEyADc4QJlVAWMxt2BYsqh/xFzO
Tz7jNKw93JaJaJuLfb+e5UNDOrxU7euIzpBsUZ8U+Sg8n3AaOHfzjtRiM+XGd2GO
kQOJoH/GPnuDm8AdWyY8dNMX3xpt1iD/QYZ3Lb2gFZqulwGcKN4L+lc2lDMKLqOw
nEkrev0deVdVR5DfmwjO7kZIOP+IfQhl1c1Q5EMnpw5WkGkXl+p9zKU3VJ/JXUV3
mBO8YOXQf4qTJ5/tiK+lM3T0ndAPLHsgH9P7qn0wDAPpQprG94wrUpIWShzAP6iT
AZL/EwVLP1qvsZcZYSO1pZa8pqj9UsLJyN7Yw2Y/rMn7DSImJP83QZ978TaMzgBP
RtHuhuNEUjpd01pCa91ZqmZENtc/D5uO7jhjHVzs0m9jWwtTuXgFMppyC1oL6FHN
6+i/NY0WIynV7iowqABZ726kAkemjx8CzU9gSRHkFtMO64UvAWe8L2ltd7c+Ymis
fjd7fJwNNTY7ULWCQpYmZka7cGhVExe9ISpp5fpx/ctT6WDDZZWtStVb0JvCJzau
GefsycN9hEOyzqzM3UjH3j+mqUfLte7c1rWnM3Tesouf+qbIqKN/JBOs3lbS7ZAg
onn7E4DvdbbaiaAZJu6vTT3sONjqWQbjvoYKol62yCGIKdIENjLeJ9/NdjnRbxsL
P0aZsqoHZ6+anvCcSTFxUP8XdOzBvQ0ICxycAleAVfmnPhsztSIWDZ8FVreuqwBt
TA4ZzuONcUGqfjkLwh8Um55LHTBSPGnZRCfGeUtmDgbjgSPd9egGJD9C0Zj3hW04
r3e5Sq5B0rh1TwYoOPm789uj5N+mgRUXZc3mJejEWLqTCmO4ondoDrk4b0xbRdnJ
Sj39ygaR6fu835jIxvxHkz80Pp5czeYdG0C3rlRjXb/FFt7VteT1IQ87rOm6GIvm
eWdmZgnjQlncOR2dc+0HrD/WhqsfxR4xdvN0Xw5Qb0BEDBPId8pCws/VzxiQZCoZ
/zASZBwyunhYFwpO499Jjxt5UmrfK/gKeOF8DDQZp8YvhibXd2WwSJnre2LvJnq+
Ame8oQunpGSknWdwJJ90XQg/mpRGXz4lvc2eScHzai/MThj9U1QVMwmZiik8UO9g
bCD0MdCfRxesElBXtUO89RE7KpE0rIhs+jZmGu0YftnoKuHQzalN+p4RCY/V+7NY
HOc9v0WQKlWtIEXhPaUJPY5bn48sk4s7ENVWKD4kF00QwYOaTxKEzR2iqxn9qMRv
/u1mx6Yk6xwY3p+4ahkM2zhD/gfsCt7RlfAv00K6DN+/+2XIrGswqQJZYDEVfQIF
yqXuhCOlZFgmxnwEC5eoiaOvcLp8JgvSZK8MMfDmMxUDpxILh+8O7dRdc+3T0plQ
QYDN6J4SeK60m/ldte2p+zojjpcahRazpQAOZOGLqaP9x1LaxI5RjWmiWhrgC8e+
xBoq4nsIRt9vsxtL6cPbMT7dbAb0AaQfCd+Hvmvnqr5JmN3clg9vAVAzvrjzkF7u
knGoyupiQA7pBdss2R6Aila7WOhn6SQEQ+B7YrRVrT4V3oYcA7dvq1epvMREarn5
OtP2n914hXvkyRvHoxzLmq9ezbAOJSxh3O7td3X4Vk/mqZX3WhCa8HJmX5ec7nR4
Fy2oeAHo8KUJ8sIi7jkDPjQFeA/PMO/wdnJs71NjIZ0QKsACoJTZ/4sluNjJrlMi
a1ofvnOSH68axtrowpYqonwMQOXtavHCwLWB2OvonzsKSM4TFCOhqGhAM74Z/Cki
91t4a6PnwOT75c2vvjNAR4hNw95lLXpNJsicBV4a4CfgaLShhzUXEMW6UYQQy9fL
QA6AnE63PoTofP5nq50kFifkOIA26e07vdcmmZj1tP4+PEhRmKwyCemd4BS/NS59
zypvV25LoP21BSLxgqC0mIQjIdt2pxktyjtyE/e6gbq4PIHA7xctAsUKRqC4X0/a
veKwTvmZpu/BbJZrwKpgxYabBawQglmvh1t2ycbv7vO9l5ynzLbqowx0HxLLg4+A
Xl8T4GUSxBRShm47glewC1gx4bzQaJPaCUC57JHbcyjs97hs156b+UJNFhNccMfM
+9uaOwC6LWkmd4ogTHY/d/FTPb5Xu7EXoSkWsWWuM/ythK5lq7ajBqzkYQj4Ev2N
6Mn4ce8AADp7VhuE+Z3ybtiZqfACGnKgSPb5V9g2v0aGWwvPH6u3JskeTbF+vkLP
LwjhlpAimi7G3qzBrBpoor8fX4AhNAVXj3YsOHxstN0i4mbqavrBpr/PBj8yqHA3
g2cgIYDNtGWDgtKGyMkJvBMt9JrXhQX0mKBTj1CniLIjz0oiBrzTpSPYu8zAVzPt
kkdNMWjYPGm230AqJ5xZyxkvyjxOktgD+pdsI4s4mwcv/15K/6B1buMrhUwLea7v
7okYIKVFCnYOn9pea+uAh3XJDAQMdAo2TOjoFq/H1ooDImjGroRsmIwaxX/NBj8U
Gl+iH1awGxF0yyEwEhA/qArujBGTmc22Ry7XFSUFZ79X3GKidI/lPpAboubdxT7f
MTHp7hY+EIUQqoXJYpsPkjeid/9l68Mi8lqOLmQwULclew/CTmqCdbTJ0nwCcXRB
QrWp3wS2mTNnRWNsRKz6ccX92b88TMxDOph3Z7k2pO9A9xSEM6kpvBZtkUJjSfyU
IIOC6BaWugaQCEFxXRDQO5Ltl3Yf0oFlHpIm8gjz9JHpPDGw0/PSKS5TcXPKZVL9
T3WHSWGXzAWXF7OVFCLapTJMbaSx3N+aBeM3rH1BS98UFef8+3BewB31zhjaAKMs
CGiZsxVE9dc/nGhQgM9t7HroJE9Av6pekYbWgPD0xdV/ZcfYBcCoKFMREsCLO32D
/uZCQ9vppPT6/0HP6DT1/l6HrBOAGHsO00kp81LT5WRtI5Mk5BA04IN1dw9bukyP
PkcHVdthBRj1o9aU0kwCv51bEcPHYAs4835ZV0DIIZvQJg+JwpNwfLtd+lhj04Js
lP7byfGij9P0w5jcRlgTbSjbGIkPC65d4xTvu44TPB3WXQHWJZa41WUNI9G1PILE
w8HJ3OrAZwiPQqvJhyPoWQLraYhXa9SoQ1r8feIo69KoeR+skNFGXfr0VsmIAjSr
Vy+y5pnWfBFNB8tnumw7IiKRgi1MB3Q2oaXeJfXeBm/Vx2gJxoIIM8W4ZcFoimor
YdrJ0KVBxwubhjhXIFfGW1bsXZ08JiaRiMWPjF3v3xKY8VivtlCVoEbljQiI+EgJ
/UNV/aPJ9lYNHFXVxnT7BNoW4Q6GQDbXLPEJxjDpdIhzIo3DngfDyy9fxg7aCGZH
ddQgNzyWduKj2AI60B1X5aiaHK3pV9Idm/A5Q6qK3HvsY+1ufShhwXfpNpnUBuDQ
iwO1jqbdKgi+DQIrvfnmZz9ExYiWC14DWC9EG5N5nO6tALA0mbnbAutoQM9KBtUM
0QB9gULlMtv/A+9x2D1xsMHUmTJthFUDrJJfGkMtPYtKJEHtalFEhSIklId4wGu6
W74wwjcyQiVjPDygJ65LT/C023Q4QfzMAcACN8Q0Z2uvk/zemJCbFrl9/EgQL/an
75wjark3pXrVsDnnzUIs+c2f+E7l8d70hUiaoAJ5YQO7mRzzmGdPR5j/9GDtntkx
27aZ9dcFUbFzKU9evBEZYjsWilO2wlflT1cdOASlYO5hXw22pUBtI9Nj/H7p9ZbY
nErvLvbElkRqaopz2+ehM7K3LZurH9ez2p7qP9fvRvlTsTIYbX/WaQTziUOG2VGl
tj4pDISRbYqU/Tr0TaY4CF1GKSFeWl6bZD2sEF2jZE4UtVDM2H7isEBsDrVbjHOS
C+bcHIe736U6hewos2TUf4wlwF7mZYyG3d53glsbBeUFFPEfMwiHMMb5KyWbunu8
NdvSdqfCQYxjK1nVwaDL+/+tW1ACmV3PfB0PaPNSC/IfBudk9sjwm5n54dEOGFMk
+VG5OVQ+kab3nyfQQpopBeYh1YuJbYcXl9IG9vb/Y1NCEZR5LL+xdDnE3gme2lT4
U05+g7fz0Ro81t/nAJiqjvQb+uW0b3QvjArjKA1dZVRYEXtEiStWb/moUkWGtRmV
cy3F2ulkLR1E8Os+2PIiLtjyOfri9VJQrxn7p+UQ1xNtvPZ22yA1XTMGVTLIyDDe
f4aGBDs/X9xk6ekg30yX1yMdVO6IjKyezrR5sj0lX2QVD77pQv9TOqiC2CNsc1i/
UxKc/S63ve9gkNmnS1zPyQfMLCkOy08jHaQRSGAlkfnjR+m5oNEnmVECxvNdOoHt
1fN70DpFBC/2Kc4xLU3Fw+l0DqZaEL3ZFNK2M3fqHA1JRf4mNBDk+z3yWfNLlD7l
njyXmGlMtRQrhgIPoWUqtu7r8NEaipHd9GXJqHSZT9FYPKPpyn81IkR4RYTlcmtz
d1GX8q4zPoxV4aXMhMdijS2zvOw1UjRdQmdy9htLCvji+zpT1DTABj7xcLILbThR
GnIOeTM/nr+LPqrf9xDus/OB+RO29I9COI7VV3M3DQisJMUsyap7qwy/bHHRL6vo
CX3g5CdHin8b+rR2av3rpQWvmiVvwVTMKNB/btzv203EnaKfzMXKCEuLZAAI7bEB
hSPoSF9dm8TySLWgvvp661ntzd/lIbuqVT7Xaf+4KQWEBaap3h3ti5ay2gB459bU
kFEogAd/iYdoophrNvM1KICpe6ZV2YxObns8EYzIki2TPip4PAva57M8ODfFdNU4
reUNfwvAK/5EeBabk057Mxmt5nA+V9qPi1FaM16HXksQ/Vt+a0It7sbmIJNDHYjo
OrLtFmRosQKa049Nn4W2bs4ImzHLSR+vO1d05rsvhJ/jAxKHK3KHKgJ7CreMhfhd
2Qsf6g5CTqex3wjXBY60MaHtxjbNN0Z/FDZcYV6ht9n4sYlpgPw3SGty4S/N7Lo5
yApBVYmVZDWxTO90+ERcPRb/jfiMhkM+cU6Tv4IWmaMXApklobI++9zuAP8AfVtm
T6U3bUk42NRdfmtHYzHXhgfMHgwcquY4ElMoBHRaiCtJvwfq/ovIe/xp5GKu5QuP
qhm9PF1bZcXd7dDAjBu4fyX+kHQb47f3n1MLOvSDT/u5LcaQTfKIZhkqiPE8iyvH
p5E7/V+CN19QB6+qaMlpqO28clMJrsYnWinlOGDBN8dXAGWxsAn03qys+0b6uIVF
oyqwLLoGhj21J8qguLfd/RyrSECpW9WKacyOMRdqV+LOL9MOWfCshwYgAYQQOeO6
A3qHs+O0ZQ+baijmvb+Csf32Mt8pE8beJvK8/fzftiyQOPDyDpAx0GdElmns19tg
3RY95pl+N9cWD8mvOYEtKLbVDghpm2B6ezFO+3dN3KY//VY98VKzMv17RdQL6Ggq
/1Ijf+5Dyy0GNY7nbHO5iZI19j6RWOhOE2MUAhGe8ksJx481NHPChEj6oApDLyyl
30rvNxYqwgM0KbXqOxBIMMHKnS3edfKosBEGiLGgGBvTmvwbOdEdzh5X4L94WyUG
V2AymrZ4ktbSrbLEKcihZSdmgn3/TcYJwUsQ2mzCFAJam2d6hDEzTELq7bctBvYI
diM7ArkNwoQGirOWIn9cchqU97QJvVxgvz2rBsVg5WFwOXm08IJUxCGEbK4n9T9P
ZLfMelDge03c4wIQug7R5u6w1sRWUKz+kjLlpU6f4GR72psyqqNe+XjEeShpM0q6
0T4cd1JIxP9AK7aPN4hLzld1Z+4txhffc4wkMqMQOAHjXov9In8O2jsNQptEB6Ky
fxjaPmK9/svdhI6xrfhHorVta8dxzWzykIJSbobOlMU25wi1qRykrQCO0gSE8flm
UDGIMKuWja5f8TJLwuw8lHZ5IF7MIcmniLOUI30cWqSOUOs3WY0jwv13ZVcGWi9R
xxlL2fiu69adJ3NsBW4csg8gnxFSuC8gn/tAEIClcEXjQbr5bLPuBv/ah9UCIAv7
tCPT/vRl8n+oRWer/+ovdq/rGiL1glT9N9faY4+EnEmLp2B/yvVJPEBdKpcU14pN
MnKtPZlg66eY5pugL/SqxNa2RPRYKvc02VgvP/uoM+f+N6YSOxPmLgS+C8KL9C9Q
mKbjpu4PICkhISb072MxxYONpPnZA+misogPPc+pdEMs48MP1AViJwHsuWxUogrN
laAe0NM2cSKrOrvHxKq7bIxbRMvtn1EzED8qcc8oHgHLgRpXMyyi+Zfeoj4xonsA
IMTorzkpT5OJPEHzNXL+iFz1eabQelwRO5xwLKsFO8NXcxM5PbqItLzS//NMGZXX
G0ki9+RRa78E/4aDQ+lEjcVT4SY+2bnKb35BMGs3Hmr+7bV+sEIGgeRNSzREQnEN
wl7d+IpH9G2B/neeUUotdIFi/4qwaqWYGiCGrWbTWeCxcEF0TFApGPgMeRwJZb9e
7nYZ8iXftfSO25DUr8G6Gm7ZzdtDRQAKFExElvLqtEO0pTN+oZ9YwvigEsULLP+g
IKpMhs/vSB5zE1iRfoslt/Yr1PC558zKq+xXy4BegcQ4sabsH6PYO5mWH5VxymZt
Tehj1e55ZkCHa0OtlRLRg3TTKpvZCS6y6Bt6Z+/MQTfG540OHSeoyDE7EkygOH65
cbn2jVw7oUpwlTRozmM49/h/+09hqw6bprG7p31IGioShNcnVIbhirkEWa7Nx3d9
a8fA8j2J8PnQOnYiDy3/tog3lmCC1UwtxWJB3kTROvLM59yeMdmdQg6Gpcwjawls
P5var/1K930+Tf56AyM12xFK8USn/BMC5EnXPll/S1GPtpgacXYhJw1Hi7lhDtgP
PKdWAbjVQ7rY99D2ziJ9+O2alirfofP1yeXjTN1pNY1q4bjcUVJPdPrwjFuAHyuB
4/D0ZVbbvTTNSxF8VlO6ih3oEnpj9Wg0ROOonYjWRwZM68JhSpptpx2CrTYBI/TH
kh8yOBXCJqjC6d2DF5PtuospQBh0BOxRxT6CiHTwJSsVoTxFqoKevk1dgheLfwew
xFeSep3LjKL1BJXPt7M2Fp49QBNAh/FpNXWJvO3OkJ+85u3vQ/WW4yRLxEjG2r21
bEbh2qQdaXUpFkiUSimdvttDoejiIV4cFv3lezQW+Vk3+aZ5jyrv6iGKwFJJRZe/
Qd2KVck+JKlFv+KPRqcK515bcMM0mj5CO3PCHiplCnMbyOfYzJjcbYzYbDTVABtY
NRMaBoHpF0anWdPpeMnmrKj0aedLNaU/PR9NA/0guoVom/Jo1vWTI70T7XX7es3h
1OPnTjsTwvjTX2/Tp8dwJPAkrRwvREmzkmQ0b3zeOAQmjq5gw+ddY9/QFL4oaX0v
X4EnjLwuSbDg1cRFXjrGRI5orzATdQED190lbCnYg9bWW8lWLYr1c6fHyjsitcK6
bho+vv35Bp3e20obIeQtg8ZYx/YOHHT0Ugodu2wrXffh0NuZjw4VkAu+JGoE0h/B
eZtfarFu31geGplGtcHfL0ZQuYCTI55YJLj4GgGgieZx//a8BgEYzQ89EN7UxRan
y81rKCSnPeM2hJOMbn1zOzMLwt9CkvEi1Dd83NitVkroZd+98tSr3dp3zT1z8xJ2
53hA4s8rTTnJct+6W4UWRwfVVbYddkArmJr8SIFYMAh2Y/iK0XXxpttfQp0JRSst
EugUIwprXUkna6wmZcWLJz1hu8Gf02Zm/G82+JaHJY+PZEpk3ytg3iDSeFGPobkR
5mZSFVd3JYP+BWYaZBKb+wBKNpH0CPQPGbHI0Gqq01ccX4gonSeGhAvrgYgBMVNX
Ot7TnGg9BnUI1Vn5189yYrTGkHefI5cNbxuZc9JwMeiAEH/uLzyo2Up4LKlCx8nr
c0GUiHjeEraMiOurFUARdos78P0Nqqc4qFs/U0kILy8v7RhENl3ukayAqhZbXzbf
cmjxdLGHpkPxM0AvD2bU1EQUGN459T2BzSSejjE886/o7CCIHzDpXLrFV9BllDBF
C4BFjO3TT+dwJrzYfVnvgZ5vYmq5jBlY/VLNx8huzOFKztf1c7R8wQXJEX42j0Om
CSNA8m9/2jwEqgI2Om+lhm13l7PKW8mZE18m5I1vYSw8SYnkIFHlDDPXa8+yC7j5
BHWWFE9oB9NLP0HqnK1dSjdYSB41NFrFHcecNUPYrd2YH3l6LvfqSf4pWnwbx+ou
eg1EqSK7fZb23I+B36oPupiLh7xMEeZ2G9vFLt3Efm6af/j8n5KZlJ7faYSsSy3h
a1rNPY4vL4ljgEiElt+zyE7BJ8ys+QvTXdBIjypp/jYp/Q92AyUuhm6MCdHJLF3u
sU2hWNvdXdYMUoiiVt+Q92f2K9l8jJSQr5VcA0Xc69gbiav9YDjy4CrYHNrYLsCP
sgApfYIf/coPlMX1lhjwkUI3Hxqzz7dS6lOOI6SeVN5cg8+rKtaIyWo3kOFTgVeo
BI79QxmKIy835CNNdeLp8YSyUHq/S7KvgYhh+gXfrBHch72GV6pSbHa8vFC4vQQt
FbOfeynEbaTemN0HZKvPhadcUZRoE+BYOWeLAaR1njRAq8XKxYoKSSIFFrUsM7MD
IPp0DhA8DiN3opjtX0xVB8yw5GEmlT4yWgSSzXV0LIWM+HRTjxjRlMPPfv9Cf+fU
TElbbQA6fpdU4jL2JebHBvZqrI79O+XSCcIJJzUhoL3aD8AmlPn629pgLTrCe5hS
vXJL8ycfAnDC2Bzkg/N0ryVvUx3lj1VLsc2Z2cr7+7fM5IScZcw+fKOIGRXSF8bj
vS4iDkimTtcLsDjPe4zsUAvfQ87HEAObP8sWBI7r0NOE43FTUknYMqkbNO0e6Vni
21+rAX41CxfxCJucQADIi6xSJ9LDu6QNaLqhunvJY7Fw+LDUjpARuvtXx0q9b836
hYAeR3qEQvrG6y+pOIMkXsCem87wt5EYIUhP/mmcKyRVTzWF0cSeSzfVhvOaLIoq
X5Dh+xkxF/WtS7d29z2EFO/+WGENgqMTjI48vR6gitr1TbGltgQVfNeAQ8QaV1dl
s18iRjQltgonj6uMzZcSeEzB/xk7cK5S+bG2HIFJduLTfKJHOxKsZLl9/F4/eCnT
To3CuPfjOSXnNa8Pr5U6FLw8LzNbVib3Tsc1yzxFoSU+BfxAr5genjn0o6vTPFHw
pJrzLvDzteBwBEUXXUlbF27QRezQJNMfYfGuDRE1eIoVN0DJelExDpn9YLsbf5dW
jaCw233FRMxn4jVl8JUdZ4ff5qdO2wUJzC825ST2KYDRl1EyNDro5NyCvavMQlH4
znOE+x0W40ZZd6siytj8bPi+KqSBJDjuZc0pCmHoqv7/h+33A6fBpPhU7M8Hf20w
DI5AGsOUjaJoH037wUB3W99xYglecMA82G1Tz0XXyRKx4PG0OVx/NUlObOslq46u
GlvjururEI1spLZUifS2/4ZPEw6bYFW8/4972mnhHVZn+xsflbwMG+9vqrBB7eyt
pCzTpH6LCExE00/Q3zfWIxjOhHdJpbB/SmHKi7ZNUjvbVkDWcIRantqgr2spXrwa
fHgO16nCfyyXWQJ9Zs2nXDOqAgO2/kNW9ZjjzEx6x5E34cDDlU8rMr9v335M87Ak
log62KXOP/5EqPKGwdujPSMhCCWIAqIc0Wle4NQdKulWzkmBie+v/PLTXC/nTd0W
XnHzZgWljSCO5wiRuUuEBsK6SPDL1qUw4T7kjWZIMUsD0mrug6zmCj8WiEfVKX4Y
kG7xSMC5RD/TNgh1i0qg/BT8zAM82YD/3CQlVNrSeffBtsLCjrYD6HXoroN8SSnj
CixjvfZAXE992Bq4Xx2Wnbom3xIaw8X6/6ZBLS+TpFMMbHvgbw+QkFqKIUeKFXO+
r7SE4oCCa2ADpliu5GYD8251/i/if7GnAZ6VTeGjdgjK4QSZ2AF3HLRIwNk3UPNt
fAOO98Il1caH0qiR+Jw+HOM0IDd3OC4rmZRe6YvHNOPEuZUE1QZVuZycFHVgsUCV
/4eZ/Huy0RSTky1lbzUPv1yhYIrLRdJFxMYNfk+q+i5ySDOTUwBh8pFKXdc8jhPj
2M7EOiqp5tePFbDlN24RoN16NSV/Aq7WhZGYl2oqte3oV+mPWaMp0830/JvyYjkW
hIjHxMkYiSjCnFcakvCsT5gzXNGUon85B+oOO7v01+wE+uhBLk05/azlntq70aLm
VX8hqExxykihGdXIT/ysxfxrAGE3qCGF9lX2SvG0ubDn0pOWvJhrc/+rVmiuiWJ1
HPzM1Z0We8knRKvIXQB1bksnAnH0sLpPnliCo7B8x8yX9J5r8OgSA5tSnY71f/ot
nQG4NqyS0UE1onM3H9hU+2Qq5cgVyIQ3sHewxE4o4drcze3W0e4vx/7URG3/76Aa
H5w+CGgRTi53MqpbBbgwl4ezNUyOX1Sp3ZVO+SgZbxGvCqh7XM8BFgWdrk4TxpqA
MTEk93TSkYI29d1TMy3rkOcAdFUvPAtfIbcJxJ3gVTA1TiJqmLgHV2EbFo7h04q4
kgtvjs91yZMriA9wXlM6vwOrHodUQg7i8pHeMknbDR53xOaE/P6owRwRY+2OtrrA
fPYji7IgEv0wYN21UGgunzwoa+G7DPG2vZ8h8El3r/eZ0UDrBy2qG/jHXXOTipuJ
7ZyTgOWZfCY9qMV673CguXybjSML88e0DZ665HByB9IzJflruSvP0fHnzcRbeXfD
JDNjmgVHJL5umoMJKAr2Qx2P80f4OKnKMVj4zHSZ+LOIWM+szJtoVLgy+nRgoCvC
+BuHw6X4XpQQNa+7qpMKD/uWvED/pFyNqT/tCvNTSl8EBzyEfvTKIeB1GH0H0ocp
5naffLDs19tvFOD8HXVKVgZqSgStogR2sdaP8nujDuYZi2Ia6mVT51BPkEY6Tpnb
Y5nG6S1uTDw/udGhdg+qeH/gdGlmAPHrbvUjQF2AhsjPGi7scMN7RUpgqw6LxK1c
/Kvjg8J0HJ2FjsImbxVpHBQB+kMoWa0iZa0oBG58TNQrMj2KyWMXUJ6C3i0m5JN5
YGGp64MaV7xMRBzwE+bCrlkuU4T8cqGUOICtZ21T9C3G7KDUB2RHnpjK6o2DEYTx
7rc7LQYsmWjEbSW5hw8yWqUQiNbOzXWhx92x41U2McV8Yb0R1m+1W5Orn9pH+5gl
C9zwOJ5RR5NDTQlIXwG/+morFJYzQGz9AC3Ti6Mtn/cMS7Q3NsvFIXGAGB+Ts3tB
TTZxPDQ5Er358iC2EwdI69V+uK9Mfj8pJh0koEd69NdqPE6j2W62ReJt2JewicjT
3T/jRwEgj8LUL8uNYPSYB5vq7sEcvZHoiPwiB2IZ7aF7YlwZepDKhh5WXxlohDj4
bfd4UHeOiPSerCkTxRLjLnNfWS5tX8KvJMsq5oycA/T677pqtQKUwK//thNPCy6E
6aSoPBGVizTOnIJ5h83C3ylOqa54gIRugrSobwAXrxoad4ZhqKKjBlgLVjbMyIFb
NtoI+9wcHIksJOyf7HfZSBSeP5Y4kCdAlcVeGaO5nHHhmcLPuIpdlqbxqQ8yHZGr
0V9hzJvVw4HfKQ5y3MSq+54bCgdfNAaImTmQQWzXXqgXjcGMvP3U790NTT0Zdbjq
vbZS/SIqfus380QuSiUIb00AQYz5uoIjBN0Plri0Xl4miutnB7VRcN6oVxLLN3up
ya9zXtN9ZyDHDkuJr4Hdk0rc3qLSD34gJdB0AYXmkJ/EoK6uhLqGv+ZnDkaIdGZt
+tPOY5a6r5W3RDgfaHC+hS9qyF+bLx/7aJ9ec/pIVRBo7tg2bhhBAfyDH+K9hfVI
rIBINXlWNUikNN6jjlnmj5wj1QNPllG+ga8SigTFMl3G1P+jPmkgmZhffFC4dDPS
idsg93mFMHcFWwQDTV+BbFcArB/qjDCShAGzLTzed/d0HrdVBWnHTcLbJsYt12yz
jBLsPlIiF0ExbtGg2LEyiUT328HxyFfqrAL3weLcPz9lp9XzyuPkjTn7tN8hCXB1
LzsMPn9UQPBJ0DiwtS9qRbXDho6q7Ksu+uG1ETu9NLO23utTTGjbkEPHrwBSif6Z
tTA3aNWNHG7MU0/t23H1/Wgd7RkOimygb1jlV3Hu7Lp/5mS0cCM87tu3phMCQYLd
G+VudB04idu9xqEmKdeqlwe4Y/Dn3ykrupVgYALaEVkmEy6rFizC7QS4ymuAt9h3
TmZsGDK1oyQaPCY14GHHJSGbyZZLSzegg3C5SjRVZe+nlcnXcBve6d+mqTElCOQu
kAvyPP7gOCPPLCZQOHSNDRKRfOAs8YpztHx2Tm73pHXp4AH5du/+W3EvCO8xvdi2
oNM15XEc0V+DSrxdyCKZ0m3800io3to31xlI+YM4dJ6nNfMvPHg6k84ue3+hK37S
GNZ79tvEAeD4OxyYoozsy0/cQUImhDiJc7W8oF0qX8+sMwKXjWhHT1ldXT5Su7Um
NheXGCwcKDwA9SYj837uaCh211iqljVuklmDRKti+cfTTLot7QD53YdeskXk0wDy
MyPKwZstVLqnkFcuXW907p9BBX4T2EDfHRuB6pbT9wabSIp6/z896A7OAoGnmCrm
vF10S7P2/HLgZBWQtVWzWwdKJKlp1MP4IBE9QfsbUU9A6kfC0OwTMRo4M/jT8bWO
y6kIIBaPjJdkoLHUguRHClqxPPq6i55nuIIdDmBtYPO9NXj8wqA/S8pbhN7C8Dob
Muu+sADkyU0fcHkPF7+j39s/ad53R2XWGMG0A4+Fd7j21RP8WbRRMoA+wrByVgf9
xW3aEe5kv5hlliqZtBCw+nnfXybFN2kUXPCfAZsbNIzt9I41XENodiaTGRQ5luMo
h7hyabLv2RFDAAsH+cy2inEaB6l/Njo2KahFnz59gGj37Ucthx1jYsbyulYwBGNM
UHL4Jxh1Ca/UeAzjqXTTXvCWpWBk1pjTzWv4Llyxq2lJRPWUZUJmr9onon8w2k9P
/H0D1+JnFgIg4ONrWC8rafwKgmS8L/5jOXSX+eZZFWeCK1xcbRi+nr1/iRnnJ63P
U9+iVw1ndCWCMqR/EvRv7DH36LVYWYxtWVNEZMXlj70YV7XPSQoAmItJe10Abgj4
lTQLPC4yVhl5ceumA0ADMN26RUC07TBUpbO9fvBKONTHOOtAsALB1fE12g2wVCEY
lEgfl/eoC8gK1ZS1V2Qt50lXolIUgPfjgi4/z5Qb+P3nFphkI5lsDdjwpz85AIIw
JkGrr7wzDNwNJJPfK9HkiFSs1H2OkrYxE6U5A/Ep0bQH/3gcPlGKuTIgL77M/8IX
44t3FCkTzF+8HJpGgCyHmdpEkRu/X463csUsN/TCuMQk81loIrNcMkr0+0HPmoZk
DutI7qK5uju1IrAf1gEPQ4O0G32ww23ym+H8Lg5CHJ9W/5eWzOoktXXYQgSBRDfN
2sk1nIhhZqzA1S4Q2GPbKc+28P5ewA0eP2hEeDMfvk2oJ5uWGaEzIvsZ0mmgrTai
Dk54Fyp2sMI3yEx3omtdYZa4+jDjfk4+89xNhR6pwmgt03RzS/b44obVKSQHorli
lKIyq9pCZ1p97nKIk6nyBSa6I/pw6NzjyCrJZAHlp11a7K7p706y4NzGTvPQ6+Df
hTKpSTsprpS6NokHAl5rvLZLe6wuAdAiGBx657Cey/hxpppjNmRzcTbEPCceLJ+3
JTiXz/xXKUFI4e4/sD0vkyKynp7A1AigT3d3uQPOILQLoU0Qu55MVyCYwJ+fgdV/
hScHIZlv7rdPNSXgThbDUiqLnofxoTOUXimD0xwbwGYwMRfvwvHmXTC7XX2M9N5h
SVAbXYSPh2o3FKTflqVLjinsajmDCQKJZtlacNGNjC0KDbz+WM/8dS553mEjhqT/
ugrxDMd9hxCItrYztF8SQjzx8He4rAWHfKsWNGt+BnlrwppPxWlBS+p0faQYpeq1
K67jOqEnsnUGxvr5ZL9z+zg0Vn1DpyJkrOAWS0e7qchGYEwn/qgEqgkoX4fIl8cT
XrDMt+4YYnPdyjTt/2tg0ZPQybnTGWsjmWvdGmrssNpfXrJfbk+AE8IBa/sCdyi3
x5aqqgBJIK0XKx5taew26U+tefQnVHwBbBtepvxY846kPfW4PDTSJc9iTHTsz7zW
5m3EK0Wyb0L1Ms5MNIYHLsmD18rkgfbPPfF9kmdvYzHKHonSqngWq51E/S2qOD2G
YCaqC8jOJ1LPZLyYDvUUSDTqi79LNczr54vgJxPDSV2KDB0dKVQi0QEOKscU20yu
RoFAhYpFhyuVpmY9x96Q/JuweoJ5RdrzQn6TagPOJNcLaWpFcWDmIDvwHQQNctvH
+loYglb33n/iKxWosut8tyIlBPxVB0ir+FtOz/1Yhw4wDY3jjUkz8W5xrdkE73aE
5jCoowyhAaN8wooK17sm49Pw76flnEJUJ3riU0QnSF7Xgq3dN7O80ZhxpXPFV5dG
+XqU7WcSp0Oq27xnRMiO0exKPFFn1IeEzBkV+QuJVXJcz+o35A5iVwTT04xlFuf8
rFq688RW/wp+FbVBhXF0MgXSA2oxSZ4Uuw1xszm3Q1VFxvQF1SU61/ZeQWmkYUl2
EXgCsxo4antLdys5dUNuWihu5trrUvKtNtWrKFHMsFvAG1J2JjwZKtKjeWm7HST2
K9DEXF12XNECNbOX1MlBDygZ4FvRAgS+DlpjgkTXfV749gp36JQEVrm1jglPJUEw
EDLqlASQIWT2Qi2tj8BOzaJ7/MzdHNrfVn76N5kIONiivldbnjYKmHGf96jNcpV1
OFdwTkh9TAx+8DUmsL4H0CbS58N7rjL2xTqY2LGnljgiXDS/+tsdQAt5k/sWT4iN
OHa+QTrUE4iN8wCHOv+ZykjOF9zuJuMsVgaM7UJA9i7hUQU54K0Q+2+s7rYeA0g3
1xw4ZPSBlUnZRugGmaSqwaL5USPZy2vwxoH+1yc8qvT9Uzh9db66H7a0uiEJZKkL
DDNPsfqDdy11emTaiqALbj/p0KPFz//Zv3P8Nqu5rkqe5fzAVs5gRqvNQSIkv+NO
Eal6zyTrnzUdUz09mDnB5o6CP9Hz+LZdrW6CmshG10MMVeI3MvKcytHz2ID7+zcZ
l4B0WFe7f/ql20na07t21AsG2FdSe+LQ5cZyFW+F24XpCtsfDH/4e7l0sN/N3C9R
Easd1xwAuLWhE80i4fqh2jX5bExGYAFl+nMg5JqpgX3uRqLfgmno77pnGIE8GOCM
bV2L8N4RHDKmH5glV++YiccmmvJjKkcWUnap07ulA6kKQUaWvoTpKmb+V3KX6qki
7z2/wuAWNYVCqOfw2We+/bOyVt1OiQYuCmk/usGhA9Pg1BhqJ8eG5wM1lUn+zuPp
mdVvbCkGUo6uvwosbyCkRuOcRPkR/NS+qSwtVMs0kkm+OCr4wEaESrFkritVZ64a
qxpqTKrZjwsfdY1oMrcJBotgO7DxGSFrBj4UqcFREk+1bSaoap5r1FNxPtobrQVd
1Qq7TmLMTU5bTbsFlQCHh93F0ochYYcJQBzvVmyvFnR9DsE/1FOsGtsbA46CU2uU
MjGgaihgpaiNnR8JOnImpljXBEqrsqcIVq5d7S74cShFO97Pm3YqC2HXPG1CWfj+
Czod29ekomzUBAU1eEdlKX7OsYjF9s6tkILiRaZIzzDZ3VoMn84t9Rf1zTDDx3ww
Dr9L+SYUD58rXGNmHbAnYNhGKA2Ee4LCB/+a2E3cQbQ0YEORox3Rt7faJGZ1VAg3
lfOB6eIxNFB9PrILLA55es8PlmyN4CgpbSUOpT2qpqqlKaNO/4PV7Pah+UjncebE
5JpJ1yszhpqjJKRhokUte6PbPq724UfrKYF9zxGIV+xTLRckDDz6jwk/1aE3Y+Tt
UnABu9dCQ0nSPNfB3xtWpyNUbcP8HGDJp4Ij6ftuNKIEEfwU/4dmTl4mdWEK+eZO
D3iVHl8JH0ZGdWtUI8chfb62iisr7+0Uh3ifL0pnOYHP7wEmplFoPrrmBAQygbpJ
4ef/WGw3Q5o81o+dE57w/L3vAlY72uJ0YgEZqRlzbq/0T/RZ5IAVVW4e+CIWHtUd
qMhmMhmdT7oHDpJ89YwukoROn8QxB07Hd6V/u7MgcZYFh3AtllQmCA8I0hb+ihJi
TUBBNC78/A+DMrUMsxfKWi0YxcGD4AP/U6h6smHYcB6HP+o0p3C3nL3t1+RUz1iC
GI7t+oQVh8TwfryzRwHjuhtBNrmR6FdZqAaZAuY/fRqyBonamhEmcqVQmKtnU64f
QIlmMIK80D04ecb/eJNsQJozUz4/Xld1+PL2QCVpYe/vJ1EgOxI17h0dnM91T2zQ
cywkkHWMdWFhgtmilByjaB8aVxYq/WjxJKqa9i0aN/bgz+9cchQ9QXXz3moHupRJ
0APoJPqsXDlXpIMh3D3qj2+mL4hdC2ZfM37OMWLTTQ0IVJhdBBCgagxHRyQCdnwA
fPRB6LlMoWfTvSCJyVLEZqmTG4gFNbP0k8iTzcO8D1lsl3W/hvxUWFpglN0ZKsTW
5VKYKxbOxCC/e66KfU2vkxUxh6DUKND5lapgsvlukoPz+KoKWdsrR2stJNFeYRLg
zc4tFOiNUrQaDc4CPMzeZ5KDq9rA//snTdD1Vy6uslFSwBDNXuDAA9DK8ZdWtMyx
hoaJgbOl9Ld4R/3mUwR5YW++CQgdrLNrj+C6ZlIZy3ZqPcsnCfA824c0v8hh2+ym
WKhlR8iYywYZU2QaSPyVz/4Q3DQQGM0ziA0su1XPTv0AjgdjpiIwcZTWjjjzq8wp
8+mVjJIuJ0PAB94BNnGn7KwHGGVfgSeNxyQUqQHODdMRZhY9b9TV3A+Y0MDjHaCC
7l3c8554Iv6nHZY+DaObFw3g0uY/sSQIxyXRLt/8FF3ccK57BdcAtXXz9AZzeq8T
YUuEdZvtnpnHGnWgiy6iucbnEJy6FEdXrtNFoOg2eu3Noo+dr5YPFrQqKirUjKKh
ZwXtyCfuNl7Lm4VY7tOQK2HHqMfxKX4jl/FC9aT7dO+xl7Ct16JyqyACl6OQWcmy
fz2lNbjemO/wVIxsk6uKP2/sQ9v/jTOF9WX3JehiOxWMBOBsGBrTRHBYLJvWHukn
VIQOL02rUmOAV848un5cs2GHriAJHdKrH7n5KtmeXfBcFKKJhfIy7zU9qWfpk7g/
YGO9+1APUByd53DPY27LcbEMQlpS8rIjoh5jv3E86zrexnkVbaBcOVtiqO7z/LMk
2Hh06XFwIfDz0P7+QRo1zYhb8RjWQcMrHwk79Xkkm3ASKyITX0uBLeiuvh5xHDSi
tRQPNA2NQPf10nCQIITg1mtQzQgVRMGXl2rOCx25NNeJUADXtGV5D0JjILx9ccn9
10sKkhBFqsLPvoueUS9HuPE5tWz2rMckC6pE951P5ITf30YNBPDuWsjcbtVxpNk1
ZugizlLL3dzRil9TxOfRKMaGPplPIwh1nuYG+uavPRC47dttnF9WOvP5fPwSLFPZ
uiFiIb4UvSgOuq1Gkv/t/f2gVXTgm3jt6fjtjF2tjHo33VuQeUPza63mlAJU3yFO
/t16ZGccAVpayrODWp/V8qxjQXdUs0YmjcXKXy0lUL9+SJSvGOhM27qC15HM3qqm
QFQ9Bk9R7hNexDBIX0/KVlrbARvTG5Y5E8AT1tQo40DkPEbnsdd6YridaDwA0GhS
sY+uBiaWE+6rVHYO9rSqzMNDK6Ge+ydgBMEvjJL+4LvGlXqSOrxGr3y4i5E9v5pU
p97JurDLVVVefYWkrr+fZuhvk2OBo6pEIJzUcHfLWDh0/gGP+lKh45t6tUph0oSr
q4kXlo5CznOrNSN3Ly8HbGIegGOOENol3Vp8xt83TN/5HZgqpVbCHrhwPQS3AV1w
Q/fQyMgOcGja3T0NUYsC9kcy41NW6L0IGim1FkPUm46gByK5SW6G7exRekxgALvY
KG/QJwqXNjlImFu6h/bVkiQB15kachtWmit5gAknGLBIiGJyRDb/OztYNn8wl3/r
R3fU4dnlWFAwaT6wxNtRU+8BY5lq/VJybgfdRuFHPmHswzL+I+1Opui1VGqxoGW8
Jbqq0PDJxOM4OhJ9CcfE4ppwyQu8WiFM/qhH4N+10mm2gm8Ht42pe4bKY1V+RGOs
WIGEuF9h1s5sQorc2fwH0FFWxLk7jT9o3HN8INL5ZEJKGETnvPfWnPxdDUsJginJ
Qf258SHUP9rsSHSTCSyfN04LmA75f+207HWbbtzdLvyc7ZR3cbpTvEBVGL6XWFNE
CYOFPxAhOL+wit6sojj8jn5hjMw2KETJ/XiniYn5uYxVqrF0w0WvzxwG4oXoCnlA
mTlpqL+djj46mbLSGUsdel1lUcnfkdX3TVjF9sKmMiOVqdrU1OjJftuEug42zlyU
Bx1T+gW8Zy9VXTbKhMH8ieIUnfD3N2DGzFIe0I42236bcLtJrAfPobGVzTEiwQud
h87Dy4Mu0u9gVayaxeovS3novYqJX36k5zx44czdzL7nuSx1FBpbJDxC3HejJldz
j3Nrs/vuqvNTh7f8FAyJ4eONa4gA4KehkH/R71yMqeJaauomnM6H6yVSsCVEVSuA
6LQycOXD8RlnmKYiHFwf7Sn808f+mnrW4fNCL3yqRPNpinp0l3a8cbfsRwCdnhJc
wa3ZBX/fSrl5JKfzSRVevwH7lXLMz2w19K6rYDPBBSv1lM5aonfXwTQsT1nvkeTF
5sZ2nl8u0OZgWt1FjuDaNKfuw1LbB2QGqdjXOx59EfGBxI9xkk2P4UH4oR4gbaD5
luq7TGnsSjuYWUpsAEl+EzLYG2aFKJ5MOxFX/vfbcSFZdG9Uq7RUHtNsBdIrYSGC
EcKHek3pWUuZaIQLzW9w1aqcCOageZoiam2wwxhKYkLSjZRz2F9DWDDtBtEhAf6J
ri4m2BqfUoqL2Qid6XBcese8c/RDAdyMFhckj+nqMJ3cSBpg3aTNJroa6c2h/71u
IM2A8tgSX512NgUUlBDh1VKp7QkgiYF45ABN5DVO8/7Qk3EE7hOyEPuFxE2bZ8kB
sDk86SmdjJNecwZbwx6TkakNJyJNk/gdaQ/rpr8yGfOvEM/HvEXqmGbPuhN5/xL0
/KJYE+rOCGkYNt98xm3DySF5trRzwCQzgVWYPMjfSk9o+yhLb6i/9GlLJH+WXISQ
z6VBIfF/ikplyxV4sSnoU6VhhU6HR37JSfVWvMuEEAI2JYNLJmzFbx+ONeNdAX34
OOrYoicC2NhE6X5mqAZX+VmdCH8oMi+1ETgc8sZA8vUVYgQdO6TJyanAh6HQWusl
lldqvzN5w2DMooRyMlAnonUSlCEIxaGZazBaiJS/IxeriUTuifsOKcMiGy8czwtV
fxKyRXN1mV2GCoN2YQINkb1AKBCQWlZvQTpD9IO2Ef5qqxnDO5Zbqndj7vmJ421g
47XV4nRB2vw+Pj/6fRj2EtQfWm/YZOdGpnwvcW+ex7DXCCk7BKbsP1vM3sq8uRJ/
SYT4484tIci8dBDa5ZnSPzzGfBQ/OOMCiHbCD3bI8Jzkzar9j1NuIEBzsUrfB43I
SSv3wudUXq4fIdKLp/RlDBMyN2aF0PQzi+ge+Mp/PCK3XECN5CTxbYVOPT6rsyrq
0YOtq4YgBG8LtHuZzQ3NiE35GRg+5b6TjzHe7zC9wcmS2XLNhs+DYvHnmKN4yoEa
pJFZTJOMBEhpwGgAJ0gEicV2Sg7vGlpW1axBXupJh/6KpTg6Jxk6MkjzMXyXqDmD
xVypayy+Sgq9dzotMqa1sKaPL0IwwVskUO8PwS7iQwy5fJC7eEn4cnEJblhHOXof
97Dg+kmQLY89mOO+o7NKuh5hsJHmK2Ni1tIhEfZvvYN+jrfmqld/B1a1iGsSCVCr
AvDT2GWPO84PSyuOk/T1Sd9YnQGajg+wdvxZnj5nV+Y=
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:18 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dXx3V3oKkuuBvYEvGbsXabxlqkTeJs/6S4TBvvj5AlI+q//3AhoeudPl9CMkqZBw
MT4hdu9Xzys+C7AmmiUdec6SvPyI26/o+j3tebIP4gh6Xfo2lKV52uXTVL7xy4bG
m73iNhx6IxuLKWEbEPiMqbD2hhuixkmZdDh+o0MifuQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28528)
RBGR4SIyAbhsUzOeCvls4d7T7rirEteiCoI7xQQaQFSmb+SN2nc0X7Akn1OHam6M
C6ypBt4IGy29EQMzFoacmVnQ6eFihPul4LVk+B6Qju8j1GDB5ooeBN2hey6XtE4Q
bHFCgIllUdKvF9fQFjVNLq92VWIVpLwE3P+yQjxIJg4l7lx+0kd+24T5JRVQaJox
QvqbcCvkJ0iaLZRP3OxgLgTm7WZXzu9RpkbQ5dHfoRB67njDBg7Mcsykb3elZQvx
CnC4Uc1ii9p0WgFX69l062tnHnIArqUzHXWgVLdYyfdFmnDDZfmG979lsYkM/FV/
mB0OcE8W+aRpcrXVEQzVOTRxszNFiK5Wbe3bD5iMQJvRtI62vYsylK+ztLeN7/4G
m+IzMscbvTpYeMm12Vwu5Jm7cW6zIojUsP+88uACJfIxDCoJpDST+T7qmBWFe4/r
ffjpoJLiFMkMR7K3cgjGUMvx5p330ggzox2yOQQlxRaKZoXW7YiuXzLUMIYquwJZ
8a2JLB5j9BZFEM5dsHoD3H6CXHqs/CS78eDEg5buL2XlTcOAeMVxtY6Nui8JirRX
SZ+BO3vsaa0YAsoWd6a8Ts7+OlW+tTreF0DO0SjcUMasCme5/300sB8J56E/SNgY
eviePANJBvud9sgxmEastOnB3O72EGgs3TJ+yEXV0kfCVZossPJcLgbryz7Rt3ca
9lzFtIk4FOuWHkMpijcr16MqwZ5gF0aiGB1QW5DTu1oBUWfr0mNAKx37hik7lhWY
aGYm6Tcxh+nhkgHhfYQIdHzjTzjSzHvWCY2qg05MEW8iakWboAa4rkmLd0eFimMx
DW3993ZNKyU/uswCulS0k+pFucxHUzq2wq3kW4psBJ8KqWTXWub4/w6cVY6vwcZB
7iZwdBfi18Ha3+6ozNq6CwW4v9I6aMwhqTi+2/kAeD/f3aMNSlRYyZXXlb3vWG8C
owxv6EKdWHWr8M9hOJJBgPJE7jNOqWYl67Hhg2ix6X5H4j/U+rm5eVOWT69LZ+wR
CMoEzCC19N+SrYj1S1m8HRKGtdCIw5BsxGyfB0jIg2c2iYjCIFu+ntsQ/AqFwprL
629n4gEFy8CZkU3SoM9krAxwzyjiXB4CUiaQQnhWw2OscjjyUV/ZPk1B2viADnMS
znOymWTor9oB93SRGkV39oCG7lSxacL36H5qJ1qjZGshyeCNBHGFPsNVTLU/8ta3
mzd9tB4M2ctBfksXnZYCCF/M6ETod+OHD1LQYYhATfN6qByI3duw2seOw0OOYV+Y
TtJmK/xMtzk4JJ/boYWQ9SbDa3v6epHaYf59bb8Uk0mh+l6zUcE/KvWs2Rz9/DqX
m8cRiRe/ajIoDS2R/hSTExzfPTKAYLFxQ5Y5Wg1crR3iF9bxfoiDhYiZuC9oqdao
0EX2LhPykS/EytpzUgdHmjEbHiqeMtwk8PNUnUEBKhkwLHVhi3RhHOEJ2/3xoBXU
u3K6+y3hrEYJTOexb5K35NOEYgaTbJJaQibJWdFSodkQM0P4PL2RtJ7ms7/wVqTy
Lm/IUClycK4Whfgzz0mtreI+1Vqm8Q1+GcSRaza9gUlWzQnMyEzvJRq4CNwy9KK1
t0XpWBrPBSXnThJXrGC/QiiiHJ+UaUGn11gt8txhNzpr+8WqDLSGeEo+d6gjOXLp
z0tDTM8O7GfA+o6niL9QGaMFia2ZQDrtbxrw6Ry9DdduBrBoeqRrZMVCrgkn/+w2
/DxLQ6UMT8wtaHon6v8so7lxXV3C33+1PJKyd+7MVJ28yMNInLkqvosEUJ8uXcER
hj/Ea9YfW0f4p65fbLYYKjojwKBl+a61oqGfhgdINUIpeDEzwuDbBj++Ne7Cqe8s
FKUOcPlp7UGrmVQ8lGwJp2I25KNR3NLWD9KGL3cZLMQzTtcs9ZSt4D/0RArvbHoc
omRrsAsruWBSYHf2icpHxTq/0wwN4HnvQylN2eYDRyzrD0oFVPLIPdBakIN5A5fL
A5Z3CCWAzzF0J2wBzCcvxjA8xKEQZlxfE/xvjOxlUKG03u3XreTy6xTKUTSxJ4NL
BzcWl2FiFwkEQHRTjFgly+pkaaaWMmgF+tac/n0FT88ZY8STigtAl+5OFKOkBBp5
zcPXoPzj0CkPqH1vJuJbExfkTO/TCLGqRhvE9de7Wj87RYM9OKoww05tED1J8kSK
OixPreTEUN7EyS7UM35YT35yiohEHhTL6vtqlhQJJYoWXn1iiKNrJ38TMRuYU9Ve
TkISVsZJr9C3OtfmG1putPHBo1EiNADYQSiKFrhFHtCPL/eOdz2wvbQBe/2jnIa6
YeM5pQ8Ld1Y42Iesc46Gfvsq6uUgHWPIrHFnRjcLCFSlhxnP1KwePz9rYWAbKzXO
AwIOW2ubE0jUkJrZFA0SnCuuSqbsl6wFaVfAZGtPNS64eOEHpHPraWYNwbkwO3Mh
ETkrGLZYBSRZqmjnTCq8aMYIbMr25dDW1UVUtUP1UHpWI23Sl0jLzF7kMnj0ANo4
bhoe2Ud8zVSgd+YBBvI+HW8CHRW1lWWvy3qvM2OBsGsSPKxAJl79OaF3NLF19ES0
I/CUQ8CjiBzO+kOzePgfxitd3n9ULPt3p7goEmwHZY3CByatdT6Gyn4DKepIGBaj
9H65bKhPmNPT41/0fyJZwCEn9gHkM1u1WxIuazwlS5sM9Q6HV1D4rom0KxAD4Fvd
rHg5IBtznt7DHrhOSqhTpO+zdZCLZgi+gbVQUmxrDnBxr4Y9S9lMcfJ4gK+PB3yP
Ciw/c4O76T+40MWP6xsztryOZVRIP48oNxn3hizMEzpnMW9T4o61hQBl9TpHQBNn
ZomWh5TYNnOmNJxtXUcFaeF0fkEArqePVoUJ0nsRLuwyD8l8wjJ7vX+qRJO6Z4Dq
tcYGyRpOAprmhkCuiT+CitEHwgzc+Dx16d6ps4icAAneFAdW3O0UeqBsZ/OySjxl
/I9R3GX2jiHby/d9B6RFuVuT0HgJ0C7K43nQ9xR0eiG8d6emfJZaJgDI5N+Y+9ge
nLz/hqyzUYwZUDQWHZuI+A3tdMXyFg4VA47HZMkURX6LAJCouh5Dvma+mtLERTfS
StOS0HwI0Te36izCUsUX9wyhsavI9TnUwvzGh1EmRU5LUyGoUKeoehFVzvHfqZzB
1RzvRjV/CoW2G86Kp0mAZu73FdB6PF/4sjhikxmGI8Kl5XD8Sq+5hHEfTDcAAp7w
4xRmkvHH8isbYb1sGpC54TWBrlxpj3UzlKuc+Y/FCIzX0r2EO4vgjZ3om+NtnscD
iPscco75oa+59udr6zS7NfZRn00fmJrr3630sBmllTZFaK1ZhOsdsnTp+ufvYqeN
ALRv0Jyy/+JgaPL4ZU2oB8/dWNoFlbjpXWyicxuXwBMCSQjCN2nDNe0XhMYIw3Lt
PMPXGChEWX/wxldFT53Ouc8moAsXPTgMA09e1m8uqAxmZ5I8lPkHeECPXc3CLj1c
4x8fUv7gqvafoDy/uFTXdfaGe2iTNHvij9LQ91M0KWAhLwGXPnQ54Im8bt0Fg9C7
Wm/6jq/0TUnFKgFk2hpykJU6VUbgTfaZrSch7PdxkXNZFksJLH3D+HDSvV4hZzGW
rok1Pbqjiskk/4RYHUGIGHCipPj9nPlXVR3IXj6zojjw+/3fQaw4XtqC9K84M3Lk
mETKtkKlX3eE0x3IZy5foV2h2nF+vJMB/NGh/Ze1301eIoS/AdYXCDiyV4r60yIG
hlZtoAOSAM3am7bbApgrIyqXccpPMGJoRJbU/DGvaaJVyg3/rTaL5BZJZnYGqXfV
uHqN5JXE8C/PEwDNAxbFWU0h6avVmFu/8iHh2ThWyjxjmLecBn/oZouOzoUpHc8r
rIpNbELnGmecaEyN9gzKlanhSxk2cXf3Jfso34uQ4WU9SuJiZV1y15PweCGrWAvZ
DENjLJoVu+xL4fWYWuvTovOc9znhkqmC9CatyuxHgqd7GBC185eKDNEIzqldgeAH
6MpLtgXhacdyDY+x2z73HTDE78BAL+iFBjklkxiAL0tQdKxnpgip+l4PZlpHpqC7
0ih29vV0TTsLpZFlJUP1oRthkAt1Lnw28sFXUf7dXE38wkspEoy1AHEIN5ZywSWN
tqwQoAqqYRPmrUugMi6Hlo6FEQZf5PoK35DcDJ0z9WYSlJ9e1kgeBREdwxfKX5UW
X8OVWsJT1MWsUBmN5wIzjvPjACpDoLRzcVRJ9x4RH16LnfTxvm7PHxKenPiGlbh4
5GjvLuyYHlMoTWbn9THVRvKgwEXWJagFktS//fDnujXph4p1DtztDz+wiWIM9s36
+GwTCAV9e+ZxbL8TseIoH2mfrYZ8tQOyPWiLqEplibHudIPBukgtsP7bOaVCb4ap
c7LTtInlzq0+HVhG7XKyaPBDqk7vJtPhSI+2PylSmmQkP0PDQ0eoCpyzz1bP8UY2
+mn8/t81sIbn1gv+6zzeFYcxRng99D4vHmTzryk3asz+6PnScEZHyhUOZX1g/lU9
/4X9fNZt8ZPaSl2OO5Lbb5CLSZoTUDkr9jUWVu4NycsfYreHB1dzcn7wt8h684Kg
sq9FeWKVcUQuHuEgnnX4aX0znLidzBJUcUkcx6BfQVgpY1pLzB5Slbq9wia/Qdqq
nXS8JPxGpRcJKhwEWrQVYfOSyiVDVgRiO29SFoSLgzgxC3psnLmYGLt7RQlTiA3m
3Fu4mlINn9zQByMRTmZK+mNgLgI/tsbZSHtDP4MycVSa8hpVwqbx/7/gXmWmjop7
9mtC84hum5YeBWt75SmQPkPScJBxaxFOoHclfXjbu719cr+kAdTKFKq21ILjXplx
ZDZPW6M56qd89fAAA26fMIWipnaXkwpAMHkhIBaT4OMrXzJfoEM+DIdGND4VNpXv
oYRFefn3FDFWmVquuKC/RZwXZGlJ1qx7lecXjJJ2zGbwBcfhXuAr56+UAUcS23fM
il5AhpeaudXJn/8satqGdXNzQ6/h+yN+jxNatGRZkUKC6Z6R1jrKdnqBRtdapXwz
9QuOpfTY+D/x/pcX4R5bq3KY6EOlhCtDh2FrX60cvpA8QWopRPHZrZYIEzxkavFA
WI7LYm1epdXZTf5oO8PxKt6EtuXGlS7X9pliTQyDeWW+npyhaEYvI3gjIZTwk0BE
izsvkC2/Cx42Npnn8erWdRanSwFUT4wAzpR33ceaKdYfVFwNbiL2ZPzXEeKff56f
V1FBuTjgXYvnh1eVn2cfy28FkvhyqyYylbDv4wwAY2AV1L+tRKbeAiaINpD8QCZj
Iap92O6wYDDafEZ9RFgD6W14WhVHRVy+73BpjCJO2ietUDVIE1dwNVyPfnQNZR2S
7xTIdQKm98m1X7YT5a7A2Dil3NyD8Ui0v0EHlid5Zaux1SW5uyA4HJQfmt2loyvT
Pt2KptPhhCK56GFMgiND3m2CMF7+iGolI5wBALwqywMYzZndV8r7MG79AeU6ZpYW
H4Ye2Bj/iT+EKyFDqJIvrYkS4AR+5rx1XvYAWL3RM9KfIlKjck3jNvJYEo7yLXBF
sXlkoZPjynW2Xoq+Rru9OPkM8DlczRH1bkPiASv5a0RaM/r3B7JI2Zr9Otd0ZGRQ
QrJSCp5zRF41sRBuMDvTQ6SJe538Hc0EsggIFEyokU+L10kBbk1LqeOPQlDbXaK7
QLdMRWwY+UXDsWDRaFJaFsd90wAK7DrWqPyNVcIxUrlbuvxQKz8nxOtIU6y1JEph
8+gCoxFCTmkv3YdleqGXnbTOYg810AfA4hyoCkeFEYq4iDcSP4mc33ERq/vor/UX
q6jHC+pLcqLuxaRgamnHBDal78GSg3/f5ZrmaTG0aFB9Uq7/Lpf7sWCYeGcJGWv3
RwdtU3F5FRbXD2ly3Ay/S5dHMkowYPe9qvscCZlteA1XefkrU3O6IYeoWUf8G0Bn
nqaGqQJLBUtJYKzmUi07gSCxDTrnp3tvjPawW0/yt4j6Wf8E7f9nwRvmd2RfKbKo
QDm57kFdZqEi6IQdjd5xIhjjC5R9KOBQ7AeuciQwoRgVY+l0BKAt4gYMh7aa36vK
JTx14wImaQERmQ5zVZew40v/c6X7jmUM6HQN12iw3BuH7Tk9Um58P2cLHLTdaGyj
JMrDJTLWpHmijYDfd1nc+GO5IXzIeqgL6JCS/yQIf8P2VPJAgh+JckMPbHnikwtf
31V8GvL9IjStNjdP5U1H5iRKorPXgnx3qkZTIUiPXz4qLGxFW7HPI8mGYkodTcpP
D4p/toZb+W8DhhGbYBY86F7NdtHK3cY+p9gkLrCdoTRFNAsCcsykQOcXurrKl5Df
oZ8iJRzfbQ0jiXD13BB32WTYGmqW+he8TcKAdvCxJng4V4/8ugHWjqRocJeIOFQK
R/orDpuBhaC2j0CnrJdjWF6aHFK4EcwUjhtzeDL5tSX+4OSWwB0Zk31mlx4Fa91L
+97ni0Kv/PCjKPJE+hKqUenXUcmNqS4qKNUDLfIVpo6YyAdKdrLDF/8pPlXX5coG
dqBWN4jDON8Vn9Uw89nqj4US5GzulxoWPQNxNastvio1hrS8CeNB/oO/N2ybrgml
2MlI+5ryJYCUCvSlUzkcgbjDpJaWr7A5hfReCRzf9HL2mfOXsd8ufVsqFOwzp2Vn
yXgOU9oinGbFEa3zczttc24qtB7MowIUfM83mfVhGEJ1EFNQpYljvan6rzVaPR35
0K2rnSyEukLiWMr6kqkxLXbZHjFIIujscjy1t4OP2LK+yB21Q+kkRABruzoIr+6o
+U6t2gB1NugN66AwwGAEhEp9vdnx+CFQWNaUKIOAft+SncWMZ9HWXJQAc7/vEWaZ
MyMGD6z6fsX0nN6XwtE7CS06lJWlUf9tyAWHmF9vmhUMTwGJ3FXsHPohzOcy1wld
TQ7ERVFYXXxJhS6uJ0nwBlO/4rOVKOeD+JIcewsqVgrCGkxsfYay6G2aYVMttUwt
KctOs1tEC2S+tQR/ArHenbpzG8xa0jIhT3bSlYa06NEou50aWWstkpSTuaB5CQWm
rUncNf8dfuhhs7/gNM5GvWfnRqhNpYuYzT/G8FTv9h2joTLaaIcxiby2rrAcQFH4
VXfb+x1+X4rfuBQlP15vkkMrm5FwVwemRgb5Q37E3EC/a7X6/vqXW58vhueGQv1X
wPMytctakmIpcL2pcWxMMgTqpk23BkRihEAfQsAf7TsPWOp66vRlbOyXr411P4zE
H/pUbxIKhHO6+wyfbXLeoiY21AVF7c5u1aSwSDLImVwHBeJ7RnSEimQIwlkAf1IS
VQ6impx0y5uoPRGD0sJ51zx2vA66AOYMrvol6fRurQl05aJEm1Yxytk7O1An2aYQ
txLpZnwMRr2vPmXQ32mK0gPhX3pKxKmioticBn708y5oIdo33lTmE8pY7pedpE03
tHgjiBAgzodMatfQAtGX/tdxxWINpS2r/BZwiepOY9qbMvG1zxyYCG8SmQSw1ayE
jB6rpkbJbvvgUT3eGzrHKeRO69De2hRr8IGHRxEtCdmbk6fiijVvjp5RerGKOcY5
lNRZ5eQObYBKYKeUZP4gzj6aj5dhXzTYPS0LdqEg3aAj4NZAI+r+JxyT5NcyB8R8
9yB3S0vZnq80eq4aH/pmEITL3wujv0ti75eh6Hkprn+wfvCz2Gc4imNEG5Zp7BX6
5Vj9oL4ulc1ArQuhwR6WFuoDjxDjpWRHzb/hScYUOhDm7VvqPok2VJ66yvTSMFCL
5iYi4dM0rsD8OBT36XOuz3VQugRljwCMwCLT4sC2n9nZgHlh+WclYc6bUx29zWnT
zDPdbMMZuXVPGpx0Sph7b8yCCfx4HXYEtUUhGTZj+mJtqSnXBfJoXyYMn0ME3oIy
2s1Ev5wk/bSBGv+MbJMjQfoIKhoqBBlb6ZVEzjpyltcXMO7OWiDa2I9hDQLZnEY0
rv9WFTWM6LibVjMENkD3r1IxEhQtinaB377QCUqyNpMW+lFbFt9hoRX90lpbM7hC
Z9WfqzP/G6D6/xWvXtZTQ2RpEle4RbLt25xNLyNcjvSMwtQs4iHQBua1FMnm609Z
+jE0cDZ0hkm6z0kIHga18Xh69j/uvEtCs6QLjzul2RZGaUHGVLhQR9gclcS9TXVI
wrDkF+l0GX4M/zSvWY6Vrh5khzqjXycZfkshKn6COawqsY86hd0UR1Bwy801/JS3
MuRDMzwQW2H9HZ7/Nc89ypN6HMK75dcgGN8g/eHltxRKmGXx0Wh40RlFMjFRinkq
8dEjep+IErq2j7PLTN35P7qgIZ6bRXte02GQSg6GmIuhJOtnJPQRC9TqKDTGfnYW
ctMq2q0YoCrd1oyaLk2tJrxaJPLT3XNslp8bTbdyiXkWe9QJ7kVNnF/CmL9ikzoN
jZJsbml+ZzDnUwqkZXjyvYLpnX4IS9Dda+NZ3JnlHCGnj9nuEw3BNJa6I+D6VHu+
Xrf8+1Hdd8Jun5ve8/5tLamVvjgTKXYVdKbfGXtexiXIAmFxdQ0C2U/Yqp7rTfGf
uAV3VAgv2MEC9vAzz/SgZvpgrJEDLSevY6EBCC6J5VR3LTt0Go4q21Q/3/rPJqEJ
6hbQkaMdpCzsARGEXfkOqoCQ6aihL5LrpcTIZrL815C46VlrhTzPLb0UcQ8L75JG
8ni2n04dXN/77qJmt46jqY3Jqo+oWWgvg4MUuix8B0qjUw+ywDlLLR2FB3zN0QJU
fy2/Uh0WIgru6zuh9DaFbgomrRp0921oXheBHm+RE/SKKkEZDCxvlRCJBcyQ1U8A
f2utF4qmvsGJYUvA4wWrQDEoT/rhWUMqaKQ4HSUZ2wWcfaaOsfAGCYhIzm3HaioE
eYW2Wc5SLl1+nkv2hObgJb/tdalawLH3q4S+Tn0c74t6lkrk7D/NB+xSdA0doTJa
2UmmpWy6s8Vmj9x3joXd5mZGMYmnyW8K4BzkXDzHhPMiU8fYWHkHVLRAg/WXyrhG
gVbL1Ktb/nMOFtJztjGjGY8i99A6U/HVVFupAQUF4gxU5Agg8xL+pv4v57aawKr2
ieHkr4PomCg+CFkkO7nyNzV9cbg7ShpXvq37QVKzmm3DFKdvlR6XQRN7X3Q724Ld
LltFkEWf0LOZx6sdvkrUacnkhjqHuNPi8QCVk0T4ItA+2h2UfHfCO67tuJXNCKCI
b7MQtXsCTGDcUFZ7fRrhG1d8S/vYden+R5Ilv6DE1bTNuEaEIgvsv3tIrPJ3cogH
xiETK3LB2RYgAjQQ7xYXIX4z4nUp5rDsWTd/MoXTljUgToNAR04PkOX4JEHnmbXV
NUzbsCbvWEAY37cNzOHEoT49g1i0kaEsadyad/U51SA3sscVujcqMLvI8OumMKCp
4mRcdHegtKZ0JCQgZW19tfsKmQq13D9iNL/iwe188MP0W3p/Y+n4lv6YptfhAd09
JbJVfB/1ipqKXtVCPe+5b99OkcFZH1XKKTDi1EUZNMpYnQVvs54op0kAsP4UVYcH
lcu6Oe36Z+pZl91mntqdYUHtYJj3JW1a02AXHRQa1VL95PFpDhAYPbM2AUkVTQ8D
Wo25F1LOqBJxqKrZwrViqpE4Y/U7UNU2YMI2Tw1XT84J4w++G16SPBxPNfyVMJZ8
TL+hO687QTMjU6QyruyxJOfE7ZvtvyiaXWoWaKHLfWQHrApbkvFQiTIjVzYjFMbH
px+4SJAzHr0Qp2FPKDThNwhxVQhVdm+BSJvySeNYszbv2IbWRY8Rvu5IXMc+JYwb
RG1zs1wCphPnqwxyahFf4pkckULStY6Uj7QJ8XIpYv/EAbgK0OkF74xpdpm4AUH4
M/MrZWt78RaH9+ARkDh0PEnWtpyKY+JRNvrQ5JICFkiY/Pv4mvxhQasNrO2fve6X
hQY5Gcz/OAGrg5G2rlIAgw8eCGA2o5asbMzBb1P1EQwzce4DuSfefwBYETplWhai
3FNFY7ahC0+FVna2DTwLEdzx2xXbDnPhn3FNqYn5SU5biDBfp5uR0YHs4DCk6CGQ
yOH7rBb20B3Uvp5eRuRSQnuXWAhGDO+3SukFKNAFjuQ5fmc7tgAdK41QYKJC8lGS
Ho0FyjG6DF8FDmNEKK6aCyVfHnBtDD3CryY2nSxsxNkowbSGDWCsnSpOG1B4TK7q
DSjxiNYiAmvyxb5ryB78iW31cpDYV0Fo4T7QuEP1TiGJvah4uqbK2dY4w6yBp98D
7WYWIdyfggtXPm0aNEw3S8CWS5m00ZjgD2dCFlic+z5UZG5Qaz1qUQiYzL0hIcH+
G17uUtz5fN1EUA595oJLtcZhIL6cKIv/r7lankXV5JlPlRdNkhqhtDh90J/o0HSh
WPzST85Lw9DjYm9F3sGSZ8sAIjY2d2wl/oSqsxhI4opgYXtEvToAc8pcNppQZg9f
+HAt+JDWtsZC9+rF8jAkH16zxzfxU/lHTz+8iAO3KTrtbJEs4zB0kFGU2grMcq5f
XEvvaCbL+WHrLOTtPR4ampUywvZ5hR9B/bc0OJyfF3+arCsAmSVfyzw6DWEJSPDr
t11JT2B+omofZk5D2C+pa2upMUtp3tWKL05kul51h0fXusecCKqaOrsA0FUPixtz
zjtTjpduDtKBQt4yBdihLtEQFS8FuQZTTO/S58Lmzdu/b9LzcCQU1VLo1m1uV/3+
7p8/MBMHhCaqjBQHXzM41kvpkI5JNBKk6ks6nEtFsnivFq+updILdXapYmydgOso
FJF1Pz7q+2bGBnK8ZANWhHRqXiJ9zfuXIjP9Vr3KyLGxPX5RSdoWEBkrEcmmrtPC
ZdGWGKuJ5mQ+QmYcUSk5Vtki6R8HdgOELQ1XV7DWjnmLDrBW+4DXwHG8om1WNyA5
Uvx55DtG/BrGAPfMjOmnXMK87/7n/99xwM14JUXGDDZv13ICIr70IpC9lwXRCDbW
sDuvfUyfCc8T9GJVp85OmUIYOl+Q1eNX4lDJ0IcXjwC6D0h7RdRO+Z80XKnTtYNt
MbgNVtit8dS4SspuIVIUqcU4y/qwHefK6sWGyt+MHWHuddNkPI+7Ov/icyliaebd
MMgIYK4vLir2j7Y3Yv9tU5FQ+DNzoSSUNl7gJThNiOVVlhwd4Nmnlnj5VaL3FKuU
s6fHeNqJRd0u1j77r0d/X55vn3XWReIqfJgnNLhPshZ4Wxld7Uwb8+8gfhRBFYrS
GOUjBRubxSM8E1IuJnlz/VOTyBxjOY0LLwM4p8wz+5zIE/W3Tt4g9dOR1ZbPIxMN
CWtuSqx9yrOpJSa1xB2ZwSX/OuU6vyKXqmi4LfwelNNQXY/3ePNsW6ypk3MuknTR
dg8W3ZJ3x5rxVYftY14I3L25T7JcLgGFwEk34e3UhztK7UxOKGewJwx+p7nhk4JA
Tz8BDUUiKUtEE5AAgGJZd76lPK5xue82uVh7gh7GiucwhfA6iIKAuMdD2o+VsDZJ
D28JyKh5stoHd08qbjtc2EO946MXOZ641uLR7UOUujn9sygvRwaQNabXmqsNRIZO
l0ZsohIccgAL3P7KTY1e9iMS/uJA9Yl3HbEhdG6XEOTuERXn18V+D4PRR21z2vUP
Uk2B4fta9LPp+Cjn9PTYPiJBJXTAMkutg9pK+r3JAXTrWo3HVLxXNA6eMkRRY9Zn
p1YFdkXOieqkJtiaALfLuo4JzrQAqz9khzYSWj2/+J9rXM518Vvx0NCods+IkrCR
1JNip/7PmngkmxT2cobQa7Jr4yc8DbHfu6HbW5lwBAm76hN7WgcLepXlhXg8mhu8
dFTX5E5PBeLynf5C0rhvRCLouilz0g/18WLcyUMR7Kp1hgetPtu41jItduhYW6gD
OTnrrpE9L6htaMimVXEeN7oEKV7y8tn2DTKDXfyNdki4ZJH5Rw4yYi8YZDkoYziU
kfPD3UmVKSTU+idwCKsEVhOb9Sx04Z/kV2Qi/PZa0RDHwtWYMjk9gr8ITf2HoEn5
veY7j2EkL/0QZy0KLZ+7571BqY4eYUcZarLSgYsIhdBUXwplp3/nuYJb2a+x7LnK
Be3HuW54diIPdjrIkYCtg3ZkDVcFns2jDgOUuU8aryIh17T/yhfELhjxp3TixkYg
7SZtH4HMDAX2r6ZVnZgRzc+TtqMeiETo2QmRvLW31dQdqlcTJU87xHFbFHEu04eu
UDazj0Lt28YgNWTRDHZ4v0Vm3g58mqLxF5FofhOEktg6pCq4eqSMdxkMRaSxv4TN
QaAQg82D9RomDNxiIOb0ucQ/mTE6f9L8Zcv6ZQhUCNBTblspFqlJnnXJzgzRBKRk
xQtVn1ojnjf2Ld9v/133LVRl8p7SiDqfcsQRIl0IJ6ERUQEGV4PF1h136IN1uAHN
HKFDupcLL2HDKyK+H12UFQx6uW5FMGr9yboM88/SbkXs/GuFlQLggtnQTn+nhQ0F
old0QmeoivkoXZfOsSWARrMecPZZ3+mg1YcL6q90FH+HRuOQ4wLDZgU7LBfiF0G2
fSyvOrq3LsynFy0MFwekQ5Ot9DPzGFuFSHiYbJw4BQiW9d+y0lFFpf0NF+bjyv1P
LKrxR/k2GMcDUQVj/ZKddNFweR5PtS/lScazhMWMfK27wL/OefeMLiqPyv5KDdCb
/hcN4Pm9w3blyGW2M7fPOifw9bkemHeTHa4FBeRIqbd60d3mWNOlHUOYGlYezgm3
fp2tFcslcZ/ZRqhtauQbPe2HJFvEvEueChFyemobSrmUwuXOrz5ZLOmdWZ6ivA2h
03In8SWjHwouQsGFZEpkD1h8ereSE2JTnfGdL9jDL1+JIJrhFwgEQfnnkCrKVRQs
x0s15OvOmtRpl+xNH6r5uFFeaantYKEJZpLnipndN1x38mDQWJ3wR85u5ElXOiSs
Vu2EdEGHyavUWWFhPiAHou9A5Q4w8u7Gkmf/6Z05b6ibMIK1Ec7UaGXN88QlZO8Y
Oth/Rw1Zr2w8+vjCjJ/PFotVjC//ZIbalhKHR1rZSLHRKJNKzIJhGOS0ENahKHPL
md2TDhM7L7TiJnVRoBE2d9rXPZaZWD197qKmYtm3vPVq8YTPs73zw0ICi+noohrQ
VeY8WyRXnd+Q77Jpj33OH3E/b9b885hCO/3evroBrzMPQxCO7I+HxM/qzeZEcKjj
Ye3vgT9YBBV9dwqK739PayzSJ53fod5lnluQPHRutbuY/3KHDhEiommYP6XplD2t
2iWJn1J6h3W8GaBQmmRUFxKvq5a7cm8rZPP2w1niG2laT3YAZviD1r7DKd0yYZZd
osrxLS4eOWMzvZ00SrX8Sxdv4jkdf2z2ipZH7sWAFThq2A5B53P/SZsPFWYrECLr
S5+qjuzn0pI6TUHzouh4ThlZv4GrnHrFLl0XcLW3AkGT2mk6Ztv+G3yIrUKO7JuR
Myv7WipEfsWDdbDxVQhgvSMjTFxu8T4Tj5ri/YrsnStTkO/eCpPK//mjMz/ODXuO
a4VVjKJr3DoFJVuozY8bPvSdTMT9XOPOmzZfPehziLMgIXvAx2VIB3D3Ki7b8tGV
aM2lb/UTtDKWMZ6G5pWTMEc3IavIsu6pUe4E/5kBLX1AoYB46dV/c7td0Ngs2EHU
FNSmr2Ua6BzWK5Nt1nWK+7xFdZG8sQFc6fK6pMqrVOCJ2b4km8c6nX7NimDitZY4
pryPDAFRivO31LfVvK4CsTOm3tkHuxATPZo69RHmw/TKJ/nG0EdR0SV3QEYYFJLh
cqWT7TpX7Fg80Ydm5EsUYYiyotUN1robG2YZRLKK0fq/z+d2tw64EMS7nkP8tMxM
r2bRjBwdO83kQRhJ/mqqA4lfiQqthzXtBM57pmqKwFKR3Zw94ZdN00sbbX8dAdIa
QppNLhnx5xtDp6iqAwv5pPI4b77Dprr+Dhod6bNYmsPBzgi/dq6XDLZWLtARNOIL
pO0Lm15VnOfTCcQwuDNVqFTucxTvaV7/l6weoUIT2MfcCJU2cxUquCNat8FTBOaU
m53/c+rt4f96sfVzxfySmsyYWskD6l8kWEeVoorNRrB+L0H0+fCkxhfXag3nHNHB
UXoY0RxXFOSbflAYd7HkaPMSnvWIra8pguN/0GOrlSMigLDJX8ublt+IRgDM0uIt
OWOMVNS76PIoIyQoYytFkR3Ybr8BDnR36CarcYWKpbPIU45awZg5eapq/zIpjQ+N
bdeQ2SkEgtlQMjCdXpjTxUsYZjnMq4WvUjKNGF5id1pvijdGX/6p384Ahfae8PdG
vmh+uFvOsDX2IdbQrxQuwb1PrPThAhDrhQLkifCSMl51ldK468uu0sl/JJJCqB88
guaq83lYhBHGYwW92Ip1Mmt5qJC9COhtwB9Fng/spDscghjFXLCeg2kX9vDeqOWV
5jLHnpC0yqoJviovfFuhNvg5qelgiZi7Ed8NT53J7VYCTSNjPYQ1wclzy03aR5dx
xGzE8eIr+RNTdhr4/VIW6yICS3MR4GRIGzX3sXFWvujZcdseonjKkM9iv3BTkntF
qsNnLADCt+AYp012UhnC+W9D5HtHjRMrUm7G3I2XPBdr+GEjy4kWD0RjkAcc+/DP
QQoUzRqw/UND9VCHI15gsiab3JNTSxwKPKoDQDv01wkNIvCbZWjDV2PdVgF/Jv6D
UD+9JQmSZwvVqzvil6CCgV1wQEQy58rIjdP9Zro8ZKQmNx89Xhlxlygay8HfkjWO
/oW8EEOUFtZKWmnZSfoXazyo/H8FM7AFVSl8U39KupGYEwfwYlfNz7aEoGi57Ecx
6mRoCySRtprYkwlCqeV+aQOm8aNWu587aHE1wrNXbXjE8CbMu3F8jchCSMWA5i5p
FsbGFmCGQo9Dno67hhEWZb1ndmXMB1CWxVRwytNEHI+/4TuXS0ZXagSQWUpDbJyv
jdyR++HgPT5gIJ6ZQ5qsAlTJ/OALWF/32e3eiaFvoiW6sHRO6kxmdHE6QBfeVHHv
nZXQMQB6ZmtGtrVXC0CoO+c27ZIZ/wqTilxUdNaUxB7qcMbVKZjUXF2QQ841HPg+
VoYZokRgJluRKKokoCYYAdaIflb9MLlEDsjtudQhjlvjKepa9DlmmbB8i7YP1jHt
QRgsJajjfjzzLHske+q2o/6HfUUgP4PvMttkcPzxGswGNMPIcPk7YmbEzBj6doaG
7JO00St6nyMPF1u/PH18SbyY0IicSP1UoJd2XfUZYMJlfNIp1wwbmDV6BZhbBqGr
cK3QIh2lTF5VFs4bVJvR/AyNfvYnSl/guQUF+3vhV6WWGsmE9EjO5it5lGecaYra
QN3vYtzRJgDNpP9Ok5fexvYcJAJGDLBZyBIRmuQIt7+1Y1hGEaLkiMJEcomnQ7kB
AY1WL9iwjI7pDRgGRU6lrWyUQn6j8/URMZA55WztiuqaeU0/AZAMeXR3NkJzQ2by
dBuMLGEIoFrRJN5G7HS8SFxrHPpTFiCQ866LLzNPLaqZ6tC4cseIlBk0aFEieBoU
HxrFWrLvPSQEmpaAPs2L3UkuUdxX6meV73KU/eWfhIhqyTbm+JQk/edK0px2Yk1m
pbywvKCQS3KjHqFlHqpxkOhhPvND7ObbV64ywXMwh0f64VXbfrFrs9Rhdt9VjI8k
tJNr4DuwIBqzumE2tnlCP/BxJOHICsH6ctVHWBQCOxqoLp0cQeMh1m7umFjtcV0I
vRj6tbAJ+GPPa+im4evu9pmAWO/klJiXNFCKqhtQirOYDa9hfDGrLlBIMQ624NVr
QkAp9W5nov2lzkl7YuqA5sVYBjgWjy+H9Nma7jfnXff+ELYSjQKQ8vdBj8z7iIb+
7FDwp3CE+xI2AW+A4V3Yoc44SGEnMNFjXqN+Zxo41I1IvEbqbLREy+4Avea+v8/M
FPObU+Joj/8NBFreUFMqMABiP9D7PO5F4gHadp51RgLkN9tlxhFqvzKGZpSMUE2d
vgkTBan3VLi9q79YJ1NsuJLnvT4BAq+A71uABT6B0dvAs1YCftYPzOa+tbTYVpe/
Vroa1ryxJt9hDOU7wtXzjadhusapZHjmgUTLvYqAsGeD+3McjyH03Zl9K93q49l6
XLHQGgBQ/ePkuqxqKPzKEOMcyuSYL90Nvd3zKCCsqCb2amiEHplGcIpFTOmgufw7
OfGeIcmKa8aJWR5eKolYIuIcZY/+96PNmsuZdL0NyrpuqlPw4xRqGpazsWh87JNg
LrWABNsnYY7LExVYRrksiFsN0CpFUckEPGhP06e54BftSPy6/TrEbnYe0W725vZg
aPkygY2ZxO2ifrPKW533B9y+i9EeFmeLESC69Sa0a3b+ogxv5/unXNQXi/HeszE9
E2pXIIAyJs/XNhJgGq7zHJ+orCrXkQIHJuwiMEZu9H1aRl6TpMHMu1zCF62cKYvi
+iC1zk5RUN9LhIj92ueradJj6nAMAALVgnWq/uj8i441zBJbju95IH3x5JPHw5Ue
dkRhclIcQzOb6ibIz3/FJndZod81lSBuJU0xCkNFdoBOkkuf4GQBl6a5Me0xVfxM
ZDZDoXCp/snlRtjwejuzuH7th3Us1R/TJV2SoCvax+JMma9M795zLG8myIBw7EQP
KvOXjnNFUm/kY9DZxEtO7cagdwEb8yPA7E/rddpmNCaXxPmMipPY5U6+w9n97q7G
InokkDpdc69pniFPJvwDn0HEKF5bKK0gA0zO3FxdREOnXf0KJfVdTlXbgddVnPny
uxkx+qOlqNqrY/xkSNRzrwXJ1vX2PktINjHqRXf9ZXoUcyDjsfujVNTjLNyBCWvU
9dZi0Bc0J0CebJsHvcam4Z7ia1XVySZboF4v6X1UU/r/hvXiMq+9UQpd9SdGvFMV
LHYNAED5Cw3jM3lnCitlqfb9GTGCARusF4WMb4uNRUqvNiwOo+Uo7SKthOkObMLc
pRSw3vg+STFsIpUdHhHp1oVkhBC9aqm5J1NFnXs8B7+ewnNfTpTiPjf8GqMzIxGT
gIrEJyv4kyr3DaoVdopmBlImfrn0sOOwhsmXfi0UjfE6ve5lc2yIqqoVEPUKrNF8
7H9KthgseJx0WdlIe1gb+KbigT8eDiw/7Ri8Na/JceEdkxSlSBrVJ7T2oGgU12J5
sk+GT80yY3EWaOzTtW+M8ktJpXonzVUf5m+TWiTmqwcB8ZUy6CSlWtMi0bgpiUPq
k8pnCkL9pdEiXPmfHjh7rs7NzzU0rgX+JccOCAn2pBmUsAd9dP1b7tyaiCNAr9Bs
6Z/DnB6qtgB4TEKlMTdf8Y6QbAMmmpMaOpx8h+l/8zJkKWxFr/S92hgv/8wgmJkh
/hBbYRTnnAvIyWO7Tr9vI7ikbt22U/nMM1maulpors0CcdKmXccYjCDJ1LJJ8/Li
0mLCI4p6DKkeTjNlSax/ly432pRQpfsG6G1OkhLd6LEcTwi16DqTw3qrLhTtu9gU
0ydiQvjPHCxcnldoSU8hWbeD6TVKWcw3Y006rHbSOLRDqCMRrXo9uJyaYqZDORWv
/f4ZmOs0uHnK2kAgVgw5jxd1pkAcgrRa7GdgsU1qYSmuUOlV7jzc48SLeMzxiohV
HriV7JfXlGbz3Wa8+PJKF2xlnvLsE7BmXgexGZvbM2uguyT4gGx+n4KgwdHtkJAb
M9/Fszbdn5O/IpTpWgAINY/KufeT5VG7YFnAr/3OeYE4WASJlPmTGox7e9XKF3Rf
g4YKjZ5MYGWDSlPSt6aBEExyjumLkKjXLOCCnoCYWPZVacrzoivB5LAx+gW3vwD4
/KBQnuJm444v7pUTMuMiQ1YG4Y2CuuLA7hrF6N5swMQ1X3mb5PXv5j8A01TtLGtc
2qWnUT13Yl/aqqliez15rLtJc5CQNCB7fajBOFYopBVLtubBqWgfXMPOj7NlCoGo
csVaXiJgAmX/YLiWS9t8uLZo6G8Lc89YOIi7SoYIiWemH7uhzbnqTJdAbxqhZNVS
JXZ0RUX1wgeA9I5kOJUrL6oMoJW8byz79QYqL9Lb0IAwVDyP9FjL5HmtyPipNhOx
nB8z3k6y8GmOpcesZ7Az/74qZEsTxaARW1NE6kz45V8BwZ5RdXFnqdDtS/Aa2xfJ
6OMbRtt3vG2siWaKtqG/1xDhP2ik2kv+9Z9dVArnIJDpXKH/zJGs2vyCnZuR3IdG
RK1fKIihECXSB68qadyyzZ2MAt3bFxxZW3QJ9PjipY0hJ8Hlab8wp4TzMRUHfd3g
xxyOT0Mo9f9aPQTFfkL/yFSnyzj64LoaQHe0P+olDJ2veA7HF35nJea8dPvN7Qr7
W/wKs6RqyiFgIfV2xoQtZfz5ER3QB4byojXgWMk70CwN6uuoePNARFx5rhTM7nuI
tNr3vNw33qjNrBLYFCHIz3I8LvERh2PrG0FX8Feh5+YoFPNF20TKWay7d6FGi54Q
n4ZzW/U8dQDpeLi7HrAlFPMf8sOdvzJKoQ7ua6QKj/plEzemSGtI6jWA8hvuDzAG
d2wHxMBWN7kPZFB5nIRyjOvjBXtqcoblSmjdT6hFXX+Ga8ET0vdsvn2J5pB8znx8
MRfWa1XeudUfpm0b5s/K3Y2zoyXog72qVpPJNxhNAVh0s360X+6XU0/d3UkBcTp0
wjhItLBEjcjO3MBNK0kxvduFiuGpGKrp/JkwkRSL+Cqsna4+2+0jPkGXKZglWHX+
okusmXKBHzIu0bKFCA8e3sjsrGl4CiBnqPppEeNQC8zLOvx4+D+5xetII2URq1ui
WoSy11P38Lr6u51gIX7rMEeOtYX+UDpf9HNmIMY9UgOtFGrrSlLcW22ztNlVmnsF
3V5t0f1WTueK7aPtUqdGnOqvzs0czhJNv6gLC2j0v9XduYWQQoyfkegr3zlFy+dZ
KqX9JedtyA7qTr0MztXXA49xkj9CnJRYEMSgInwbwh9Ixl8C8cV9Ap3s8I7GuWnN
UA7vkZqjLzx1/pBwKPoJPeRRBzpICNaMvEngcSZ/yIlaI5sr9EptbpCGl3E8a4uA
jdWT1SRDke8lxguvK8DM0u4ik0DmSax6Rxjz3f8S6EJEczhJNG8Dd+Fyha9RFsko
LEVBHKZVsOcZaGgvyR0oipE35Re3AaKLvKkLWA4JTBCZv62AcNfpp3Fav67y+lzS
KtVROo/b4OilsPit5ECv5fgZiySH15BMhcTKeBi2pVqTtZu95pMo1Ry8BKXzqLcI
xhLamY4nl/qSrRUJ34BfsnmoPo79iJqkTIHL5CWvZQQ4xJP5n9DROL1wFFL5pd/g
tvePFPG7+aLxsUHfQ6y1D8KyDjyTbd6cppi6nmcBKCuJi6R4hgby1vB15SPw4a4e
QmvYI8C/gskS4X6unyHFHgOBxWZUQelEyx1b1gBpsgychWXTXYWH52+WBaUNdZTS
CGH9wMnvRRH7UXuix56rvqeCv7pJfwTbMbryy1TK5VahMCpQDJloS+Yl+L3kYKHh
0t1q/ScNBseYqfI79EIAyYaQdYwFVKZ5xw2xbifZD3i0h5zTB1dv0RmDo0+mX86c
PQyWSv0gZz/+0nNwjr94aGMJZD/IiVSG/xm+e2H9BoNomAYYB2z+MG47x1Q/rWoS
uQ3WNhlvjlQv1Yx3FCkfJkXmsTXeGh2k+dhQ/aaDrOzW2qXSh+8oFsXCciCtIeem
NUR1iF1oGqeoQ7ZfcGcgEgXEerkdtotJ+Rzn8o8f3kjnm3/qWw1FHFYTXMOKNSth
m8mjtOTZXYukPgUJPQDlHNPtPII9WnBa8NpeKCIsokp6RBen5nu0Uwb95/OGqINS
UMpCIK3GK2b1T/ytlxSG5jzc/hzxI3ESsdDZ1QcknAtmC1bYNZWxjSpFoBlaGHhR
B/sL6c+PHYJlPxJNubIzm3n0/U1kTNjURg7zvJWixI31YkjCxQuahOTkqCbvpWsc
DrA4Wx6sNvOnymhmMDj5/6bL7F0y/l87UyuYTvAythqrQmOPosXOdjF2rQQ5sjl7
IU7bGxWjg+caROS4XkmMWS4a1OLbn4hoIbfOvfS0q8+RglxB8dW9JRvrty7F0FTI
Ru0J2FI6sp2dHX+R6LglITc/n8VtpSI6I4MfiHLlQovp5F6fKDprYEa21mswca/x
ap0UEcVL45txOwfRgiTKuLG/H8tLUX976Rb6b1bM8ChjNIRi4k/pioDlGtLOdEg/
kwv0svdoYguc5Koxpav4/xjnIvWoeGyVhaaNuq1qvZqsGnhkS0IejYGNvNo3BC/c
xM7aTlsJPQurVYD2s8qZE7DmLM2iau4UdeqQIqtyZsb8TeBJu/EMA7sT7sMled9Q
Z8oj4zRsc7feEj3xpY14Uj0Z6s7dR1clrwyJZ0d+K9DdxYNlzoUsBif2sCCxei8w
EAVBDU0OjtsmYqw9arbI7cKw5pOR7vxFYl23Spq82Gb+DBhiBTjzgVidbcfxhOSo
QoRV93RocftDU3KFK7Kf4a7xX80B0E+QN6QB6Mm3DBfSLd4Oz/nzHM49PJAIxd+T
lLq6jpKF7rC6s/rhN03a+05P2dKXbplrXP2wy2mS4tIUsgqKlP22eKgH/dqsj8Gp
H8xu7BiAPJ/zT3XEFfH2uVQLgegokR+VVoKWOmq2WgoOLMLI5WC57Iwz7nEeujd8
2SvvsrXoZUjXHaS/GZUuu1OcOB9u8YjkovPS2SNv3qidWK+4UORHJg+XxlPFTtUd
xGKx1k7Cd3EDz8yEDDTtbxvDrcATqt5cHmTXEQQpwdFUTLTnwrkwdS34ortf8adJ
YYKQVF82/tGKje5SA96nTa/sTdxk075aEEn/OwVf3mLZ5y26jnBI76KPBzGUbe6I
/OdmXY9c6g7pc9c8PSRvmw4/d3Yczpc62YVyN7Y+DqeJt3DTrv4kb/mY1dt6SM7o
iaDcenjtM3mCfDFD5jsnuBFgdiC57GVb8iJ9+9KdkFzMFZM4C15Z16XTsfulFUoY
ZeyGzPXeaaW3/JImuJxxjN+i29k1CgX0MjOFifIFOJgwWQiUasVFw7BQefD589f1
JotybXz3sK68K4+Qbd/eYG2A4ClTprgvtvAYGz0+5Qs5oXB7/rvzTKDF/VVOBkhI
iXZ7cS2BqVTjbSQT205s+K0wlVk00oGu75fgt2rLXm/y6V3Bhd4zKVWmxmUFw/ok
yzwgw2/YbBHVS5gyA7Yon+oMnEPzjGlN6GXAfMOBur9UixPhDDnMMSyxy4Qxl00v
TcOozmDT4qvArny8OtTkP2dlZPrFlgKmYunIe66d51S2NGhW3kS0ia8vUtpNC1cA
P4XMZm1vwc1d5np+ZNPR5SsBXbrhopoqXh44Jz0iw6T8uX5qBlX7dd9W0FRxgDL1
XLGuA0VXmBXnzUCiMedpRFPPHKudEUS+yaDAgJaYqqD9kSr97sW9LlAY9YpDanhc
Wy/hisB1m0en5Pm4o8oFypZx5bpH0gxJdZpyBVs336z3xWZpaj75B9Y/SAKqKFXX
qXhT3AtObU0duqEziWZ2ln7vATmZsZ0bMdDSJWx63HMod+Gi3DukcWxmuU8VPHR7
CVO7pBO9XVgmBuf0k06VgO5k4NjWFJ/RJHuLavW0nE+WHmflZvtVw627WOHt8SZN
xtS29rQp4AXfYETWa4cK9f+dOpa6JCL/V5uHkmJ7DOev9wskKl/k+9wUYbaGFt13
iNTaJbEBaHnaBBih5ooPURUpRZNYzuNu0kSbTQMNdHb342yVWWzlkvTgajkv1v10
XKc9ZuoaIzS4VhWdbdl4f4Sg089J0+1aIdPJ7M0+cyRb+194gnr6iun0aCXF3C6z
wGVPuGVLjAwOhbJybZDmPfdHA/XWt2C2C0bd7S9FVeVBBdr6afiru62LruDjvvCQ
G/6Khw/BqGlGfPNWqGDhJWZ6ccSrx0kuWi0QT4lSgmrFqISiiLDSdwGTjSUicBj9
Ih8l1Ls6V5hZ0ujgF90aWvuOdn+IzWyqyE+xR4bEV+Xyyil/D2Bd9iY+msxoVZBy
NdLzMZApKypSYKSmWZ9FpndXIjYfJ+4Q586nchbrqrr6xeXQr2zPN2w5J7X8HOMc
IuJpt2jiXia/gUDS8vj1vIL6/9aLDczNc2DinoOvYnsS2JyAXhGYF77t+LeJt0FM
ZqCC6T0QqLPg7mQ259Otx/0SlCqXm5lpDQPG2jMB9AB/+4+TXHD1v3fuiaFjKW2t
PPadmNl3rxFU+VM39waCGp/EYyQB7LL6sfmHCgMN04fBlzMjoQcSUTq5iDDjyfiv
ttrSiio18TiI7rKeY/U/RTsr50AjfoX0Cg+xN9obfWHqTz5BwC1eZD6NZIvqIN/s
h8pq1CnrhhAFYxyQtMI4l24i/NRYV+/DUZeBzw/3EYSeI2lfiTKeNuoPaOqVYROe
sH2wL2t+Hp/PkACAGoZ4lQxlYzSwgeUdpP4QpCXTZMHCxa60yHba1tMLFX4LP4n5
NCtNBJa9UhsRW1TEvD7QhH9bhu4dRIR634K5Uv3RgF8UwbpAG0jooMkd7rJkbYwY
dv7MSgpQLrB1+3lYIE1jbAt/55f6GHHetL7UWQwrNd213ANHMzveGih1cUdl93a7
i777qwI8hvso0blWOL9XBMGojxuIyHb8d1mt8rxSHN2uzb+fRUBBkEr6a2AU/UU1
K9l/n6YK9MdZ7blvkkl5n/RNjHLvsqOhMTibx+tf7bsEe8kmvSzIdEQVjnGzDlFS
nm9G0GPgs8+otebUNtxq3IIxhxcpekSpghCL2R3huv335vOKkPVuFDoWn6xll+JQ
NJziQbz6owpltTWO+0q5IFYNxOMJzn1DIqHKAaAc5eY09ZJJZgNjzCMhTFoyp7qG
yCnzg25s29cbn2kkj/cntfv4KNV0K9dNBFcvcAajXH6nOzXIgFEJJG2dJuGcSTl0
oU3KXW03BNQ9G+jdbNq4tVMDkydW58CwEaaZCjIxlhJENoKJrQ4u0/GLOz/gixua
Vr6ikNJxlu0Zox4YKOMVxsKKZL/sEpJEfFdx/NAlMijqT0I0O6yNmMmm7xB6JHbD
CgAwjI7MqvGxZ/XhZDLX/q8IkxauDi89vJmFwNu1W5JZbLUfV7JRE2kFHxhZb6WH
QXMVyon/Dakm+tgfCRaCCN65K5zl12wxkLQjhueg+e00zcrPJeae3Yf8nAj+jt8+
aW48/sp/kd+AOtHoQprneq7DI+EoD59Q3QICPRoejmY2OwsYGQeCZubl4NWS5Ejo
hFPotaFdXMHhyZqEbPUDfblumhUuFa4o7ALGLRmN48ilVzjM8IUKyWYbCvL+99Pb
jID8A2vjngyfh+7klHpxnWBz0gRZ73s92CSFwz4oB4Yti3iILaK3wzhK3G9gHt6K
Yjzm5V6q9hFEiS0VCrKaGuv8yu5TdYjPuy/nP9DhYrZSsScjMrHANc6QwmpuxA4G
ryxkc2JXpoeffRcKlaNIe3AiFxP33I3a0Nz36sVJB/lOIu3RndFtkFfwAK2y8I8H
Zp4tpKoGidkEyfD364rh5V+vaXLFhI2yxUb6fBZELDXh3zpB2pj4RtO0o/3DpHRD
Cou9l4WjafFOLj8Fs06+PcDgPPtudk42oe6FmJO3pzwvhKRB6Y/6BCc3Vw1lQpWd
5D7LlJHulFnk3AvY18pMLJ1OPrsdG26VtPtPlkpF5plgr7juQiTCE5/7lLxvoGcN
HxypnxCJ/B9NojoUHzWhmnEpUsi+7qyibrKVQcq/n01Xxgt/UfRU/DkWG8iW6r7a
j6HLjRhj7teAlGPAuhLFYfwj8gRCI/ZYKdr3VuxnLwTXG9rX1RlJy0zRA86MmBMy
qXKD69HBxIepDDdVgD3K/b5Lq+5tBk5V4Sj0K6CDTtVqJoBR56nFMjstN+uaXRTz
wCaRr5v2ZCq4gPJFvtmFENJsQWikgqkTW82ytKROpUu2uZj3Hi74L6qW4uok2hRX
MNKLRy5kLCww97txNdAzrL0jEOqL6o5+SxOwrYCB4pBOYHYAZZUqZhNMkehjefiy
iJv6XaWziAKn4o9XKf9atw9Guizc4RDAQxHKPwNl7AeiHzaLh4njjFWtUAWl+bDc
W3BVIVf3eauMOCuqwicaBSpvTvFuxTNar+p+utBWhm3PmPepIZjdWS8znv5SxeiQ
v9Fw5bV+4ywWF4/robQvFbFY6OQiolRNmQr8NAdxXCuVmuFHm+LieI56DhYXO7jI
O13tmorVBp0p8ApG5Naehgnxy8G370KD3PAyTT81ZViU1MoMucGz197HZp0A1dv4
wx/8mJtMCMM3L3E+LEFM8gKZBARNqW4wHsmAiaHNpsp1usxFUjprLlth/9Z68rRk
jKxTG5UUbPqFxbKQweyQFiGPD++2MAOOrA7ss9r1u4V/qcyLBzOn187WQ6e705NC
y2RM2kxyCImG0dzZ2JQzDVzH6PQBW3WbxF8yiG1nD5OKOjS5C9c7YnK6oz6os5Gi
UdXZzuiCDhYtq+1cB1zFeI3GoxpQLj1H3vSabpfGux1MJdnJqiZnQ5m6WJWRRt5q
B4pyYG1VoWI/YTyTcRM/ud1we1Nk3qfm16PDguapmValEeE/8uhVK8dp6dxdhWR3
yRpM/lnyRUT4t5ZI0m9Dv9fAB3IASnYlNSqKtUXickaDW+ttMRAsVKegtlwIkdEE
HTWxfKkoOfynP+ehfOUVnEo/nRs3cTMB1du5GT7ufeU4VKZAeQ+sI1F6hSgZEhf3
sEeelpfRtvJY/IXGWEmIcOsCw1SpAOCYl0z/yEJFhGa1UQ31xUWb7ZHYC1qRadD7
9eCBfGIvRb09xp5JnW4XvkDgTy4vUhusgdiPqvUGYhEJzq0lv1ypr5634TV5Go0w
sL4ATaWw0/zjWFTcue3eGVcam7vbAJjvpBVw2Eh2CVDOSKHbqVbm4+Rmlr2fYi8C
Gou75zr1++yenfhHC2/IFjJqnOJy9Qq8bu/rDlpcXFPiimc/iobKmWhwoqPPF755
y5tL4GMy/NCeenKfuLUwR0ryuljjfX5YhwTGlsTjMdj2FJi8e/f5bH6YrpntOs+P
tte5fZcqmU2AWUdBAU2ihVSFkIG9IE/uh18T3sqkvtfWua4BHo6pB/bk37YXCxZT
EjcqSigMUZl0BAgE5ftmma49qs+nv7KEJj9YvOKCouXan+4MqpIOuQLHEsHe+UrQ
KgLbD3eudxqEsFTFMxPc6M2+/42c8HmPggbyAPG1LIznGo7KEFBcV8Kn9+8jo9H+
+962i0m5jygmGbkf8hR1BCZ3CGix0bWffgMRe9dZuPy7wW7HXGWnpp8Sj6/lDUyI
o1fOCBJyBNFPuTA9uKVo19bRO46kCsJ/uH5+8G3pEcdqh4YeRkF4qjtBysc6E5aW
7/HmNIV9NLxfGds8MVfD6zbQk+zPuocipz6VI6Ehmbw09TsVkWdGyP+MepM3tbs9
20Et9GZErho0uJ0fDJ+93A2IGSF93Jbs4WB8I4PNSYzoVY9nNJQvtwuVm6OqlUNh
7vBffvTQlA5MVEqJvs2L030S2AtXx9nBxP4OcGfQtcIvi2RIo+3K9gz3RJ/G0HG+
d2TEw58ug8XY6ilrACo3NS3T+oE5ZLkeJWyAP/mWZAFoCSk0zcjPWEWDZ5M9VUqZ
GOZF5uVsgppeDTX9nmTm7azNJYHWyX05+eF4kWwwt2YwPdj3dzUuriSjraJXwUL4
/BuGXZ6pvzd/VEpMFN8p2XfmLbqWH/Q5duZDD9RSNMRBTwX9zBzIsNbdoia7jZAg
vox/fiO/McH2LrFVXF9irSv6Kd26Zf4qxpwmMI+qeJykH3jbhEJk6Z7ssI1/oG5b
uCTq0m3sQMJpbGSuPIhHfidiNJXtndU/7wPqvdeaDtRekJ4q6rPjPrfijGshVduc
MJ9rhxJcRHTLqwgTSZub4PReEfg4C8HcZtLSF91HDTRUWk00/mO7/ZPDY601wlnc
NPFoU/KWwv5/cz1kX4yo3FV/wU4aIJqk+8IPGIsz3Mf7fKFxUuzcrGCnpu47h2l/
8etNdVzv82HJo6Jx9dhcXMXeGDW9n0BRivfEyCCXm7j++crB03mmYLK6j2l58NiN
PJNValHSGEZ51frDlNZwXX+1RVI6vTes6kXNrGEl0mBLaJ9UnlqEa/xz2Hjq2Y82
vTGh8uLp67D63kUp+9RU0WpHx2Rj22HSe1GThz7CisUGzVGt+ClOODlcbU0eNvcG
/bx69zpca6pQ0WWgZ7gWJfl0IgfScePwHkELVvBc3FMc+mIulz+iJQE/xqHLQ+Fw
p5nlmNhOeXyQv3OjA+9DER95VKSvaEv3out78sJbUaqaR58CauBftl54JvOsWF2J
JDUZ9sgWNj1Tvvrbc52QY9GEBqB8BcccCKUKC2FIC5nU0BGCFYc8TGRVgMHe4pM8
J1KgmXWr9CJKi7AFZPhyclXvUoDT6EGT0/hPL8NSCE0aDe4K9nHdV426FkbpK3W9
o1Xb4Bp7qbkuq2b9Nbzf0kPz5150OYVIjvy2hYUDDDoJj9W8u1VjOhhur9th28HO
OJGbsaTRvL/+9NciLjjhcLSuIivsOCivaxOas+j9d0eyA8XKPULOMwsTQmziWCIO
SG54zmA1Sx59hZMH6ILI/ql2ikzFCnhaGWOlzbrvGqOpql0dkd2ZjkzI39HhjZWF
DxIHGrArXfeW0R+BcqO0vlJYVV6ACLqvGU9KmVKSgp5uv+AkfKgKGCXBNV+qXQYq
7qh/nCVtnz5IAOHIV1MG3LdmZxPgiMY/aN3AJpCKENkaT5NLLfsAuJoE49kcD43Z
EaR0RWUS5GHp2+URe0F4K53g9wi4T2J8tJ8qlMZqa10NaTjc9j+YwifmimF7gIEx
MAxn64LqR5kbBLsQ6OP2HtG5sT2zHn561PU4q/jy1Wv9xzVvehfSWnZ25lAjyQef
O2J8WDmLaZp3eTYdatLOvPVDxRDc9Wq+ZltkfWd96Rb5a4d27Os0BBjizW6HxmQ0
Xo7q/qykYzSlkoEPNt4r0qSCxciHhXAWRjG/5tnsWlXyXjxyC7emsrtNskFrLOzz
H7ZT//PMbtDBQKhyaEUTYTLj8Dkqz9wDUgZEpf/tXSrLUI7Jg6z115oc478vZTcf
VTiBWD4PMgAsin5oroe/QyDQC76q6GXCUV0olNvW14iFRl4RBcW/STvBaosjuW/F
c/Oipmq4m+fe49iydCW0Mvc2BzCHyukvGOI1sJDdgB1VLIF6J+ffde64GX5LHssQ
pCD7P4inpeiu5dTl+BuD9PgQbsdDw5zCiatFyPYChYn7bYF6tUI3snAMcdeDFWW/
RvP5HLWXHk8gF/AP1BPn+qVZPi6hkAHW1N+iLxa0sclksthTdSn9mjADFD18J3mG
sUDzML2EkSFe0cZRhGCmOMo1rK/z7t7g6Wacy0PPdrd+aOz2NPFyvFuyUP9E3FLs
Sy0BUXf5XXuykL2XC5+ZPTlEdX0pRfE93h2Xd8TYBagrIaxoclTE43IaACCElwCb
s94zMBrZedP9dQOpKnrQRe5E67807779PA/614Pqm9epNbAgNgkdk7pZpCJAWbXP
1dGpBBl0t7AA7MUL5D8LeWHyX8IwOVU2XINzaBjErL4YYifKF1G0M98PWhvG+RgH
KEAM9BRsDToNNpCDOuX2A2Lq+9iM5Zqqk9zDqWCfJJq4YV5+YU0Z2+P/p9EYgZod
x04iz3ix7B7ZPTfPud+4S9jMR+qizvjJ18JkesCz7+/M0uoQgDr+OqqIL3Rmf9h4
DRE+eT1RKAtWBa7hsIr7DbhrifVeiwyHEQRYUutgpjoze9+HvOyeFSWUJquMdag8
/QAF8iqguozmz2M3B1zDCRhslONze6jlUpYF2qVqXu+Wzf09VzmeonCWIVpfkF+b
Lr69e50DoWafzTXujZy3PBMfnyLsngNak/L2/J/3Ya5QYZ/0AAFvDkeIrDNquNVV
eUayHEUE48yqEv9nzRppmh30bGGx+e1Z8/DSJdkCi5Vz0YfOhW0DaevbG5bUYmwv
els5lZbmGJZWHsYsUGjlwUC8j1HD3axViwMOo5xxCZIlUYz9V5AKPE0u1WYWKiaj
tND4i5cYNQEi5JAchfsMCfekFJ+MP/TVsp4OBaXhoHN6DmcDnIvLS1R5rFJTQmI7
u3qSVNWXY4ja7O2xV+D0jPGL9hmQWofzkPK9CYqKG27DSZvVsCHjOHkFcnmzXZtI
YSAYK6XZB3M3hZjeSWobsPyO7CtfJ+3ySBTDmofOh8bUwyvDb7wbv2MEh9pgGrG8
ZhGERFWZrq/xzWlXP24RHeOLrGiYunmjXqT0m90McIbvFSIyx1YvPqFhGO28i03H
4vxypeHmN4fUsPoMAeIjkAgyHh7RdRQeQg5yrEVK4LLbBrc/klY76xMmt4nKbsi9
firEncVoNywkbv9PUmRJfcrexPRzphzs0DuJiE0OEz98xDGSAB9TKp8PyLfQ4tQ4
Popwffwm22uF5tQGoyEZ3z2ztaAK1vR54EwF1g2tmU/1YFKvAuhpPcdqDdfQXEGT
VnzEPexaK8p5+a1VpaiUJ6o2uqXBpugk+Ac27Olj1E6kQAvnqyS0wmnyTTVYAgSi
shbYbnU7V2HZ3+AFHDoSShYBrd5zI/GxTaGq1SiNiPhf5BBrhUpL50FYp4+aIZiv
hXN+7LQTZ4ik23dSadLXQDdkZifsJwJIJiaQz/VPAanAM+GsaPfh4G143FnmmZIK
MBBRpZNrrOjY+fiq2NJcz3Xx3VDjxRaeUNFjuwDgQu8qVJogWHZl5ZI1hRyvk25N
3hPEnsiEcpG8wiWrklv+v/C4ULNgYAHhTnKdRp8OxN1TmuCWGjmsjUWFF4juO62z
3F5IWOYBinpOg2W+75yPQH56qKW4r9zyObW3AaVfQ288hqZIWIj1bxGYLDUdzfQZ
/p9KwlXbZ54CrwzzyB0Ie7BcZujqmoGN3D+r76fz0ljfjLAtJ2q+9S8Kp2nzBBgq
tM1y4SW7XwacQTyHN/ayo9rk+n3sxZbpfrRUM9FDCer1jThOq1CZseLur876lobI
nPYFct+F0wFY3pFGl240kLVoVRliKV7EVkkSaUml7RcN0LWBoBKbYYHX0ofkrdKm
OdgDKyf2CZHA3cFP8q6eSPt2kKxganG8w2PasmpcE9NncccPrPPkdIDlZf6RDIpC
QZ8OA/g93VXzb+O0g7t1LAXpE/iFeE0lIheELTB/6T0uIVW9wKiEQRXwQG5gufZl
TJzwLrDPZVJi9VPDb2oWt584hnpfljs9OE80xBkM2xlkKHZB1vpc4J6eZwrppdWo
/bh9ssYjVGtESXDYqUxT0pFkd+TwlU3Li/JBJgJzcim6jaZl+yuI+ZUIzUkPrw6l
omuqLShNWNwLPSYCOJ4+zXTazYUSuhbKaEhJRxjqQxsNzncamyLUjowNpxXRBL6o
DND2LYcYLsaxbL607bA14CRgBMBSQOlh+2HRyLLaMMoAwMsBhOJOICw5tUVVfFjE
7KB5vOXGX6EhZThObgclJ44YfvKhyWo75YzpdeKoyqqZty/yqDsNHWg8EGpuQFhM
IXb/L01ybIpTv3vy+a/wayuWaznFb1rzlQyDkA4y1BovvQn8rJCRSNtzqw50ZZ8X
8H9VbBpFbxubgi9gYUKGP45dzYahF8cb4DhObHWAAa4zQ74ygzfQ20NQy6t8Vd/A
OzMUKHBUbYBAQjb+x8Ix39YzcRUiudeDHdTqlcJsuJOH00ivufSqi3KXG6KbDuul
owWVvqzR8xWr9DaF5GYGy9y7xeoN+Lsjww5532Va8yHfsLSnnLsNMKcQuwYqXyH5
O61aDwFksATzWXoEnlGfu4OvGI7acfR2tW0DChCStrNbmDChucAGlZp0az8jMDuk
5Y2m8N8KgcYqc7A1ccwkbv/ZOWyf+t/uN2YYZ4kKNVSJfs68ne2PiWdpx1puwoWi
KORQCEYlJ+olbmOw0X7hPKAHiYc+N6xFZz3lWr4G/KE9QZh9NqL3eoOztqVTb0BU
COoJSzNiLC07LAYUhN6/c4yCZk1l2Cr6pxbhOCUK3eaBeUrjYneiogVYgpL1W9Qo
SvZLqWO3k+TvvFYkCJhwTFezxJfen6TERSerlNKeNqyx85AT5SlXjyE3waa61Bpy
31vGvJ6EwZwVHUeYDgSuHd9yTk3Z/44AMWYQ/5wN+kekBRKxVFUT1vYVjPzHiImF
ZeLA0uRalo0lMrWd/KMn2USmb+pRq4NhJWjuoCtmi+FJFodmtyFNX3+V+9bqj38B
Dt8NjXTyGd2UMjOWoxzwWcfm14Vdl14QrAXRKqgUnY8YhXjEZ4Q9OqjGDZOAK1Bt
kzPyAQSDVQi1BqU9w8PM6DNZ+Whq7uvzlOoq102Lc1av6CRSuPmZ1zYtj6b7f1nD
ctCyoQV5IO6+1aPpkMVB5UCeilyrgKTvmApotlOpI0SVh2nm0xFhJq580q4LAuiN
HCZZjkuIrW1YtHRXmdiwwOnVUpMO/H3Vy/8dLG7VWalxp+ls68PyDcUTXJ5ZJV+j
9T1Rl6xD5cW9G99gEblwgIELvnz2RyHrjRjGW/9datj9t7H6W7f+O7g+pt/z7AAi
tAOW02uaWfkEIVEc+B+mc2zs4FXDrJJPHIdhmJAznKLxoC4l/vOOQgDCTJDKbQ+0
EM9k5Fg1pGgThqfUsCuQTWaBcLYTBWOpyNrO1fhh65JeDXlhHwQV3Jn2MUOlqM8w
0ICwnmvFDgpZ6As45xoKVu3enMI63wN33MizhKfeKW7bW7+t+lEUAkxc2+yYzYcx
ZzM8e1V4/Dsy04J3n/lR1GLNMS6orDARpIQuARWlulZcINjaEoGSOy1uTQcs/k9e
zrrXmg/PIrZ5v/21VAhNh1A7ochVhEXRVmovZmX2/P6Z7uN2YYHKeVTzNXewU/Fe
ZT7Pc+BfMMzajp7ZVgq29CuwYdK6lcl7CtESvWqoSdPNnjcntjZWxR2clhiKU1Mg
YF+AM3NH578k+trckpTgM7BE/UBPFGEMApaOwlN0ph6omfTE6sT1LxCyEV6tEeoa
trEQybs3/xZFzA6bHZT7pvcuX+yWTi4s2yXbd+tkyIjNlkoWGAoJaRxGv+9PdZ90
wH3exgfBUcWgM+TACDVvR1xbAFsq+SI+EK5iJ3pWQGeVfApKg38JXZaUq1JqM2K1
RxWT6EX3RHQPrgerL1we4A2xhr/iFTyUlp0I49hpqp6LCWrB7UYKZaOh45KMFWfC
/Nu4sXglLQXBDX/YWlxENgByxGJS7ICK+EJ9/arRW1EFyYbRLYwOmf6q3I0TqkBh
Ei8XabY9WAhN9X4mIxSjInNrpbGPidoDztKEXI5eLImJhRA7MRUFnVMFjy5rRtDm
R40IUCEb5XZWSOezCRui7ACONqPTr4ZkCGwTza5F0bUa5vatc1ePOQSO7krvJ+/j
z5GfZaixGgNM8mLn8YVzaHlq8u/lzFnJmNSY73nABpQ+rolN8ZCkXCv+BDKbylai
KWAcUOytILy4WSUzZaW1ShplOKN4XozNZG3KHj3RcZRAhAf6IcjYgl4f+bWuh117
GII0XUkOHKIY7i/HGQtwVUFWloBYg/EoXiOVqCVE7lo5YihYzYxL6W/uchxyNnfw
buPaaC02sXxTi+uWYX6zd8WnBQd90ERbAaxNLlqHH7NWQDwW2+iSyq7vDYPNRnHV
F74mj0qSNVYg1KPzEBR7alA+P+xPHbWeG6lYsMn24e2AYXu1BTg6amUVO2YeqBEk
f08zWs8gsUogdbIc3Yj5dkz2CJKq7pVLf6LJZwnL2bR6Kx7na2Hq4fE7MbjYreD2
1he5Jf8E87Yrrlvkf0meL/QX+YqyBk0YQ6F+kdPhalBpk1RhTqTcUbsrN9uzGxuX
zQkphoZRY235T8CBqhEt2rvctOD8MRoJcs88lVdNkUn8xm46jK9B2TrTR4az1Vrv
wOvhWGqRVYpgsJ6z51oMHjC1LEaHbCVyK5Bk1yOVNj1h/NzaDDKZEUKpXJKOE3Nf
R9ygHypEQc1RdzIG3/X8Gp1Eotm7nygG5jcwqzkiiGfmh133j5clZMc1KizCcLHW
On95p1ou8KZ1CHoVK0HIvfkezNqFB1x1SXYq0mP/ZjpFrjz1aTevHL0cqLDIfPKs
Dcr+z9SvZ2rPeet4WKgfeh+Bin73ervUTJGRPOT3M/ettD2T6szbLfj+yDN0urVM
/OwML7tiTD3TlRzqOh393S102hIDSjALkkCFrgTLhd2tJsP+rBpyTSp85BZIBgjJ
rxQNnoJGXlhsXok2kyK9p6oyT8SDHb7YvA7lZqrneY8Xvozxs/FqdX1P3rRneb82
VZPhAtKwKskCiyCcMtoBRh4vP6uiC7myzh/pYTR9ZeDI4VyBJeVoJ9yjTmpaD5kA
DN7BPs7v5HwFqO0yz3fejY/fmTflWcgY7jjkT6E/6geNbIzcgkRHtDCtE3CIw7cH
2i8XDAX9BU745xHaY19e0CmXXbf4kXpUKWF6wBBxrj/Mg2vNy2iAkve5dJ8iG+lX
eEmuWXPKgYkGGvrHI/NnDMM9g1IQCi99wlO4MmPTU2LJMo0NMiIK1T0/PZJr/v4G
4mW33ZsbA5TsSTtMyjhnuU+oLq00Y3IgrqkZo2VgQwZxFB9DdHuvLuwYrLzM2wNj
6K0oGzAhkSd37DMv/1TPGSNrkUI/9/D0Ndz1xWR9OT1uGife2WZkx3Nc4UI2PO51
s46WyTaOkCc+Gh0c0+h092S2ZwYoL5sOWvLbZ3dQvu8Cy73sFe0oExjiWKsrPwIP
29UFqjo0GYP5BaNxodhj7dkAi4pd8A1rRHnnDKcedpVVc3Njcd3NTepkgqnKtrD4
At9fT1MMaI1Kb5f4HqP9ddLRW0Zln5hNp8T3GJoWb88qdD5vVlv8KhiRmSI6Kyqu
ewn8DcwL05wu03rw8aEnNLUV+M/OozXOaSo1rgMdYmFljOu2wBtbwl2kWTdSGAqr
qA1ZV1zRzzEpds4x+rtpqhgqoAam7Z5RyKhoThHuXT7tiPF+ebWNZ4iVlYoz0PvG
n205NYH1FkO3hg5yqbY6+Xmi/GvVsZmWfZQuFRFWvPBop0Brpg6qagX+1WVKpr2l
oo4lCeos74U6QHj/HQlwXxhralVDYeqQLc4uGgzxuzFVG1T6h/cdsBfmef4i5MZX
DHadBIjCUFBbkXEl+LZz/aiFqLQABbkaB7smapU5uw8eCju+L6IxaFj1rcfFwVAo
8bOpRHKpEeYvryHhQN4YJjucHa8P/+skCYB1q/Wzhl8ztc5r678KVuhws+o7k1tc
8rP6bf9KpULp3ZNW0iqb+inl3nOm9DqMAQVxOw2Da3sK4U5PRyTGLps4N0KcBtWH
QiTFIgeBLYF6nFAqLAuETxxrh8ePvj40dvIRtXGnsqM44r+DqPKqj3s+Jktm1UKK
BfKlZZba41WkeB56NT94icJIpq1DZmTwBztKc7xsm/hCfd8+gbY6i2EOGbmjjqrJ
N2owiM7WDOqkXh0sETmLh+6Rn7ySIPalaArPG0pd8+0TjmSnj8X1F+SatWiK1Uju
FX7Q5NdKwOr40miO9Jtq4habHuV97+ystK1ZzAKj7NPwfAFIrSlroXT8KZ3TWqCA
tk2KN1RARKKL+2fd9HBtAzow6xNEFY2apKSFJkXw6yh/AYaNYivbiUAUGiwDHfhG
zCjr+AM0f8iONbG1ZblyC2lxhxp8rHalT3UaI9whXS9HgVewSNwFBq4z3H+JSBII
uICIF5QirgpiVrKymieDfNR6K4V47BoH2njmK662vhzW+0e2qB9y5c5LWz/EM5ll
VRxzXivClIuxfu3BVUCKaFmz9Y07sEmvO0KTzyA7G7LGkSLuMD6m/4gN1Ug2cD0+
x6FnmxftBn3d/8H4HHD0o2Dj7107GUGrXU/q4/tL7KC2qu5A+GGMwgMmNAVyqUQZ
Bh8rYlZZO0n45foy91ypvr9avbbilsMZ35iBChL97tYhYXdXPELOBP4YS4FY4Weh
9srCuSkNueb5JgsuC2KfKDorAvf17midlkgk048Mmt+xUVXEfCWzwcHPoqUDyIrK
nw8RzTwl2S0QXXOiDu10xoaSYPyIUq85vSYL38XjNodjxNvtneTr2j8Qm8xwBODf
KGLn4JWDpkK7enw2K5S15gaoh6U8esPLnuxJXsBkxCsGDJkbCdgTjxgLo+WtlOba
RunS23oMd80HXegxTyMp3F/A1f1pnVV0TvM1eKGdE6uPmnXFjEMi9003SuxvlMpb
k9rPXxm6RkNMZJwUmD+3mtma+eSA3y11w4tkfBK5yPPKkKWekA8fTFoZbPm4e9ob
QgG7USLugCSc/xLwDt0BWhJV2gMlN5bS76yAWjj2aorfSSyVxXGGEOJpWmNkqOX7
NKoa3p2PRFk63BYpXc+PLKDf7298YGJuxnkH5H+his5jWDbefsnnP/KiEkSkwOog
8k6Qizgn0B2OXNye915Zcv58tWfzp4Th0xYflky0hp4S7WeAj4MF7OaC+SOD5ZCu
AuF+HFRTYZelMI8as1pdi0n3D6iCS44mOxd41TlOP0NXk+CSRqo4qZKSWqA0ER0p
HJwaSqIL7PhCtbVaQszTX+ZA+w4DaC8NlHChwP88u0ruDvrmVVH0kEcS1X6a1CCc
Nlyaf4G71jkuG2bzEIPfaxOxRd0U095hgnDhqSrKy9by2qy1ICzHiZ7mARl6jJgD
x/w/JdYb2dHklQlQou0ORxWU5T2xy2aJq7ONlbsRU8mGsW2cbNB4m3mf3ynsL58F
NoEhp7JtWiTR9OuMHexGYSJ6RDE6sxauumWMH0gMMs6dX0KKtpEE//lH4sO/bqk1
VCKcl4vlL4Ivce4xwH6JKGbmubuIDbYfofyqrXWzMlrh5ltS2A7FXR1YQlnGuRG7
b4lxHGID0qLz2W4UQ9rCB8DYfaHNPX8bSs154cpLUPNPJgLi/qHN9LGAr+ZyIejU
fPOm38LN0GbDW4QQ3NTO6G1Iaihe9y3aDf+nbzKrbjF+pWo2LKfIyUP47Vr8Pyo8
m72aKxTFgfrvxYB5tQiiuWScB7T5GyiVxwJcrZkfZWpfbS0KuDSosaMHNz8QdRik
hpCKRil3qv3pJnJ/ppgxHb2pWTpoJrQW1SbWbkaEogOl+bA161uxz1GkznuC7gLH
tSVWaW2yOcJzn6eXs6wwTuFCjvfEHHA7k4T1dIJ+o9FbBXGtbmHa5/LUZ5Qq+WAG
zR0Prj9jtmAO80smJUOivUvBm/A2chMDfYzWYFg1FdDwekb7gcxsjdGLXgFidPa0
3PPYXQ1Y19SAb76+7N3XoVrvQxU2iKFk7AbuFQMyArqKWvNYJD1/h8axohcB+SDu
eraHUwlgTgv+T7Dh9XGFqBNaZCb65KZrwiFBWcgtpgeZH+j2Xm+llZP/oGmAhXtp
LnRTzLGDS0sntDCtkA5DQOqm1tX7hlosEKkuZasAGAlQo8X780sR1lLPANHSUHXT
NdBftpDicTQO5XO57R6L6R53ip/hGWe5BIkFSM0BExJ04UO1aa42q91QXJ8czECV
7LdVtlc62sT+fLRIhj4Y0IkWatP0u9+ubAuErd2j7TJAqfX4DP5PLDw3ZeVVjQta
jH7cx+6zOL2XnjoZ4u1TEC7A3FYTn7zyF8XEtOqJz7Nq5gIQg0YVofmMaLw92T8X
2eZ2DIsUCgGyr8fdu5Ekpt38o7Kmerk1oOcInMmJhVGW1YeJ852RbLyrZFF8MjZN
Q6+igKdbCwzr8MFqB/FvdrPVZM71wx9u09jthY+zYx99g5jtZyIUq0F3NOH2Y+HE
OhDg07urRG1sfrdaSY8bQIX2HZLROFKhn2YdVUgxxsC8UoZqyLVc4OCK7p+Y+Ya+
m/vd2TLZlJTGBbm0r32M1O2mCMP5VrMgC+KCXJE8Qz2SKTk5Tmu/zM+IZm1bHR1y
fCTPuJhedXnheE4oFzRxZ+V7ECaK6AMG7sj5UE0CmBmXpOX0qK35WLNh2skV8QXf
Mzme8a3HsIv0x14MULP0NG/VD+/4UyTgvotoHc7l4kMT5dfKakDF49LJINHWQTd9
FxUc9XC6AlvC1J6RdCKPjfETw7O0N7GmtcXyPVZ/o2+0FCMsp2zLyWwdX4yaXuOQ
yBMxVg9uV//auxMt5cuMabbHN1mENTOMcZLBus4d9jBAbEEinX5nBke5LpUdIyFV
ZWtm2/dwbKFPLmLWjSY8TyE8rPmkx7GUTwqme7GToqprPPz8JSnwFrhRFAVPDii5
VCivSkx6nrJuF2XqJtlE4jZpu3Fujdhd+0u98sQmMsyKXBK6AO0Tu4Vj4W1T8NIU
fNEn3hfN+68Ek7dxJCDMpzsZTdw8hpJZVn2ufC7y7oFhvUKp8dVZMD7I0B+fOLvd
2wxRnoLkQKz+HNZG6QtDcLnUp4kr7HUo9UuredTaSw60CMSoUK4BDfmcS7d0ABfz
zTMkV1vOu0g6r2Jijp/qiuJcBOGn5BQpLR5L+um/e+CoutOg3xkvZwmo2x3vhTNo
FAcGCVasdckWoVxqyCSTo2bzLimUmG1kPQcPttmDx4A1rHk7/m/MpshivmP8MuRy
gN6L6sr7fWURbCgjmxht6g39SKgYL5jSs8UJQQ7BqZQzvYgXDcVtGqksTLZR3/Oh
ib/FZL9UnbaHpVGjSt9KsnkZwt0saRlAE9VES3S1czLeT2sWD/EjWBHO0mDcbRuG
AkYvOQJ+Tif28TdDlhBk5cHKSTfSXNbX/N7paFJMSVvg98ru33qQqJeH48UtKN6C
nUXLnrVnrkMrrWsBayc2pq11vLySq/ot4EIIGv34nPwqtOoS42MyhDEEpN0fUbeb
g7w9ZoQ23aEHyG3BUcc71H+unUwhyZzRiy136rbtsV3Ng3WQwC0Xm1xSSosqkoIU
1V+M5oGRHQSmYh9Liq4SlL7ZS6lk3kxyqZMbITRLZV7QZOtY5mcYAaHKMQ02RrNf
kjKjKqFh+MkdZ/kT4hYQtHI8ASJcHTtqHQxc0X6/SvMcXxeIm8N5ZAoNTrMFoATG
TvtAVEIda5PKqJNkUpVzVy+56jNaZ1LPjetbaXgQbZrKQ1mrGpmTSmFEsLpB81XH
Imu6ZeHMd/gcSq3XC6NzEV2GrwBDenmzi+6bqTNmTM6qB8TLWmi7EfhQRz+AJqg5
UV5ves1mKa+jl/6jg1tf8quUQ7n1qibB5cO0S0TR5YX7qA2KisyQgrNnRTUosfRb
A6SoaDwAljNvTGpc0xcU0J+LXQEa6iZRh1iPyi42/ZcU4e/VYFJXZHsn0u6kIcOg
80GoZ28LSPdqnhx65OWLHJMMoKoZAIW5oldAmbnXWywmhiG/fYklLTAq7NygWcww
LADiB4+H0c+ngz3VPTq1jKbl+lLi/np0y7WY9kJqglhFKaDOxfc1qdsn+8Lh6Wh0
TQkQBCTHEOz74erTl4KPCu9kp84VBdyHp18zbJL69ZUpMhGajOcrM6QcrfixNCy+
B2G7RtHsh2/2RVospNvSfUmTdLwfw5XYgpFYfMvRwxM5/hwrKOxBGgU3MMJrOj7O
vcSwyABgJTOlKz8XC2EEEr7VIkAe8/eml9O1dt8sxoG59U46+4Cnle1V0wl1CShf
ZTUpAawuiwDbae6dRmkyPhskvxaXbV8mual4fhySygKpHFDOY0jKXVcb/dglAjW1
5tg4qAil7Gdk2lELK9bmrUJDgIwKzLB126+aWITE5jjMrdrPV5MkjRJ6vSEPR3TP
Jar5/npDeAEj4dpe5VgpZI4UhlRvCeJRoWjIJ0fbG/5omSyRsnOmo+S7dhLq3H3l
OX0HuoN7b1GxTbrySu+UzcIGtsOohCpRSDDC9itIwLY5FGDgi06ZeAQq83pWPeSQ
9tdevfm4ZPyrNLzHM5hlLfmo8xrvUkrnzziBrlys24WyLskQsE+6cdIe66Uuz0js
6/b/YOyIZ3Ak6fQFwKPuzx6HBTxsQ8w74gslHOAMfICBhQIbzT5k8s9aO2Vd+Qbs
V8vuGP3L10+mU/zfE5oKjIHzgTzxqompYPND6n0ILoaYciJJDJIsWLfJuQoDmPcc
cFc2zUqPicMGmNDhC4nevNc/M6yrQVOaxBuMKnz8H9Y7geP+wZxf7je56mLWc18f
X/l4pMxlNd+MW4ie6F9qPxUTd6Xh9r7ZBUqHQQbaZpN3qqIlWK7YmthdN912pd4h
fVypGAPE76e3Ng4a9ZIAtiRQfdl0bmfnD/+B+MFOLq4wQ2rXbLw8SAo/ZlzBeRoZ
vZQWUYfz0dGsM6nuJ5HI7L2scJWuRbuDdYH8Xz6w+3S1cCuJDU8OV2zU+ETRVwtN
wAH3dNSzfGrLMgKCcyQPtxFi/0PkhuyMqV79IKvofCBnhOLF1s/mQ7fE8KEFAs/3
tn26gAkL6oajd9zNBrwFN61bc788np8uIxAL0VbNO6zhrFmeOb0nwh2yaNWKtkf8
TvPKOw/unrQsDNNBvfoFrA==
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:29 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LdWf70B+9ln7LS4LrhNXJo0Tigh7gp1w2eWqHJpCIosTL/thKmeqy7/lFLYJkqSi
AjdG1ps5HeVrlDIHClsRpawdlgh2TjZoIaiOvtZ4WVhDiolAPSwMMNukRBzr8n9H
/dVFOZTL8T3odgScVtAnfOmcNI8Nf8wCTH5QjM7s9fw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18320)
hovY8l4I8o313djNjOp1yfbRogqWiB+l6QMV9dNOGJ/L77LN0msUcT60zzScetuD
5EBblclGJdpys0Zm8wN6+W+RSxtt0B4rqr6i9VRjUDh9uSa64PnnbwJY0XOqVOyF
tizSncoib+hk2Wf2YdSK4kBHwsa+eGPgnNEWcOdr+PNFo9VhsaqTVEfhOZ/is/Pm
S7B3bjf0Knlfp5QmSg0TNRIe3jMHBDmJxurmfV4oX3eTfYpLicYr0wWfS+uM7UZ3
4MgiymNl1MvdoPAhiOfg5ZIgiMLeRlwrHBP5uwDQEed/om0cOKJeFhnt6v8DLiC8
Fpb2SPlQ8u7T8OEaJaITAYzELfcKmoOQ6eWKfnT9CdqejLVeKwSp2d1Fi2atFgaM
bJFp1kAG8WLoPjsmjnibtBjeqONuPjYgBz5t+C3D5duSbyWBVjVw+hNgXSer0ejf
bU5k2MR3dy2OWOEVUzsotShBjWFQ2b3wz8Ya/1wJy+bl5slqDwFp/tEi0sIKwBgi
81ZXHwwn7UtvhRTtxBaLEN5nM3VG/H0DV33y/OBKZEKIhaF+DeXdLUCJWwIETISX
psYMcBUzUfgvSkLtcGHg/5cYogbMxe/wko5wVv/ERM8aCACuewVOtKdc/PUDaaeu
foi0UvEME0avvASIzEfLR2PVJwDWnWYccZUcSyN/ddzy0i3ta5VBstBtw+ZGV8e3
jGfYWhmeB+D0ltIJG7g5U/dDdumHOSYKwzKoAspyx3a1wamwaeibE6NthNdoJFZg
1DEQMMAHulaLft/4emf7BbkxdbpSvMPKUg3JdTBhYTmU2Y/2mxD8ut1AFpSszw6I
X5IxEXfOr4EDzc3vn6wAPJlLS9U89iP3BUB3iUxD1XlvP+QpTtmdbpS1iHXhzA//
jvyYCadKdgD9uC3tiEdkANp5t7G7JudhnykwFvN7wv6w+nEBOJigcGBHlu1FH631
kpXtydTq4vHxg6n4Fr2mlfpAv9ciAljZW1HkARh/h02kmDt5qxe26MPzJtkI/ksu
jEdqkQZnuepNMExkxyLaGEBNx1ua0npyLTq8iIxPT6W3Xa5X4cA7DngAV36NNSCi
LOsAodOcrrX97mPxzsEbc2wlvTcI6H8QFG3wa6T3GXar1PAGVZ861au6m6gtXTUz
4UmnSgi4L1lXam2/+Ap78aBJyGCoLsThYKxtf7m2P06bxUtqWxXuyvrOY2wzjqEL
XHqB+WkeGnnzVi7ghhuFupUpKsbQSwRPUlwfei5/cOMeVfld8FabcTanJDkdH73v
sVdVpcks4RRYMGy8WoOKBl3CjicpctAyu1EvtUsPMMiNarzOS/bsjt6jnM4b9qJJ
VnvXNsdbbt0h9ssIWiOIZ3+AefC3Nu7LNesIo/hEJfJs7VR5Y5X5GSg3OtSrHy/E
shyZIML2fN9LGb+H3is53pN4sKJ//cNUM3WdNU0GPcnGNnxBAN0KXlwk+YKXYloq
GHhdrXKvlAbtkZXfPWchu5lzDkLd76oK1uaDEcYGXfu95M0JwsWNJeECAbCu/SiM
yni8QB6GxCuuep0GJV3lC6uTR3YRdDXeZnrpVsXK0B+TQbRQqpAopIxNyck0JEWa
V2P9/vT1IJxNal9hUE5XdqkrC4g2AaR5Ii2vmp1bPbfgLMMb+GAEUFFnaabhG3sM
/jIrDO9goZ+sNksv7/sugvxenun7PPmOwYUsA/DKkQSlAAPBKZf/nUZAl4MZFPw/
rHmdDPYeK38Cy8TVitS4+0fC50gDICP9J8Xi/8n/V/QTiQaKdIjX7hvX+Zp4dUgB
cKziVfK0NsBslKl+FaHHVo4j0DFRe8njnyqkl9C49q1nfcSOjGlogFioUuOn2pFN
1YW4tLGw3IdRcm98DXN4QYAOCznbF1WcwW8AcQc6mpEMoWlI1MOzG8u9f/hc0q+e
scIBdll0+KQ07GDgH18n3aT7fEOt0WbPvtwTnT3SzG3BqH7DWw2Kqm/d/bd1AXyT
ylpeQOU7v8aq9HjJJ14of7IY5ZMPO0VjJuN4jGd40jZZt7SzsQexOnLHz0Ty2JgW
7Xvezv4FGzkfnK8/5zXhc9fj98HGrXhUMwU3Uizlq0VAuSTC+BZ64mNgERsHbs5p
7cwmEJXZYpiQ4N/jeFSd/C5oDxxbPqLXcoH6GYqhGmx09bax1bTdpFbxbgeVrCZi
30wSkNwt6cO/IoFV3+Ikjo9phEs2aeyW5crDfSNfDoG/dzzaJrTTIEmn9bYdOWfD
i1zwjfHKz2MHboLJbKgO34x+S0dH7wfv5eYMQt6yAmA0S2tHspYpURTu8F4lNt57
PSZf0y3Tie/QXyJtmwGIEU+yJFBTixOk/DxQDU+gC2xj4eRq5dRJu+oMFjbYjmZF
sK3+BxbL79c4sqBZ2QPJ+w7xxOWNk1kW1UJ6BGdcMugwxD0lshOE6xuaChXV+BvI
yhXgZhLzWThGeogSZxpVly6upyi0T1ZO9KlXao78V9U8lN8RHv9CEJZ0ylJcV1R+
E5od8qrtsrqDToqi/uGD+NjROohV6vz47R18YAYIUhE9HLKHy5eRN24o8sUz4Ajp
aiDON2zB2tAf0iC8Dd/uProhL57RBduBcOpH5aqsddp8VmEGUyKdCaLvECx84NO/
uDxZq7oTDAqkc7/QnmIAFkMr9KvpQrciWaJQbz7wmpAhIc3SzJO+yd0dRMWvT/22
joToqRazMk4BmJRRyvwyC/TqEWsNfZQvumBD87w4WJe50698LwK/TWjySmuw4Cz7
VEW05je+gkmyH+VRg/ni8EOz0onFKLeYuKUFVuVNVGTaJouhahUZA7GqiT1tR8B8
4HOD/lnDHIT167njQsj772rf66zvzomSAXKgL9iyIX4NYNoy4ubURzPW/CkQBDk2
GnxASS/A+nB35pvzP00cwyzDCZ5W1mGMU+1ulIF9fzEWKMrSZpAUIQZSjLeHMu0D
v9Bk318yVzDkkWhwS5YusL4glnv0FO9+vzEkxO20qO+NfkwcCRN5yh95pdqGr0HG
G6p4qqJ/d80JhDS7cioEdufUH33nU5IdzGakI7l+Iu4fkgyhpSvvl0sAk5rU4751
KZt5upOgG3IJhiP7NflMdBQziZkls7O9qBZro6EnDMjGxjtC3M3UcICGK44874yg
SeDOGX++NsEuqHDiWbqDm9U+MSXDhPxdxWL47lzgVXKJehuzy1SGzXIbITwUlgju
di11MKxyKb8ZwqYL4nSkGro092mHzLTrYkhjfEpxm66q4nTZMaGL3g8YyKUzwFp6
y3GcqXgFbuHgoC4uJi0F9fDvY6m/THePMaZqiNEezvuilglFkqHD5cFTTphyV9ir
leX/eqF8oP/99AiPtHaVZFzsR2gdwS+AnJ+B2p+m/bMd6kD6RkWzAZLGlu6mOloL
qWvlWD5iw+i3euofSfjutBVRS3dhXY3c4R3DVftVnkhN9cYLV+HzY6Wnl2TFJVIU
nTQcbcJMjpQbVJzCIozMtVjWHsYROyNRjHZj45iswVQKquPig2wtFJAw2qKDcboz
ic6nvHlvnd167ucH5n9BDunVUL8WE7t074gTz1O4nMdPU5Hz1smgIZsXUjEDhu5e
KhdVRWXWYCaSYG0IUNNjvnx8K2t4TN8sc+M6eoexrADCMPw0PkppBB7I4RCzOU+k
fzA1SGHo+3VVuvdTQL2Phs+gd2Zh0HzXx0DJ3FgbhTXT6SPePn29kEku6DsXJlhz
s+1Vgo0RQ4z2Z+Jjd095oN5kXZZsp+zQpJdCsLvleemk7fs0GMpzbZgkyS5V2nhM
udQvJsXjhaBFEfQy5sQoHkjp/a8XDwPNLpzK42PjiycWt0ClAMJcqWDEgpa7yUE4
TMF/GHNuUs6Ngptc9wMwb1oT1bOEpNWj6nsVJSqNxF7QOB1PtApX5RojVm/+syq3
JXPT8VKCe8H7HHNcbGkKQEUET4sjGvOpZeu/CblO0kniFFYnXIWbZUEjsXlwgd56
o8spCQb8KlfOxofTCbh3dW4TcniU1QOXML/9yRzNi8iElpzW1EoQzySZ6DQMFwoX
WL026O0m+oJKum3nokwcyqLLCkgDCQdYjqZOlfT1ZaSHWzP9gdTBCSTH/mrQ/HbM
tzIqz+LRtANNdOkISPcJhK9jokO2/F8mO2+Nm3tqei49LpC3HePz2nnJ/+W5MAvW
Ym5gVUZ/NO83JhVSEpjjc5LSAlMFUhT/GGZgnEXY0mELGbXGiW7W9XCpBxVYE5nt
UEDBxzIVxjacD6opu8bu43b6jxrBHi614S1MraaHpkAlDq9KA8ZeqZ/EGSsTZwn0
/w7eH0ecSu3iGllvTLQB5G9x9s8qfuZ0LoJ6hxWBFBDkLKhkLn/F+hK+kwzirvnk
hTkkrMXexfkl0MVs+6nDA9Tj591icfY1DU7IKW9neIgFQE8T/2BCKoX7HYGFcrWn
OYFQUkwTqvyZKEEphKffoNBNrlJ02Jo8quxiBGDQmIYs/9QhrFMjx7ip/Xmm9A0i
rrTzj5hDIRg7xgp1oUln67uPkTj7aJd8D7ja9F1OlLD86D91UH7OupZtLxoBWKne
5msqVHqU0WMFgf8xJLfCQqVgjylFR6DeH0RFtKz/hn6EUCfxxGVu7VXFychVpLr+
pZyfBCFw8pwZsAnl70urnNzrNz8xoCt0N4fb068D+ekjRH0bbYWcsjQXpDXLhp6b
SY9nbYwWoUHUWiY+owTx+p8u71jxSYCQbhvBtNFa4+vMr6JyqjJNIVeKTz1n97ts
/VLVA7dBQBxMDKeKsRPePpXuVvMp0woOpK15SknxVGBUK6APrExyAE8BWEEv9MBu
ygWfqjGvT4i+CRVC78q2oTPrHRDlJLY7CX+TBc7NBn2jgsS3l+SbDH1CHHsvXEK+
cw3KulsGvTlw32GUZF8vTpOcbf1sI6tsieYVIdjcDv/GgUfTksxpTW7bY63sVHi9
LrDfvhMqaJrO+HgvpYZji5KKrX2NRu+I/ltTbNwATPKo9G4aItFQ30Sph2fA3ACp
vAMdnFly/Am7i7oYHUD8kHrcX5s7QVC/ETTxtUfXDS1hoMlMRvfK768/K2vA+GXs
WCX7Du3wQeORH1iTPzIDGay3jmNRmX370GMN3C/ij3LAisI9yHoRbWQjCVJXoRwi
U2Ylj57XwOJdT6I/ohplKDf4r4puumoi52Km72Dh+MFPjelMuZ6rktCqpLxVbawx
O7OYmmNx2HJSy8kk6kGxDLVQbK6P3D5qDnOQyJRcHfBm28EJ6GUiUjGm78PFIED+
w3etnlC9zNgq20Qvj0AN4HTc49TorokgNLN2a+E0gMIY19enXa+dgU+xuPO92bNF
mm/17JhHCjBU/2y+qrY9k2FB1ooEveCcO+AeJhE9oDDuoKWWLJbKfdTLC3WGHIrQ
XOq7jRkAFoa6lRKJ5BhWd1VDgJGwAvHiF4rCgoyssIQKtXkfgP5Vt6uNagnQVBhV
7d5/GcPsedGqJhNOsM3X0s+F9JoVeu88e1+lFyPaD/HX5N6XvOLtu+6x+l20TuDo
XAMHE6Vu5XYXlXj4uCS7Xq4+KBOPNhIXiTTwVBe9irAhQqf10nqFKfM1X238NtX5
cB2FBr9fntKUU2vRjguVBkxylgDJ06YMyRbP3ssP5RjxycxizeIfuS1UeMbumvj2
7fYc9LsvBGUUppy2bhl+IiuGFltWRkilmi5i8/zaklD7RnuuoTBbjZ6ypVCyALbt
tR1LwWFhtVfaiFS1i2J0AW22yrJdreYnH7+e0OaMaLJ1s+Y1V6Y9AI4FOhotwT+P
1Q7Ntqe/PikmukeD8j7mndUisXrBYPKum/UzH4aI2VawYm3ZllY2PPrgufVnr0by
YgyWMnB737ofkHZ2PABlbkPCywnl+pDTy9v3/AOOg8fhi15W93BKjyhZ91xYAke8
w3Kr/cMf28B3gVInP6vqUqA29YDqGlRE1bJKbDYW/8Qhb0HsDAi88UzUGTNCt6kq
RLEx/6E52KlgrPv3lYgB/Nx2ovYnCDyG2rY18Mav06EcdarSK2HfZkx3wW5MegeB
ljroMKsoTn+BluvQvDNq07y/cAtp2R+xIiAd+xzLM4dXRLGpcaNpRbcLDmUxIuUW
IbutfvqtVIrH4u+CF6ec3Lr3NhlaB2E4KEY2RrkJouJ/pCjJdyxrR4eDkTQKZw9A
e3Ka9Ucvwte5Z1wyc3knkImoC+SSPEFt9BQiNHvZ91ooqrLOSziFCTjEsIwWClqR
AtdtQiAEGgMpzgie+cKhjkagbs9qE6Mh90cJkXsgNNSwqVaR0wGCfqJwNr5z/jrf
/IVZsFWZJsaalV/xoVDtXYqVjMmJxRO4cUHXD4MNqAp+EIuiQgAhktXuyI8G5D14
Bw9kBfHJI1g6h3NXZpRXb/u5CIY0yJC/0tlKigJ0GgDn5FQrsagAvEoOwG4Hk42O
uzZHbKMOb95VZICv8Dy/dBhttXfEyb+0zOdF4eE1199ehKlNVIKEdsWblt1bnLWI
hZ1MpER+6gcpJu5isfth/w0n/R8GrcBAuIx+G1Iezxd0f3hZtLtMBLiziBj+gaPu
wWhbrVnT7Qt4x2L/IiOTneUuzrYCK04lf8yPSz6B61QsWyHwoLnpnQ7HxdGldoB/
oEOvRXKc+4KSgwN2k/Asshfp5Tr6Zt24rzIh8GyEDzDRPOMepL2sOGOn4BK97boE
aw1RxTF1yijmM5vKHTKzRHV7XurKS47HnVcIyxeCPT/4qZTRlJf1rH3BxqI76JEU
eA5mwZMOjukgQBivQNZ9grouEm2Xrk1/YADRHlpVjnXIFfM+OIin7XmLpXyZRH0D
r+99p644+nleeTdEIP4rSkssMlatrgUeHd+r81JH8LmUdzNfaZoDw7PW7o6QulH/
YXjGOtkNObwH9XR9XgoSiZ6lmC9OAsLhnu7KEowX1JxxyTk+GgIxfbqFv55AY3Fu
16zZaak6quMlJWb+JzLJnYA1x8mUuZY6jWCkIwmg3lcViFUMJy31Szp8N+6yEll+
V4449YaqMhJnG+uV36dZd+c/CVJIZjmnLwm50cc5w1uD26g52BTcwyn4ENMgbFNN
LccoIH/h929YdQFlPdnQEKrCqy1BN23fnI+W47m/c0enyUiMTjVolQUJQ0Hze6vf
M1Y+bjgKEyjlVeb5BMLgOkEv+85WJ8RMzpXoo1X7MRkSq051dBR3y8VwiKzFsbdw
KPlUYqxzoSIMKlFmFlDpAphI2OevhL7dfYRP4heI0cJn2/PwKJuMwRL2TrsQeT/k
dsyxA7NXv0mjhVEJli3Q5yiHf7aFZvmBRKzjpafBt9lgU2/CR23FPQk3t6V8IFIE
FDPoWM4Xoi3y6LGfSTbKm0voqo/Mzljds7N1ZlzCYFa5MH/2hqEuJnKLdCDbuk+D
2cIEpBnjvZ+1YD0fBsynqyt1yZqjdbSQfW3NBKcNZU65Am2CWZV3F9Mva2ZHlUAr
J3atebMg8AZRdgny/yHQFaoeby9Hy6RHZeQD2qLSHVfe70aMH0jZ9IQE6TrtsEH7
/+gglZTnk52sM7geuGEQ2Ffs9Vy6V8s8xV3vll3n0R0oKlzDnJQMvIjuWeqGOXdD
IpZ9JEPZLy+k9hWCLWvZ3cuArt+QVGo2fdOUVSFA4i2gDeTjPO4T0gjtc0NGLVMP
GuuMcQwpmQNMJ2EZPHBDJoolaMOVMCRznrPEeqtGrVfEP8KUvWdD4R5oVOYoJwb7
soJEXqC8s3qiCL8A8JHNiurh6BXjqzECc2swyUZZWCdVF3H5dJsQpynzJ0O471su
OpSFszQmhMCWOlqp8xxPDjbKSPqqhya+u32ebUNVxBQuitW+r+jo6Sru7jihHI7L
LeI0NCxkHZ7LxS/98Uzmb8/50VmcjuRjbUqCeAkvS9DNEc8PxLSnj9ZScS+4a6ot
3/ElW5Y9y4wljW8V+nmSAn72kqWnmlAS20fvqzSFkL+LJFpbnThBQWJf+D76i50G
AK68TRyXuTkFGEVB3HNBx0gfS3xp9ZjPTp2IjH1QId603y/IuIJFzfXgjSzGityO
tQxmGpPDnzuMiemN0fHCbmLLzVEnPiys9Re69n/Q6PgxNZRhjr142Fg7WdMGeo5k
J63F1Z/PuMnql86CdferiMi+4+0SagDhJT6ujor9UBP5FvkHCK51LD9/4K1zF+xP
5XFUCFZdGPCFswxN2RiIjQ5g3MozuvrvDGlSO/k/JcKoVovDvWKK0KmmoDjKELxr
7VAwzrqSvP92+fHjXeieVNJ9yNkMVux1WZ4zuVD/Q1bvdfuTkLoojzN/vgREzFAN
TWeMaAFMhIXUrH116KGpZQNsqZWzIXB7I10vPA978p1ug4k79jMlNsSuHiTRlTtg
pjDEVlsd4sN0HS+JK99jaVPx69qnax7fquhwDhiP4JKbPYZFXHe3Tw6VIFVsMr+k
0HN/z+dSjmLntva6x8BvRamhV3dW5DtTc2+GpvhjzJnaL0BsFqHq/UuPg/6v281Z
OslHBUuAYdg3SxdRTUzwsOpIGUlSU9ODn30oKN5KWrczHDcl10TcHPLd08/Z4tMB
vkH+UYD4Pex65DChKun2GkgtPPE2Duv8c3dbIa9q3m0K0l4dKKigsRjW/5/31PI1
dUtXZoVl3GmteP26QqyBjREQnD0QD6Dq2TY8uY5n0WRTCkEYTHteGevaW010xP81
s+AIZihfj5GXhFDcBdJBLaa0vTh3fg/4YZbLnIP6tQt+vyllcNd0/p68QW+Swkrg
5C0dXZRFn6ep9B2fpywybOGADeBN+B3I4R1wcV2zQM99shdpU5bGGlrVcLzsb/BS
/IpGu3xlUzV0vR4RR9rGFn+YMCKTTWrTeqh4H4yX1Hk0bQLNa7CsWNItrf4zlQqA
C1ETSltvAXIv77k7Os7wsXxJ8OxAlwcvFox9nT3sqbqLNmQEIiqv53Cd17SIsWRp
bW4msT+w0OCsylDi+29zEPiftE2foIswW9u2x/EPdICYhBGDfwi0n+OgdPXUsOJ5
95GVbI6y+plsdtNm/nAMD5+8Fu13jm7kQF3jZwP6ZPstMpMpodt1oROzNFeWwqJL
mQd2GlRonthTnbktKMxOHzvrHTqsXzZMKtmavc+J04go/8EwCl2JR2bagosFIFf6
a6mniMAAbE7CbE3O4fAHCQWWxad+Yvh4m2aUY9jcuL7RMt6R3RRRJF27dz8TIhG0
vBPFbIKi7hIDRAkjmDg+ZZI9uNsCX54v62f+9ixoHmG+Wu4LsEUVqdZWCae6kKhy
Pz+j9oyqoChIae6jVwaTUxcm0rHICxUijH/mSETszRntpg9QXE8SQeZzKOiVXbGT
YemoRBsciyJJO7h2T1IcAeAGEYys1+BqN4kNVdjSQYom77lJCWZjQo4YRkDtCxmK
4xF4hRj1tGPJldS/fMVzGp9BiNiI1hQmNKUoBcq44iIE0jphB3qyP4XnhAH1dywH
JIP8cWeUt+Gzxszl+hfbw/DfiOQ2hK0BHBtTtyOUh8G1xgGUXQ/cj+v5CnK1InV8
6dK4QO1cQ8JNp1TtzcOeDlMttBG1evu2dimXWm78VUC49/hUEqhNeXo1CFpvR31R
Ou2QWra4ktCzJrV5bW1C3aq+/NU4aqnX8I3vToO//Jy+23C86aeIm0ItsIx2BOsW
xMKM7v7q4TycHOxcRZp/jcZxEHVnCGdLFAHDPUYrVmKSbur19tw9ildmJPdyv2Ej
R/CokQb8Y4VdzPNFS9hrkOoxqtZfIwuOC/YM6IxCzT7ahsBUYoDruJSwTmldTNch
ON+i1zdipNr4JzgxlNww/rBRJmP4aaG/8jc96YvTFqSEhm7RQqMAWsCuIcBpISro
MKmHCvOYWzU7yWofpEM9WDQ662RxjJgkF03kBQdNL3y5ZKwKkkHeV+ERaPilYa0d
d2l/jcTLt3iDW8izQL2SsRscgdAVxin3DbMWrAo6fiGkUjYwPEdcV43UX/dE95eS
nco6Wu7aGVPb1ta6zs5PIszn8M4CHait6QVzl7ElphwMOTTn0WTl0ItmT19MrPMb
Ola1mi/5FdTXyY+2MV76FvRGz3zinu5Y3CO/NpJ2BVxd0o5wO0Zflx53sLomVkru
9WQU7r9k0CSqWmKSza6JGOU+NCYP9Cs3kgWK9qSy03Y8Xib8l0ULKuFgMdYgajTs
gtceLPNxLJXsIfWeP59rsot8eK/iB+cGWdsbfaRC+Ac9MP+XD2y6MyKREKV7vL2q
eYgrvCadjOOyioHdlYgXyyf0UxL0JmP3FI+bubY+/skcWm3VT7QVamcXwZ8WNxK6
K7LJxDvM6G77pdLzZRvCEccovYR56XG226cfbHj4ihOvHkrT6lFK7A6A6WcGzERA
e0xsG5suJT0K5+jWKUD1Eez3LxpfVKiLgk44OAUTfintOC+KVbtUD4lukKCoc/kD
csWyYYOwvCG6n458QxhboFzwYDJq3dfLPq9K4QWjmS8mIVTepQiifXtWoFu4RGwZ
hEtyKCU/Gtcfno5KxQzPzsH5PtQW3iEanKTLlGsfrtldAORS8IGkHdU01sfdEUSx
onHvbnHAg93+rCO3+Et8YHzmpRDwaCAXjox0aKv4us5Nwn+PGkkL7d6CCInw7flg
qsCRaoPTTlkTL4VwTS5Pd5Tm0HZujpbQzxHNGjuHnqVZ/D7EELa373pAE6g/IRux
mC7porQuhqql5L6fLO0Ht4rFgAs5sF8ZV9rg7xJZEVmjw4YPNF8j1KqEaBHSRVXK
brepdWBo+JneSxe4cO7pBtY1gpkcsV3UoEVlS50Gchg+wmwZwHFKwyEciCuV5eY2
7qaDE11riOGqHBTZAUvQXh5u9M3mhulHzvEUJxpXO05V/MIddmVSvb0YxeA0r7Uq
MBfKaW2Gpl7mjEFp4DgeeMAKM5jFAYBT0K7x2ze54tikIDqnaNe92q6fNDZANpoZ
s79A3AMh1znUOw5Jy1+7Nfao6QWOOyJAO1e4i4vWDkTqp1V2BLehrwnE9HkwRioO
Z9noDb7ONxzDW/CVE32OeVifux6DnOdIsvyp+cwnJIbkFCk8QuG4iJkeuJmi6iWk
hqky2n7GpJ5JtUnWZZZnjEFzKOMKg7t4JNI5mHYGBOA7gml4+euak/5eRn/RJ0Cj
qqc5yhiZsMrGG+MZGixhS/xi6MMg5hagM2Mn6utGkp3xHcHH863PESBQMNHKE0QF
YnxQgyAg89h/QjW0qPer7twjT02UMaohBfBoDi5obRhP3oehwN6F26ZWEBQJc3uQ
fgNoDVNfdA3bDtcd3oq2TtxJRkbHReYEk+zH951ph8bzdpGz1Lu6wzsmsNkcqT+4
gnDymv2dRNuz2KnvOAM+plohv5sK5pwFo9JYhnAmvHzU94p9Ob4ZHzyglAOJzfkq
MNYJNxg0t6gYrjHSUCvuwI27hvTZfddfzWQz+DFb/h7FiXRc4OIZNv/aZYRgNdQw
hKd6m1QyLOQG+GPmVvix6tz4u2hb3+B0ug8urJ+m2JOhZTrUGUdUnDOggqKESXMp
Axz5PGsUWEIEivb6xje66/o2HddW5fqavMD24bOoAtOHVdLdrm2yKuchKqp8IDLb
1coqDVft8haIMFA+xkHxN+NcnaMdrHId3BkEKmrxTurLV5C8727DsHOMwX3CX/AJ
iPV1pPbeDkvwYf85yHI+MNyZ3o5fXkF6Tx7zy1kqX6bdoNFYa5RG2SN8UmYjDZuT
+2VHnVhJv/+F9dhvoU0GvD6xmEcII/uipNpX6I54tPBrlT5bypm+wPzhDnFuADr5
mer+UckQ0jwzZ2mMxpRo6nHxWnM30SydBysygXSswqE303HRU2uOK8Ftd0PWhr+M
SSIgAt6ODhFPckhPDmd53Ik9jx64WCrh/R5JoGZD0wBOgo2JN97wwYvgv+RouaoK
8ohTaCRj5Ysnqx8LofCdwzDtrXlH4kPEJRHPQnK1cR+lxJFIMxMTWDREy1NcgPY6
lhYzlaPhLYA7wkVtD4yVxG/Xh89Yh0JfmucREsUzQ7V2FcLv2demsugn4E8eDmad
N1RBXJxXmAlF+xXQ2hawI46X4HWLX0Gbqa6jt48aIANZ7TzNDuLX9P37M4lGxUP1
xtXmK+ArNElsG7yCPpbhPGuBngs3NIXcB8ai2Dzs43gViAGRyP+G8xEGox1qs73V
QbG9j+cOHxrJDtqlaYmMIAGGYHxzituiGfvG/TG7I5njkaS6OmJ4Ed0PbMuDiSIM
KMY8dOp311oVJ23p6GaquuBtzFvYEJFyXPeZlBTr2sIZDXiqBjss34+bSqfJ7yqD
7hYCaWQ4bGsIZ00yophko3Vx76A/9rBNem54OrWSsNHO3Y1gMXKpuybKFTmTHSI3
14csfECBPu5IBkUOU9aw3E3zz+astoZKRH1TmEUJfC1olYj90FXxKz31TBr7kn6n
rPdI64jNl218iLEMg3ilsXy+JZIofa2ruKS8OBA3xBoN8cyH4Z7TUA+rPRvOm6YB
VSYr1v2971RiN+Vy/sz4VTboOiyupiVBA00o95KcAudQ7v3R6NVr453r84CiCrD2
ZZYHeAbnZOJRbg2dnLLjevp4pHJv/9+JDv7nuTeauHF3idBDpU5Hf6DxRlmvnm1d
Ukxwg326bVBplvUm381J1WErQxM8qfnAgtCiR8t9N1Gn/Xw0/4t92BcQ4nM/dV7w
YhMObgyzOYEFNH9U+7RGcPlE6ScyWFohXl3WsnRyGxyKuRSVhej0loGunfT84qee
2+l2FOsBTnUVoJJMbkRQkuKjtLHCl3I6rNYCRCKKYSw7td9wkX/tBik88Zpc5FV9
6cg/4wfJ4HuURt92Yx/z+NMWc/Fm8HKd1iNJRr0EVDEXKvlL+yp3ETgw+feUaqdX
jWlisMKh7Xv1CizatXe9hI7nE+PiVKu9QQwguBaxFM+O+0XuEEOOnjIZbhPP+KbL
lm7Q4pswzfudeA6OT2doydqlSOYn/ifiDFTA8Q/SnRgDQTbWb8kYLtIxBJBp5Gk3
9R/EWr5YQ8vRUG7b4NYvrgz7qTMN4gUSkB8YSMpJWSpL8gJDL5YGlK3UgVWIdB8y
C3bSN25B9y2dksAWBKIhHVC77IjEKprYb1bTMtAtzYfaeu1C9PwvjQAdzKgOyyPW
zfZKJgRIOtCB9jxkrCj0tbMOoM8echcmh9KayjGGXt1delk3BjJ3TaQVG2hE0213
GN21mw7h5eDjJEmJOBXswrDnGEJdMxvt/dYVR4lX1bxVM5YFxyGSbBQeC0Z/n2EC
oHk9LNIan7DEStXp0BEtPuuALndhdRLQMBk/4bWzaKjKGQ+Z6RVjISslqtKR/BdD
3xrZhsk6NjxXg8WJHDzn6Pzp8N01zDiG4LpgISjshtf1nfNI2x0G4ZWqOSpWMdY2
GyoY0E/habVM4SXXim54lkCnvCHLzPR1kanCPCV2n8QMWJykvqe8RFwXSKN0OCaD
7WKrhvVqVnDGdIIh4X0zzNraygdIHm8/Od8VreCkm+o5h86sa3ccUOPMTnrTYH0V
Hidm9Rr/eAf63WCkEWoSdb9wTQPMGkwdguC53q0gfa4jAYUcitPaQmPRAmhDb0Zk
fyIuyf935CcnuDvkDRPN+yc3Wcco1UIvIXnn02ySLfyRlGd4sz7iRRNkQ4brgI2d
2dGn/Pg2Y+92Qbrv/tcSTjO9rM3nujAWtuha6ooXauuR2ukKl5YXW3nQYBGTQrYw
zWuSTnhRop1QODJyzquvGU0tT5zMlU2otLOftr52sOfnOPhDrok4OX/BL/vKopXy
fasejNH39kJRjRF43uwly99tenUGGyE5vcYX/Z79qXHKABcL+rRWV+UT0Q2XKM2T
+nyUesEGj8reVuQtvP5b/psqO8gU0T99rKbgUuUz4+AJRvzVa05r6aJeZ9HgAAko
H4zitiuEsyG+0SorFZTD0Gh9tNB0Nh5+9oIbSmCgegvbMHJZ30YQuqaWmIXDe8DP
53EZ7EFFtL7mKmdS+am5+jCJYGAc8I21ERqALho2riy7ybDeUN32oL7EuM2stVYk
6vWhuc9JZwqXCEw0PvEZzHecgfm3TYNkneGoD50+Vq2HY1BTCmV9mkOI+9Te2suR
9uX2+DihCTZK4kku9mnNq/IFFf4/a6AEU4QJLZCNayRl3B8qZzTkQ/rBgFNB6tdD
IB+YUDInQdYMB+zbySRWOybxSXMY0V6P65TowZJwAAmztEhiVJ9RD5DTsA/WRLkM
LLR7u2GEsqQ/+mesKQu4und68xeEiryljk7yfErq+skEjpcVTaL7JP893r6i/iOs
b93FFCh+h/PumBGdpXhC+P2B6gqalQhrEa+mMOAXGHvLMMUNlU/d5K+vmh0IUfl1
H4+GvyNffAch/3dZBNI64P8CpyiO15e8gQU1/u8sKMUk6E9+TUouKsvVr6Rt7Gfc
pp5u4STXNBMTzhlUqF3BYTfP12krZVumqNkto4m5yztrJacPrDyHdgy3BjtVz5V9
BQsA229FzPQuL3zxGb9l4wweatBy+sVmZLJdijPGPzKPSegItSsPo2yBj4wL8A/3
95xMP83xjxWWdWC9HCg+B8Q4hBan+3vEATm3mGF3ufECdaa/swC7E31tkLYjqp6r
XOvgh2uIOohScJpkLSeGJfawUIfpdtAJuk+X2OXKrR8N8dOIAulB8cWK59y5Nl5c
fEXbYd6oCGXj0e+AD6mhvvorMGf/oGBBxyRcbPVKwqnfzWtQPnJaBRLaKNbGG8dU
gIhTWvWTBVzBuhyNnJiHiqs6pHxETqEr0cIWpF3ucn7ZPdEAIK7qewG10S5bnPu8
uHUat5el3lysO6fUts+PhDRa9d2zlMzmWekl0BDuWdKQOBK6iMo1n0r6qX0S2MlR
XrSxrgq4LKn+6Cet9AgqeFUHUXQYXaDjKEa3CWGw6Qb6tkW1Qn5dNFGCIQImieGZ
NwXnkibgYR8Nhaq/Y1rDZZO5fdEgQDFKZA0+PP3Tp5Kw2jZnmsHLb+CeiOhXNH26
0voMbD3PSnU/x8zSUCU354m6IwdJM1yHyUsB03B0Akx5AFV1/PbcZvlL/EaKnGnH
w6hl9T9wlUy0P2z5eJmHL4U//ORo43rLE3K1DW7XnLPXZJCm2OCihk/ytshErJwo
Ukfgz4kRZdT56vheJy9FwH0CL47YdBUt2u/BbWn3UTXJrkYxNkGtZySfFsGRw6yy
yP7KQ4JD5gqQVODmFjTqlL24GfGBWDkFvV6OgWL2tHwtFUlPVxCmnhWZFg2CLh87
EDzx8BBSN5v1ivXiDJK50Pi2dnrdICCcwfERLogji5XP2rcRsRVsk04qtXb/KroV
qevcL1HLHfSPxXwYv81pqPOXkQBD9lBMfH0N4ffAiNzCrU27E6Ey/QASzZ3pj5Fw
IUKlULF5bovQuLy4Mg4B+FWIVxstYapphCmvDMayXKyKe0csELC+gndtcjpFa4ia
NQi9vnZQACoBzc3xHucxd3KrkT4BJQ3BacICOK7FzZKdLcXzyridxZYUbl7QovPe
gOkSel6cW+wQFMD/WTASAj7f17PKKuMnRp9+mdGsdtNWx91A3MLjsbu4mUnqbSAL
UXOw+0eXgcXq7z6KSCvVj6pKr1LH3TevkYi26YEeO61cqd1iRW7RcYC2cIwNgPHh
az76WanlPaE0G2QPq2Xd/mIZVy5s73TjZS/ix4SueVvzbI7r1Kq2VlLtHdh4mPa1
ChVm+Go7qknUcz/P7qmnr4g28WmgsCWt9HNDjKEd+m90/BcnDYw3iu/8/UbEO58B
/iVxKmg4yXIgftfrsvItMywxhLltsKm2aDRSNuqP2lJDH31vzC9RaZi40ypM046f
hq590MHAGNZoBlMUiT+9vJcNJ4gZK+MgXvmyxdQOOe604crQP/I5/BxfyydHBBHJ
RzgdA6+cn2K/OaW6Ze9puvxYa7Qx9tfu+4VVn/rI3MOLhcThELYMkNtPrjytNbc2
Pyf6WcaiyEst2NVo/VtljxbSN2zHWn7atAi1qeIRFXSwbXMu3gXo1FDb+AFJEYxM
fDMNdpBGyd+/NVmv3J10FFeHESikOcxAStf8B5sPsMfoNvIt1pJMHMSJYvewQD3C
fFjht5HtCzBqXuaRyfDVl392OJnwbcRC+Gwo5qKeuE6UBkjQf+4gAN1h5kS7UeQD
w2VRg/yFgLTrFAfEEEH8zVnMsBxcBlJii3nYvkWX8xIxhC4Qpm7d8DkeIt0T20mh
5bnp/CG6O9J4IbLWIxd7gvem2IOb9OHzoBPAeevrRLl2x9H5+wPVmSQeoXONLy9l
9jCbnjzbqxPQc/rS7u+vE7Q8xq8jGAESkNRKHpxwUzEEQ2E8yOSf/9rQEBE2ExJw
rFjVUqBEMCA9aRmU7ECMtXC8yO7z7+H6/UUN4r7+/VZHHhHy27OPBrFou+kw952A
HCTz40lRsKuEm9tF/Wpigs7rcG1+QH/DiF4SSzqmosm0Yl5Zbin2Y97eGVaVdOSh
X4KDW+iuSdZFWFrq6TlRs9rVWdIlnnDMnzj4P+Te91ySX08nEA2y8TvpVeurjRtZ
QioMmfHMUaAJzk/fpdDLD8EjeSEKK3jUJKOf6gHXXS2usX/hTjnr0/Zmt6mLyZMd
JPStYeX81WEChIy8qYF/IYWPoRgENFwk1yl+af+HxFz8QV8jy7wpGgYdR8fL6Kjg
YbBTvZtCCROlwX6QNqGxEb7uB1XTahEiUf2us6zXCeRwX8LpiWuppnz+Kndx1KGG
oGuUy05o4h5+G7lOp5Z/4mMvm19ZqzMq/fc0Dq6uu7C4be/4xhBRxc8/BO77AMO2
bc10EJ7FkgEUBW/hxo+8vXQQtDVxDx/vGrTijUg4ZmcX/ntFJzWG6yYVRMrX+xvj
/d99mZ9raUJeXQBlXdww0FH/630pQKLXzvv8W4w0hfHQmttMIRNKqdnXw2uG10qG
vo9eHHruQlUye36cpo8Jk+ZlaYmVPCkuB+kGD6nYvqQ2bsr5ZUC0kfhvCZ5c5cmu
I7GoiS3qGI/TIPQW5BPDg6xJ/huI0AL0BnvVGWsdA3b1ZJfD7Y+0cPXu2OToXShY
yZq0hCg4sy3e4sCzdX0CJoX6ptsVqySu1w1AxxF/X5AKu37TAlp/+w64Ug6ncnlQ
bK4Zuo7P5j39PTTGrt3ppxC43zlJg0kuvR00QqCEBrZxlf3ihxDWc6CoDDfovCS9
dwuc1cYxR9f0V8est3vdvv07ONMTNpIEgX1H5+qNlS1HM0hCuERlc4DDNC0fPEhl
pwER9IC2jt+J87kCoK4lzgyd1v/KqEJ8C5WSaHBos7x3ybxEmw/dbR4gSDTGkEMd
e5LoxkeAvalDWxNMJKTZIv/XmV0TxL0PF3p/nmp6a9B6SuIt1aXWhD7Cxjfolp4A
ASIa2QVQB7UiThtHhnRk1ExDvDerWPRgmDQL7ZvYqwVtmNnf1ixuz/89r1wnEHCr
62MurD7K2b45wxzHSuN9MTHaJ0EQmv6X7mQwGTUZbplaq/iS/3/NSjKNzQkRFqf1
T+UzSNEbgkUHa7npAf3Ov4MkvkBbRxX7aomFDzr8X/9UsQ90/bGGEI0KrfDrgqfk
uMQH/3WNbq1D63IBmSVJw0wsDxbYd4dv7L0tvWZybnw4l9vHmbT3rE5R5qW843Mq
9BKNN0mPiMaKUoGuw9Ktmy4oOfyO+F6//Ib/kJxnjoSUXxBUHm1tW3VfXpX38UoB
mXR8krvD6KroJWVqIYLdZX9herMKYMyWFA5ksetgGgPmfvPReGVnS/hLWUIit+0n
ky9BD+aCPX7YZCCzkd70hGT4AJThtW4PD5Y5cKfyXA7l4JNwEOVaq9LQEji23tsn
I0k57yYaxyHZIqPRqpkot6GL908CAQO1cT1BnilxNNTOA30+ulIrUlKSjfo1ljka
Qczs9MCvn0KREK9b9isDI31VRZ8sjaR7fBVqLkHvqYcMkgy7ike/uwfofVJTBxwS
bvNU7SyHuEjhn1RFG7fQeZSNnQcK4V18DYFd/2XWJZjcfGDzu1kRr9936Am7z0f9
kklmxBUN0Q0ZQLWymBoqI9rHyX03OYZqoQsnaC49yU6igplj+se4qx+Xq0tzhtwW
KkmL+ntK4mzKcW04RTHmSpWLH12CnutKGWc0FE6Pz4NwEWWJqWTOWjgLfCImTOLp
eyk0e5cz9CfuGsYWr2g8jl/gR4p1YEZ16PZqajpFmUrmm2gar+87NsRemZU1FkyL
VfyAtdP3kVhwmdf+3iZTBo1AaXHPi860J5+TSGd6wMkgI2oXbdWVP5mQdQgeYZLv
XqXEmEE74mMkdq2iBtSuH1k3Dm1uwp7saMTBo45p3WYb2My7uJQ4yAeuDBE/7aiC
muxFxcXcbOBoGKfx4rZOgS4C8NRMkDzXZ2waeytKa4jImq5rNn10Le5mIfOZmaMj
JF+grbmbHh6KCT51RZutVKKzIkEz5g0hnS0SseyLTCHSamDRFOAIZsD4PdPx1XrL
irxlgGIqlJW75v9OQG1y/yIKDr8fu6VoExktt72xcwJwf5UqoIS955HFvhD2GTJc
4xROK4S+EN8/wwVNIRjzu2al40HMG6Q0ZltPwTp/9wqmTJVrP3+VBpHkXg30nMtB
id1VxnRlt3kg26IdigEkmqJUNr81n5fhuZdgKF6dGbAm3rsqemxCmttVG9NcZRi5
GmAwvfI8jXwBpXTfwdoZmPMlfxCp8zaCkrxSOgCmrBvOUngROxcmH4BNVQW4mUI1
NXCtcTskC9g9AoHFl13Kp/YrgGrJRusu8C1Uieushb92tBYV18TBNH5ALf3X1+D4
dCowwPrzYvWjpSbDKhzR4MLFV1ejSbFu3GrvIrKOW2H2Hpc55dD9Rwy5pVoYJQkN
Mh+aMDbQ2QkA/9Yy94CVdhX6TVV23A0y0eh7BPZ0Z27wN1GziUb2rXhACZxwqKrG
aDDNvvZCc68AmTJ29Umjmpok4xFG0PrpuhWCq6iptWE8EZHpgmcFOmNdlphW2DOC
zSvB7Uuqr5Fqa6+F7d+z4b7kwpLZl4B1aPgEq9tc2QccOwjwhzfWKK8mZoOqZE85
7Cv73BxRPWXzqw4AWOsrGv+XvqLSOEMGi+P/EHtYur8ZZl8jrH05fo7Pgs6QCUSz
4sVu/b3A5cav5NE8qiIYsneVYNk2AFYkeqK8EjINno2nvMoM/RCdNZFJt/wrgbeD
hPzSxhJYn0sqd4xsQ9n1JCir/60n6+u5iQ/B1d3aYmJZEUWcN2wkVX3dFuOW8pWZ
Vlcck0Buk6aR/2NoUWnGtgzm5hKLP5pdxkRM5FsuAMMCs+2flOED3UoDywdIC2d6
p3CLHvV1XKGYTtzptCQ/B+dR3JN+AC+zwcDYbwaTL6eK3WIYiHdn8QX22yiO+U3I
uUHBIrgt7d/giNXMXC5jNxQHm4/LbOdPoQjKU8f49wuCkIf9DvHctfgVb56sy6Fm
nkbtMWAkUizzeSpDhacOze1g5n6yzcsCJKKQNUmG/qBV7ppUXWkdJE5SLZem9yTM
AP59HKYPP7sFvmKPqO17GZrEa/p+0rukS6WurQE5DuABzhXphOw0xkvQL27nQZYu
X1Ru3ydXKWWu8T+Ulz1Br5NHscybUu+0MRg9TQAf7bnflyqtiot4/AMdLHU7Qgzk
CJtbRbPQrMUdcDNoWoygvm4MdzWPak3wGItb+gUdJ4ka4yDvrV3tQvnqpht8tQtl
N+XR+rOom03A6uy6WRM9Phfz4NZoEHXV+0HeMs8VCMlm7Y2Lm5KUHYAvC5rh5pmE
16Al5vugIjhv1JRGjWujgOA3wuvlkmyDN7KGlrppAxY05jx/C2KkxqLG6Na4cekL
NCMHoYC7nb0E+17af5ynWyVvfzSxaF06bUW6fQa6YQUEzrIV0iNwflO6hmOKAGGl
Q2tHCSQvgJvx/ZBhzVQJUPwLmLTu1Uzt2mHOq0scK+TVODwTeQFDuq+Atukt3iuz
yvIjc9UU7urpp1EVVb+Zl/O7dpcO7U3YzNY9Tb2377BnedaB/4MBAfgTVlFvEOfI
wCMNBPAhwZG00aXz612JXXU3mbdqpF9BSheU7J23qEuzijWCwqaUiembNmwmESx4
EkENfUOdFkUQon5AfxxCx31gjNKvaGON81VKl7X5wHjfAxoJFm06zi+E2N74bqPP
fu371h7hg2m5SNsLSWrkI6cJa0Kkgs/sEIBuQBucBYtjkRji18Se2Wc/oBL/aNtf
kv5eCFr99JBh+4j3lD5XJT3qUMibW4beCcHhNFsBq4U6bvbShJE9lczA/U8gya3O
bl5Lwi72ODtT+++SbeYdBL0te/N4ofgOyNhKbbuoKDGzMWNAR7GJp0l7RmOi2yNR
Td6Shk6glRK+xTQWhwbswBQupoz1Rw0NfBoJCd4NTSNYuhyvw8HurKdPWOaWVhnb
cvH8UkFVt7fQRldcsa8fGa/GkN9H2To5fkLyoXAGvdqPZIIu6Of0s/YChPPveni/
s3wtcdbjfPs0xsVkzpHtp5PS07r2gcfF8tR/y+DeajK4FVZmQ1EWTXDPNMzfGrEC
MchPvx3f66qp4l1GFeoBO+4/ofbiL1pt4sDcVw6YHj0f6E9VatgOowmbhU+1ZC/g
/+umO9y0f9RKe4WleBF/tqu5F4b0fz7AeAIfvGFaAa43w21SNkXYbGyDtrMr9p2o
317rrHJOx72/wgjo3zPFUlqlPDrxKPSOZEbIfy2YQJCIFvZEyFfLv7aMwdBfNp+d
hy+6qfZWck0py80SWGkrzPHn7OpAXgQs7X3JdhQ44rwatDDYEFHO1GfpUPOSvyEp
XgbB/EAjIdvcITvDNSNuXXWoKpUnhlJfazHwh2QLay5AALbT8pi9/tyNOyCfDOLM
JqZAPe1infWWoSNDv7CYtTtta12FkQq67ZWSnhExl2kVue55aUfIYLCgssjQapN3
rKkXSDjmu4ZnbeoYsWVpypX7wS7+dN2MnJh8Qqdmpvw3KmIRZj/xPV++RPDv6rWi
MAi/LJ486ZEXN6jqHoXIgDd3PxMhdwdCkpvWiUE+/mnCZIA+AepcD7XwplaNrk+c
6YMmwRSvDXpGHZW/vv43FcrQ1BdtERz8jcYPuXqRMsVcvEPrJyCzn54m95KGcda+
2qSr5h0/RmfPDxyxAr3YOccCabRsnfdoFFNWZHH648gRXj5FudsUW30q3OX0TokG
bftjVLaPPJJ6zRtd5s/oa8AhKtQPKXUGvEviL1Q5zJwwMMdUBSF4pdsuntRvYYgn
KoCsP+1M8QHsBQwYKKExCJFW5hMusDpCq9sqjMzGH5ihtJnVLtt4gxP+icjx7L6/
vryjhKv9Qzfc+m21TegqaH4Vj7qYz3kFyO0Tg40/ZsVyrTEWaY3rlz/BTJL8XcpM
mmI+y2S+NtRQRgaZ8DZChZIKUssu588+EMIwmKKs4ioVRra9KlAGE6LgHhv/+OEq
4aZ5na5Cl9F85Kln3f3JIKSblsJFlQMtgkQAcbSdMfL/iO9Pxqovk16iE8H40RUR
5KsRYBkT3athHSOfumSFQa/cAS1yTastDFgO3fbTv7GGElQ5Dso9KCvK1emoY1z9
IvBXXSD/QkdLKKmO00Yn5W7zZX0rRNy97E2bXoW9QLwUfCLYMSBzkqkFNGseIW44
EurCwx+A1qpwy0x8xLgObmLkM6F4bwekvUdTjo/DQ4K4uxwAztNmWsOUiUQf59Bc
0V0ZQCZi/A/WMUAMYeGWnY4XqvOhMObHUXxK7RBd0qu7qmAcIuejrotrkJCUGP1R
9csk36qrsUne3ahN3gxyW3ZwPAaT0sopwAyCGrow+CdLSP8gkoXuDgltOsXOYtTN
0L1PmJlWq+Vhb3vo4D1GgY5JVVvzaK9sL/9PId7ScK0hClWx5BUgLTb9WzzxjTJq
vjIh0LoB0nQ1rmBOciGxyrLFSNQEXjIXYpYv+90D4XLxcZXbWdJ4aXNcgW+LeNhj
w/LuTJhbIUMOJWKrEKj+EtdRmYE7TV0pO+SAgk+7Wju+HuPCm+7egVfsloPxJr71
gVztEvOIpM9m9u8AxBaWDIkBcG1akN1jI52E51k4wcfnrSG7wU27Fmnh+mwgAr08
4EYGFo7Quoe5jS6Mi7NuWvh20gsTlTCtFpFPVbBfqeyvpYj229JlGq7NVtg2Tl8O
vUgGFFpSR0gllb+ci3NZc45E2r63t2ZUqkRIkPEGkNXfFKFZzQIkU+wexkzYxL9q
BWKedSbjheNrepUi/emadNqr8wTXujBykATVfZmRvTU6L5KysbVKoPWZB09NaId4
Kbhgg/DD63TS7vnAFBHs4pRrK6aSQ0F4/Bki9SbYnPJqcAOHHpMXmWCcxuEFwMn8
0D338Hdz98fwFzQj2GYvZux09ayzGeaIujPgGi0yg9Ck+9tjxcCrq7RVh22S5gxi
xzL7wSmWCMkqw0jo9njLGtuwg1wntR9bFXM8HIwB14R82q7cE1XK7UR6txJt3SnR
ILY9+9aUfI0hGdOBXrmBwDf6pbj+fnSlaElqpGk74rvuG3Hxrd4GjaQlXoHGNDuT
FvuOiMSGsLFJA0fQR7Mpm3aEUYXXFHwspOTw/g7wbxMOFgWhfqgexdifwZFlHXGG
tRujjgxIWnjNj/vMsVrY+Pok6kuKjzZ0KzRCcwBhZ+3r+zPxOAX9GDT2KLrpU2bY
acA34r5xzW1Jj9pkgkVQ73WG2V29SVCi558ZDroy4oHhTgavMZk5Y7K1E0tOVoHX
1ucCGj8QbfhddfXx/UyDSORMDvzcBExLNDsBKOpd1lye63g+v/fYtgIiJoMJgfXB
fDenNBOTgDIXWNSdT6iYBS59svvyatr9Wago+PS5dqno3O5IIoOgHUD6TrTW9CPi
WzKC0wxg1KkqWesPyzV82oGSE+zBUjZuDim1QrABRv3t1ZiXSH1Mk1r246f+XRsD
aqt4MOeiygkzr/AyOLpX1xKdIhAd4PBRQ4AUn51o+A5M+mNeo6yb38xHMU1/HU4K
y6tmOmqMOiwTv2HfBezuQGSAqa3NIQsD7V8UAaDWOXt8itd8bKC+xdGbooKTRztl
zQjxtmAKtyc7HF3ue0vf5ecLxfbKzKqqkCDwdRxlaxwM7EW9MiqW4A/RAVuMmuHy
ko+m+Dcx1/qjhm8G3Swo1u7708qiSMqPJouloy8m1pQtyApbwhFLSTYOkwmWhgpQ
e/ZjdhsF0QhatbMy1dfQ5aOSencTFfZwueu07c5tip0CY1AKzDyggsQVXOEuVIQD
fOYU3WVALJX/ed3uQqPgdJgAdLz2J3l7gF2b7PjfLp/+WiUU7S1LBDlIppdIn3jq
TfeATTVMM8eNUemDsA/Pyj7K+Zjsr861yVRBA8WLvatv7myiJ3K+eBjEoh8HgQfn
yTLkt904KOdT4r4u9C4nkjmLYklGkIAOXvs62QPf6emlHuKxJ0BWmie3dN6ERiao
nna9jiRd1PG8PvSx8MU0/B2IncyNGvMwQxv1ij0481v0qvyrO1dIrmIzuXOBSVVa
cMtCRuuZF+p2Bxx4t4iVgd8gXpL261BL5B15U3kGNzkhFAEk8NYFsKtqULiciBe+
PE8M2pZe2o3ActEc7FZx5shT6kriL+pkNdtS82n6SpRqYESnKtsnPni8YtXPFTLw
bM0jedBwmntXEetB0VjqRQSvb/9tNDhRs0FgALXbgkbsTq+Ue8Yts7I+Ruf+DuUy
14JgZsSBM/fNg691oMCx2+RVe1ErgSJc2CCfn8avmQWrQfeeQgIvx92PIkyg7Rj5
FuvxaT2Lh2OhcCYgQhxPVbUcsq7vW7+KWM2RO6KjHVCsE3REQXUNu2v5kgvFQf18
Db6RIU5S+4Ez6sA1dRpcmk60H/sqintgLsXNej5s84VV+k3PIhFJudIdamwNZNvR
DCUnifrCEsNSR5zDx8f3UyA7Au9bTG5PmIeo7zhpM4nPe8FZCDDJlmXQQr6V9bwo
6JqkOxSbxnShJ3oIG68Hk6JUwd5ul9zqqSKhmUFlRx6yZ0KZvid882UuDGvSwF9Q
kRnbmcVF8arDCqbrauFKQoqd1YLjsd9FBwYvZAGk8/bkDsLAvwziE83oWMAmH0UD
ck98wZalFmV6e/gw8qd0uwDlYve8eM9VMLGaTZ56konoXxIvAOA2ifq667RBuHh5
L2G0EgDCqUa0VS0RV/A7WXMSbrSQcr6d3etE6f+IDsOK6Pnl9LmjUkWYM6j6ccA/
eKolBr0SowXbP+GKIS2RqCdtSzEgU5ZZ7c3nxYXTNWgIjdtqG/W9XMv8Ex+aSezc
AO94NE1P453X9JWtsS+U27eyUceeU/ApMJBGxRak35NIWUeXbXxZOz0tkKku5Cg4
zYMWqmLNbPLzeqeR5U9Y+IwafKAcLpQJ3w9fTUsikdmbW1G9/ALSZdfQr7SPDlIK
F6DdPoY6iXGB2oN0+9/2+mnKAHYXai7bqa/9vHhCpG6oUykM/SYVfVNvAQDCkQOW
oPuULq3xOY2VuHI97Na3CnaQ6E9CwgfeTBuJhhcM2e7B2lNZmqVJqv8yicKbaoHs
aZ1n1dzjN6M8nDQ1saWBWqA3UFhb0hzcojJgbgnOIgE=
`pragma protect end_protected

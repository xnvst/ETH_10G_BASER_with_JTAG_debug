// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:23 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RFkKD6SfSiC+oC5LJRBla2Ucjouz7D1fh9v/KFb1jnmtNmgSCOprwc5CdMuSS51R
LZcGUvz7npXr7RtYSaIwJbA3K5Oa7F2MvqOQnSedTtVqDVdx7NwR1ozNX1ojlObZ
bQBdjlPsu1GVCYBGJqleUVl9YBloOaq2wOO4RYBGhgc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8560)
6o9aeP3R2z3m66NQ76tzREJ++wK8c7noPG6wxnBCIuOdiIUODbS5gyNsgrW1Dwc8
J3qXnd+b8EiS6pYGMkfS/Awa+E7bFpV7dRus2fEFHNroB5fNRdxDWQKVywtaa/X0
1swSxe3b/Uxi4xTU2kn/rdflA9ZbYpEMde8u0vKyCyo/EGyGATBULHj06KMMt2BR
TRFftsIirqTvLkT1N/Ex/WSufSDMPBCEhTytmiUMSPxUEcSlgiOTLrzcJWx4iuE7
3pu/qVP4xjiFwmwXwV7cfkeKU8LS72rtHW/4TjE7YaCNUV4PIVWSFpevwzyBNgtS
Oi038WByaM9zjCqBkmsKq3sdhHxqaDOJf73KSAosDTnbB5uLLCq0UOAcc3wlem7K
Z290OWkG785KcCi0mcV9mf7rkT9HQ0POohmoGBnsYiVScwtHPuP7u3aAfQvKP79g
ICye5lg4Hto3cBSyhNYkDf3B7ppVlf+oqg0DFoZSu7VT/3AAkJodO5OPEy3WA9K3
v3tNr7D8LA0hr2nKMrH8azqtIuIZLEl10fQBa2MqWz/WNHiRafnx+sQ+mapjgmUn
UH6RVRgt02c/mXmxO54yFBIOMTvsvfGPFEyTc55vBw0XdPhxLnCu6ZAE9mWy7Ej4
JReNVQt3JSjil5LBxzzQbEz3aCWXlHCf/A/zL9fuZKjEjYYYSamGcki2Wy4L/6j9
/GXRxDidhnxDiR2WYrj8XFJU+el4JeUvwe48k+lz7UGdrjoXRM4cd8Fyc6GQiVVc
Ic63z7njsULQ/WSTG3M6cFvy8hlRoYi1H+zeU+VslhX/+imcbNirMuAALdspavG/
k20U/sQv2+dXQEKHt01idGxRvyoN+vXwjirN9ZcYBoZkP9apdw+HQ35XWpipaxpF
XVqXrKHxcZyq4gI14QtkE9uGwjvNxYmEQN2j6XymTy/hluznHsp0wOmjWCnf84Ik
Sdcw3CwZaxUtZdcCS9un0Ilk1xtAxiq5255N0JE6Bt1AiblTK9XhxUr9Y0DQ8DQh
me5iU/r5XCaMCpPum7GOBnsrUgCworfgII2AOcBJX4zKczV/MhMtkKx2DDXjDI0A
3MPrR7xKE/MIL2vWvH7WxPJ8oVFV5+eqahGdCWuNWeBJVxXfm5Dai9mJ1EtkC41F
hceJtifeTIx6A8v30Y8Z9OEHpSv93+S3BHqxv5TPSDKTbVkyDgRDfX3T2++C6xZh
Z7hqhTm2rjnTt53I5NeZI9WY/u6/JZg7kbCulET99LtZVaNtjunLe7nxMfpIWlFT
6E0K2+l6gtNaNYWQ9IgTgyUTCnCNlb5FwFTmV+GE9oUOjxmJTr1QhWD5U7EOctZs
JSvmWQoBkfgeylo8q9Yf37+cmMGNEgfuIrKfMBLz8/3HOWQLSKw8qYeFnN4wj408
NhxKjvreI6iKm8zZc6eLgBFmYnhfeABeYO1RxphO5JX0V56ubfdA4wHahYtYX+8p
rK0aH05OAZdBV7/Df4d4PBnlR6SCOXyN4DXIwKByO3UY2D5k8PXqJ8NP/fVXThjj
oDS07d/QWA3GdkQGqxRnx4k9bGfD6WjKNH5XFrhGVLMYCb8Kz4NxOyxpr/HrdQ3a
fLAdliusIdRDP6DD7LSdQGYxLQof8cr4CY7vzrdZTBCxsKGiK+SFluQMm/zvgnqu
1p4+FfCM0z+kYpaJeIWaKdZZlytg2VhosFgwByrYHONV6QiM55SYEg8lAaunkbWU
Kbu0UDMhb1CCz0se/bwWVa5JvM/4Het5VfGJu0ZtiEcMHV0Cb8YyUAzKOntyeJWB
SwlnvQW4znMyxqG+RJsnvn05dLt2Qjy2uxRnIRWwi7L/2GEkd96loHR8SjBfEUj7
zJiV3vSc2Gxzs7N8ZmtbPweMF6q3rvjogfRvnJ8sr6y2jrjZnc2tMuIUsyzl9bj1
hyP6krCJXV/2FgfhG3RdFCJn10b3hfC8nyODOVs337zqDsbhcipwpn9tHD9BAgJT
9EeqFB5UTHM7jGe3atzVXZDpBrZZIFxjOdTHGksk+GhhKq2LTFW713WKl9MLoUeY
2t8iEBSYUxv33BBFYwbR/MgFXj0WNGfXuzknqoMTTCPBt5fglDRaLfyVTRWh78L6
XOxD2jSUjzytazg0WhOL071iDZvk5XcnhK1jeqs6Fipy/YZA7u4tyvyELcDXbe77
QCi7N+RllQkwdBNkVZqE+y62xfUTIDrJGaPoLScDhxVfR5+ps/yfUK9lhx3ae3Mz
KWKKKxe+p/72lbD2Cqdt8cCsBFZkYxwHn1ldBqiIfzufW/hRmLGI4UxmeasYlpRQ
vIzOYZbiLV5O6fcHHZYP9Whm2gMYhNMOBJ5E8WxRuwE0/4noJ9rs0a81G8lRqFc/
qc7K28RT+wZTGGatTcUynwysp++eezkDOI5UQ77oXdQbJs1BvmU1lMuyjqJkr2/X
JzHfPNm/La5d3SQD020kOudY76UEjvr4eFoQLYOEP1yJX4PpBSJ4oOnXegN1siGV
p1GiXc3Eh6m7EnVY7mLCXJv4U+WMMLZe4e1KJWhI0RTeSfu1xiQjWnAHiCCFACJX
epJqJNOCL2JFTujQpPrStXj0O8kT1TPdHIDN8gJEzsxQYmT5jI15Gk8du3/6//39
iysp6AzJ8JLymJWtmDzmhrqKzYp/4EGqs0vkkRJ1dZfj8yUTOoWIySQqcWxP3VIw
i7H74QDDEQw1J++RpGML2gtfKf//PgBQB0oFC7QiNtLTuG4d5App8Egy6Egi34V8
ujNUd4Aspa9D9IFNkCz1DGtJBoypa5dUOtLxpBE5IY+rkpYCwbbg0PokBY/mTOKD
bUcdUxFjwIbr1p58y0Xo1HukpWSsubaGcAICjcK7xY7/BiecnAgDxvkvGE2ehnN6
IJRv9c4hPIwTEgJtcSrwdU8O90+6u1ti+OiY7gDwe3hCg8iYN0Mdm1BLutFP5UkW
BBDn+V79dSrdOh6H1GyHVv7KMeVAbbzM7NKfgJciwjobdCn2hMQGtIfPv7cQgGgC
zUo1fGtzt3RXsBTwSTrQDwztWsE9QYZTc4QIzI/sdAkMKLRUlG3Hyi3fgbq+8usl
ZLYTWHh2Wj7KtSFN6GeC/KhqpN+YzyABjOavgs4aVV+xTEO25557SmdAX4S9f6wc
AkQeN5H5Ip9BUKjTEt8e+9OUxeVPbs3punavp6iOdoxk5AZnFaMvFnp/7wLmDXKE
iyYMk4i4/IiPtb1gN9vjWo5jzP6PWaYPbDFeUmBEbuuEzBHX9tdli+5WO15pOBQ+
T0pACNXxqqEETr/kjLNedo6tON8nyPYSM2icRNNTkq7TJ0ZxX9MFmPqxFHXd1tqc
gImoHEZGi1+h8Dew7ZzAEOllTYKPeDwU4sSDM51KnnAD8NIf5mvGUf0b6p+Bi+FA
HChydCXJzaxfoYTg70wNZoDryT3z63v/850NBA8O5+927UhpvStz/gllOlhmTIRY
gzV+0CP0gmHv97fkDdQP7VqUtGnlLWgNmvnymjxU84e0TzN5nmqGjRal5pW0AE/D
yTLkSSMFT4/qEAiG1R1pWyRD4ki9gUfd/6JVUrL5Npqjq9NNJKhxiTVuHqXUFC4R
1Xh1JyYin2RLdGCas9VsjwA7jksMyidXcybfhxnJUswVGXP2PK7ScrxZYAQ7vTn5
QvjP6Bw8viUesvlh4hzT4mqdyuKy2WQ1bvP4Bswds/J+7L9BdRDZ6uE/xfdRuIKs
1RGYMTovJPBdKSfkqMnky4OtJcipzq+XWihrybsmpScZ7LinQGBYCEUDjlf+qxkF
OMK/hQ/XiepQDa0dfnOEVP4XVoELEUj68avdgpLKOYvo787illfgPFnofiHbG9l1
H6JEFfQB0/k4IxD3b78TClyqW5Lh1XNnn3Jx5XVMrUmDwd0Gs5N67NBZ0LJ5WxDJ
7vXIdfhCxzqUZA3pEKpQ59ZVE0PAPVROxhVCZVqaGR+0WY5kGw/M++qA9Ctuwr1Y
gbsVV3OOprnuHxwHc0vScnqpNVHtXbhF2BVsmQ1wRaPJ/byuksMzqf4E8nvVJqpr
ZTRBdh21PYQVFRAiO4x3P+2LUub0aESMSDzAOjTddv5tB/DZ3GxqMw9mwZNNpxXz
7zpUZblfeRnTozp2PYTMdP9/oL/PymX+qwjMOQM82jImIey43TORh4O9l0JV89UW
+hDwAzegK66d7Uz0IutPNuUIgenjqXhzZ8/vZRsw4kNIqKOgfRce7d+tBQSuwq3u
eM4zRbcLAfo94LgCAMdHu+MkCD3843nQaeoXW1Xn7YJeA7iZfl6QMbNF8v+mkzCW
ews1Qr3Gcuj6atMnLdnE179d6tMiTMexoxcvARDDX8j5rl13x6Sdl1FzvCrzZcbH
qcmdc/e94olAMXpoaJqaAajzWFMi+KRpihkE1F0dZa1kUjDUepXNOXqunBh9dzNb
Xf5k7PN14S4JfTNMi7R2xxbh2nliX2iGMMD/eg88hOjBMrL8mAJ2PLwj7Sj6UHT8
5CMv8ZR8sef2wakHGGfXiLFZyYvkfOwqRbERqR72tBMKS+dBF0icBatqXmiQvXyx
o+PZ4JY2Rn6monjvNRk08+vF5QaZkpaQBgUpOs7rgJNBw/XOLOqwLWdJyemmEVWa
zqcTko8pJcFrzzqLX9VRjhEWLmdHJTj08frjswno1VKJVT9bTskVizxEnD1PnGjB
rwmRwL54qD+EeYgYWT6dgmqv7Q93yCDDEg2LZNRzIVpNgtkTlQ4EUjhimhe5o6Tc
/bPM1xGrB8ZtA9+TVt7oJjp5Mydfmn4ID7KbQZvUy9pa3KdSYi+tw5vgHUOh2MMn
0exZm1dBEN0Ga8wM/0ln+x3KXSy/BWeffHJxNTjpJz4F2c7ceUMmFHWd8dgvvszU
q++HUpa05lXHIGasvZgkv+bM1EWRKNzo1N2cpGkMVHRyGovGLFgvSSdnOKyekUqI
ZQi26HRoO1ZQH5+k1D3z6RHvDw+mhxqJjWqU8UEAodSlUm6WlLULtUc8T/Y2Iudi
zBMJC/bGVcfOo8LkQ7lp3l6wU0cSC0nLPAOLYQSjL5ZWYM6RHhbp4ZTVgWNu0AqN
bpgq2P8YJ7P8CGcPm9LGlal8Nil0+zhxLgAh1KuVtATkB3Bjd+KVj/n2kcs+EAJ1
UJpz16TbPcKCLWX3prF/2oJsZOAZgfQom04xoTHXjowO1OF60F9Ulu+klrIA1BBd
hWWucqQF41w+sUxuYQgxux5DJdTuiS3oYxVktxKgwEEb3dAUz91wN1fRUmiGR7mC
fH0q1bqQL9HeEezFaJ6Wdp+1cxo22DY1HadwJlHHE5aZWtnzhn9/HMGUEj9Pb5X+
L1rURqsic5zLP5a/jt2VpHP2DofcJvFWTZ1IH0UqNDpzefwg9feHkfArrBNfgGQM
sU4EmvvPlFE3oUd8hstKT1oqT/oZgmaJA4Oplc1TajiywP1RHbywj/jPuLgxtqzs
lsIeZeO4259Y85J3l4p7VfkPtlhK2Uc4UsXo7tsdAancukNq3QRuosFurFOGMZdO
glMAFHgOntgONySouAqxfugonLoIyqgLL8n4y3NeMaMqI8Pu79XdDjfw5vxGfwJ8
WKaJywcrG4NWMrqJ/lgJiRrZa1qerYt1tcjSFoP6SnrAQYrz58EmcTurTi35NyuB
KERuBuK2hrGM3OIJYbUX4lTl93YfumZxyeKxpqzJ6CLcOAXrAPHZ4cwava+1bcEs
agNPrFjXGem7yEKqUmZAz6XaplzwRS+nK59qQuGYM3jokO2uKDAtU4kwU9lx76Tb
C+8azGdPi2b2K6xe3b4n2ZuXD1tSR7k/NXs6yhQevS8chdFA8gRl/Z/g08IOeUO7
m7pZ/o+7y+UplZbTWxWSQBjuz8TtHSk7nzYVwZAqu/loY/ZcmETL7qPFMXo+ICV9
3xjhQ46Ic5JiVIDBoXDT+ZPrAdeEk7GEYiPXsvurxsxBvYk1FWq/jgwP0xzs+Adt
ktLViBcHD9BTgJiWZeW9aGzGLmX6DsElvgTH3VUXTSXETmKMGB0u84x/tu7O8jac
NA/JKpEIGoNEasdBqdJ6+cfO5hxNs2IqnLk4tXG1Y5T5bdTBNIMFi0elGgDACZQ/
j/WKe/J1RVvjCDGDTvSB72BAIYDhKnfGbTkanFTnpgWOyl1grYBuCpd45DSytLgs
CSykH8eX6m9b/3eXrx2Rr8iTH5mzQE2YE1QyZd3MZ0s4QbyDK7DBlNE+tVw5QPiu
JHw7agD+05oJ9FqNwRMwn6pF6I94jEV8UGbGnEGAT3KpMw0I/GIWWZ3db8ftbcqk
ZZe82D2P0PK4XMElvY2D4gg+EymfZEjdyAtfQObC3LRXBB/lOj8vIsmAMQnG56X3
O/4SpQGLyC65COb+AfuRSuzrM1FkexlXIdV/i08LxeuM7TQKz1wEejtneJHGbLE1
byW73TWgT/BW9O6kTczmFl13cGAccAVXzoRPNnL4PGGdBaiUYBRnWurgbU5e5P46
9jkvG+TzA71vkTYlFPzF8dThNRyAL9sPZca7BlpZlUnjAF1vvBesccG+3iFu1FaQ
xeMwvMr1NDTu+skU1Jh6+zPw1OHPBHTiOF3Ic/3nbwAWv7KHGXBbMiVP8jUa2hnq
MKVEDf0NlTWPJGBAJzsztbbMNjRczUs43TkhE2F0Rsdiwsl51Ft6HkUqd4OnDaRJ
zHVrB5vlQmxTXH1D17uyykw/swkbd7/3f5rA2n3hHxc2NiqY+J5c8Z0Rhbdz70xJ
kt2rTLBAgczMcCRjYOsX7uEOg1n/TaQaM23gOa6g2HrUbDk4ctfuR2uo/VYLZIxg
u7MzaVLG6z4z5+24dy3JZHvTYVRdTn3535GmKm3GuGiRUirCXNhUXHYL+R3QpCId
543rWpImqCeKFQd1MmA4v7WyrqbCIhVa6vV+0kvmjLEx8iUDJAjmXytcGnbayrqZ
5Ob/5qb+pHSpgSVYki/QU/CFbfiJkRa7uZ52lWB0Ud70UF6YZiq628wbxhunQNzU
jQKOjGl0K58Sw/tqi7XOdsOeMjdhI3NrSa9gEaWext5vflxKgeX141LiQlNSu3cZ
r7CunHhNogpU0oh3aI3RCW9zxFmC/L7CxxOuUctjZpK1ZVRnSFgieMLYlvm72Opk
2ar0EG9QaL5pzpHBvrk5vktAqLTeY0PLBa7d/kZRN9vFw6qbyJwmtJLkJp5S5ni1
ohYXdL06iRnal/2Pg5k+63EWQCsKMh7cZHnIfTwOGD4weGvP3btaPJcXHVMcJFsv
071Hw3nD5+HrVp9rsDcJbNnDDdCA4dilB9OXntBB0WE2enL1aGkkRcYMBgg5H105
0siiFDjsqsVXOAwSr9tDwcF08EMw9zzfTjdamixtefpevFM146i5lsc8L97zXdHv
mmwJyO9EQjEThfQIU5+exJWib21Reg7z2AqprPqcn3n5HuApimnDmOOh99/sanAo
zFgrQm/2sMzY3qOEgKOYOvdPM8GW8H2o9Z2aLXrCdWpQfC10EJOAW0SupmtbVLGx
NWOwEqBDn8iRF6MOy5mYvQJgqvmQvKbkckKyxomiBe8qzG5ONwiftmDwoyd/mwJj
XsqxjsXghR8l420nk231E9W/a8RwDGlSN1+tvgfOB5KHUZqCtUWkTIB53wDNpHJ4
0xfsQ3DRGIEnNH8gDSRACnA5miTJbbMkVEo6uXLpHfIEx9XkL6Vga4gfZuNaCc6I
IoXTChd5iZNOaednRFWktqTCOiIeUrKhM36s61nCsLjYiEyF7+q56+vigAZnCU59
77lOU8qkEHdtpOjriRimenopycrcNBJB2aqVhYf1kxaUow6REiJW8ZYSsM7nwbxS
T+pooSW1BhuLqzFi5FY5ViGrfUOtRmP9PPjK6BeZb81WY86UOZ3QrlDR7pqp0Mj/
DL9EU+hNYePzI3mAtgZZyDbRTIUwPWFCqU75LqxCq44GkW/HvEz1mJJW8QHRbHCK
6i0NePMe4fPKa74ox6Q8IoPtb5RPHa1Mbh/28M2xIEQix1v/upHwUAyZDP9rEioM
UkY7i2pobNIVIbXfSk8femOThueRyAFOl4ZGSoM1969/UozruYnGUCqbmYfrqpME
cVz1Dgz8zEdU6FJ1WS+z06yOy9/ZpIR9cQFTtVAIYfRty5TgyWv1tmt3jnxT1DZ/
tgHeEVIJDagNeOKO0QjYwIbkJXqGe2/wZnWqgbISk6SpQOImwDQ7XE12RRhO9U4y
+4BK1gueSF2OWh1/bGw7dM4Q2B2ixki8E5X/C02Sy2D7VjeoLraIyBustL6Qn7Uh
V8JtVxcj7lqoH9dBc3KHPn93fpN/g12R+e3yRYf8OlJUsB7OuRJO5+jIxPYNAu9v
eNvyOMSEE5q5G7sgVv+oF3CZvKJMwTpf3sqkNVQUQIsfSZr1qLbMH+gTeNTeRQxZ
jeYmIRVs5MBzZHVN3cR5izlXzr6Xx0Cxs5VI/bhuLQLiBC66LDMPNVWoAwqK6erd
kzoyjaYAXewU0p7hDatZFxqDDfdPV6q8ccpUBCqp/5qdfZnK8oikOkOliVNP+xWF
YcI+s4r2FmaSZLLqMFEjW0BjTEoEwfJhlkLrMqY1Yl4qpK+ewMiJX1zpKC7REVO5
IMfPKam+HmRA64Xi7cpuqpKaNWf3XMaNRXObGid5Bszyc9LCwEbh+MiH36miQxLm
DXD7K4/xFBd93I3MoNSaf2rV5qdwsUQ5Too/kx9+7OVfWbpmAMFVWGk6KrpfFHgs
Wzckq6jYU6nwMQR9wrC/dVsMVJ/b0hNQFmzQoqXT8hLA6/GRKarylURz6MtebubR
IkaH3kS9POP+Zxoq8FOeEgw4YdkgkI1RPwmj1TucCji2uDwCxBR2zOUDofL3/9f7
1pCcaEOpo7qnwpmak/vWt17wLfaf5aYJfPIAZR+4A86gv0xuQmQQsySqsDpipj/8
qMaOTn6LXR31xpyFRlWu/V5QYT/AtNgbxurvPcyLvaI36A5zg5rLCOx55Xz6ZWel
ZurXc5jsSklg4160MlE8oOgUo3ecmkdgKmjJmCZRB3mitS283hiFepPcttRnDcH2
+A4BbXx522zJGQud6RW64hXg3RI+enT68jzLSy1fxX9f0yJxZ46JvLbT89PnD3jG
C0guuC/8qEufTSCnKm3gDuTQsDVBupHRDXTnYH7mETM4NalfDOx2JKjZxjiGL0gK
3rDIC11/7t4U1QG4Tm+uT4rerK/8IKeDUAhFcYKnmYJbet5veT5u+Nk8h8RehIYD
S71SorHld6HHYFr0k7/G+zdOaf1RdT91Cycu8dUcRpZbcOWUK3Pbzcz3cy1runJq
M8rDCtScfrT5t0ylVrmD4huGNXP5j3kcthHMJdHN4O6jrsbrPwQezL5kVx21vI2u
kg3xuR1jJm97KoBWMpKzYgIS76rfL2V/2LmOz/vMFLqc3HKMdmKaf+9irE9LKHNF
tss6bxEo9d4CLfGJHvu8lm8dNXjs+DiUWZBOYXFGwn7ACvG1RY/AG1uEdSvX+vw+
YXb8goCF7kBeEt4aBHY/P/WWMBGIOKYNwRkbHBG3SXMHl4phOJWO6bGEDaQ9z/aw
ePDPa1N5jhRiPG0ZUmpU0k3D3kfEzIr3vKSLJtKQFjokISn/r5X3rq/wgeybw+xl
dne1M6e6DOEOaRtUm2tI0Tfih37l8YNaVuCoUaMZiGYtWSe1bLrmqOQcxdPpuLX3
eBYfV+7GkFco3GMKa7st6m5SlF1lMbrCKi7T/ZqGvQBsgdPzyYqrqHo0f9CcXG5U
xNcCx019KWGGyHJIdPq0myan/RddsSTjm2VtHyfUvvalYTuvVbZgzP2hQGBWnMaD
6cUETVquxgXgXSH8gqYqQ7qORtYO278Qh1vVnRe4F+BRt7SVFMyQJqCyZLeI+KoR
zD4+xyBIGEuajGJf/S24q/4TgY9fH2IoKBPyiOggD0BmGnfBkhakJOCbV5XdqAtP
GiHuoFV+8X+om4evrt2TthLFh64fXasEYJaCJuYSgSvzXV4h8z7zfWbO+v5CLY+k
cTtXTE/jjcFcY6pbesBkeuTxBjfHBCjFyptslujFE5GMyM44AAX0arEYQ+lI/AlX
8DWQ0VEJodccRK4tFx+2Ao7wWrZOZKOKJdO4Tu8scesDjATa0Cg11R72NvDZ6djL
B+eZd4/y8pdyu9xZ9PQiOunYgtH5H+Y5SXVLu3E06IK46Ms3EIgCgLVoCt9l/fSu
oehs12oUBWyPe0x0scFbvlNOIO22DJLdu6+jtrkE2SVHjO5jIFXl2VGilHdeD3AY
AZc2TCnq7D6oM+sN4IS+wgBwS6Bim6fKj/fYAcUFdwh1MQZUZGwAyF7KS1rigZWq
zlDxC3tszgRjKWn+7huuewdospWZoHRjNGZTdK4gYrci7BvWIhhcIHvWONFnDRM+
UjYD5FkVC0Yi5wUwynP0Mf56DrqhtrYwKllZWuGR2PVlZSsDDNq3DXZ3Ifk5whtx
l1E6BLpLQm79UyvqRAYGaKPaNgn3pGDCzOUa8Bfy3Vexg08QeDOhFRToyxC3Woiu
vK1phSBHd/cZbpWTrS1lF0v2zZAHt7QgeiQ/VwtT9G3Guv2/uV80rVMdupac69eD
9T53SSF2+ARBjlYxTzNTxrBjO6FDfq5MU1BRxEWWsF5y23+8mLk1Ho2fUR6Dmk1L
jOPYC/lOJclkQvpNCXmS0omX8Al4M4zJOEKuuwTi0KnXvIOBzLrs7WYXi/tkODYw
7DVp3z5FOauboTCZvVKVR2k4dcWc1H2lpTGAZWzlPNBoSeEf58K2V/jv02zavne4
dlBwo4BEMrBzUX2F3l5wjXT8hM0l8JvH9D9FDVh92+XrQf9IkAgo6kVeiHE1UmPv
wsP3IzhccUgFcGkD8P75cH4hvsQi/ZfCnPDoQOSqdYPscv7QcxLTmYa5VKqZbgWG
iJaqr7JeE2n1/OgfSA8H9OFMsCbd1KXIINTDszUPJvQ+aHHDd8q0mW1069TX5BDd
SCMxpRqQJ2r693eUMxXui6U1QsNmPCulM2/a0m6+01sKHXeahLFqqZEXKO5bK3C8
TlOl1I4WM4dn22XfPJb+VKFL0TGg5dqVYafWBDjFdVSw5hpkYVgijuXGRrWDT4nb
ETHNzo0dblhhDTlqo8lEihSw0N1jcxYsz7p+5X6eI6qlC8nZIOH1VYfZ5PEupTJC
LOlBfHPNEk/co00SknIROwJ9AvxzmGapX2gRBiydC87p7nEdM0BCeHJ71XpdI+0B
bd8PUUdN9a8AgIUfdJJAdLh6RknEK5VZVkNQckrM1P5RnFPo/Zd4YwYaYNuUCHE5
vs9LOfMB7Jaxi0kygQ/q3otFFD385VXn22mTaPJMW3b4pRy5d2Xd0y3KcjaY/N5O
79vtZzjF9BXsxF74Hlbby4oL7qQa7fpfIiedFiGh9LdVd07roYi7XdMJ2vRjlahB
cKQff3mE2AdgFndMWjDs/w==
`pragma protect end_protected

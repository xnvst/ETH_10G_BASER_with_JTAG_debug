// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:14:31 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BnvNWr0ofvG5oWyAheh9kyy2NseOM7EVpAkuk504nyCHyNPrjopBzB4QayoQ3/aM
40QPxvQB6MPEEAIqi7gfstbByg6mAWT6EjydiXoh9vd1CJ6EqVHv1nIFf8ZK+Cf0
Nph6+pNoSRMklqXdVUlk7tcknR7zWGdHn4h0u+XAqXM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20080)
pTKXE7yHoMga8UyqXZMjnuynRXsUJcbFXU1LYCtmrt4M98icmH4LVd9Jg60hXql/
zM7dZaU6Rv+WqrV6JVb206ylgZk2mHgY9DgpV3KxTyB7GwC8taEWG4wRz2X+o1cE
y6p2V4AUlDYNwxdKWbPv2s8RZ7OiXwSaH/0R+nqzsPa//1ouPIr41YkEP78hJicq
s+XReQnnF33MyJkm0gqboYAEaVxDZXCmHAuaIX1bAJcU6Uh0V14l8/x3mFWhP7xo
DOGMKwAj0NlHEwEE1amoSgy5VLIuwcCReuSgEtXlW8Du72RwGtBQj6DgYM/CzFzA
Ub/xTEnicR/WpLkZIxIAkm8afEQszjcL7OYczWeE4MaUlJFBSZPAaCGSDFccw03D
AYarRg8/KGdsZQq+5gf6AJ2Q3WcYyKsTZrRAkECc1bpqfznQ7IoVG1t4BD7SwfQE
oqLSVpF6uDfh3dDDRwoUW5RyY+tvw5UBq/VnLX5Y4QbXsAqXP0e/1pgsTwaXE/BE
6Rnlu4KcA/1icgz9jEO8T1z/J3JT6HV60uQ9DJ2Qiz8nuIrCuinzB1GfoihXuFRl
hkpi9MAQygh5Tfn0P2eoJqO4v4OpYHioLQEBOPGwyn/BYw4bkn3VCVLasnEVXn2V
WrK0gGooVWZ9PgNVKAoVA0D/Far38bqWF9JOc8KhAptRaoKm8VGrQpZko/QBIJO+
SA27okFKj1G22P90+mih0NMEiSfuuElRQ+TPd7LaMZe+eQ49tDAle5MPgP7FvSFf
2kKE4pK2F5DSaG/IqcNx4EVZ5hCm3TIQprRa3lAsTT5OLLFRl8qe8eEMNiDwgDiO
ZyENTd1HfQSd8iYuWu4SOsgCEnHgzmPqvfkzU+gJX3bBwNf/4TnTiaWNLwcAH0U+
HCEE8RltjUnABA6LzppItamC4jRmVF/7EMtiowbe/omPMNpd2yxVakpKRRiQ993f
R+ZQMnTwTFtspDQ4z7YU8yqyAPSjKKNj+7bMFsJI/ObJDRkPZpe0W31SvhumrbKS
obRHjjkRR0FxrgBpaCnmEF6SyHTu2SxI3TlA5osy9ywZFpvZukuR+z5JbWPWvZA8
206z50mf2m+KaaJzDoTzhFRGVVhLH7WZ3y47np971w1cAxRd6/n/6SV4eLtkQXGA
Uqtn2lXugHdfiUBTtF0G+gPn0mdYgdy0+fbMOMMd0k09onT2w3ZBlKkduIc37bKl
e33TR7Lu3xnJl4BraRHgB3aoejLCvjOulyXo1WgWk0AdNmvZ+5UhnqbPZ24TnxBw
PRJrr7euVhfPY/0seIAg6CzfYcCGdSKaoYvknptD3vgaTTTNLXnX4ljixTisrnEs
oCQJAThajLbpXhilLn4Jlt7R5ABYRhkAl4oeWzsPcuJacPKDlh9R4olHwLAp+wV/
s9NtJUJlivQNvB2PNVuJDqvhV07GP73jaK6/NVOeiDxpdw2pc/31QTUPDZuJhYFQ
H1whjZkBFOQCT9q4ISwHICE38meaoQZeKcoFexihJ92PPjpyygQ7VeTwLS7Qbh3g
QDZC6OedDYO+N6DqHcYHdc+xaWSZvWMZFkYOP0dhg0BMa8HI/ClxFEssRrXHtre1
y2ME75AgdBCxjUnc++ZkQwziWd/LxjHRPSwi9vc6z10vpFVYkT6/hKvPOj2ntHYf
7q7fFh0YprRYYjONCSOMFSvauVxCJ5pJMNzE/17jPHzNKuBJsYL+DweunNARvioD
5wQaywBfsdDqbmTOVQsG/QT5kdUkYOrAeJDOqTvBfU5l+IEdGR3uokp3JvSlNns0
V9hVWS59AJ7FzHpLoJIAS++Ken0KSykZ8WQ1aFKLmb6QtGvszz4DthkA9/Y86sMg
VgOEuDw4QeKnWHiHUFIQvJ2tn7a7DGNeGaxPfV6nHI1gw5H37JGYGnjxeQiDEaxd
3UE39TTktpuCZ9rp1IvEBTvXnvxbJ6mCtfbMKkKGc19gWJGNZG2EsUx0AkAxNE0/
214vPuBSl5F4kZNEfPKo6L3++mfbPuH3CzFp27HCGQhK3v++m++4iB5VpsvLaBBf
O4YFvbtD1+VJkVgEgwRzJLEG7NybdyZtgVg3hwfrYdNxzGVT6G1FWErLfFzZ22X2
bwIKGMbFFjr07Q+bwoYRQIqEVGfFklyoYmmqX1eulCEzNxcgVllaR65ULhD4APD2
Kb2kv4IESFAXrgdCTME2FYXh2WvTSi/wAbfBCvdlgInrI3q2sComn94j5CJwbnNr
dflQ2eqzqaCOKmSbiaXjFqlsxuJAdJ7US/gvMGqeGGTgHMgbNzMH3NJcZjX4QyFY
9UyqCLXh3/hcG++b8udjKYuHavbhloIyQSXCvhENrgyNDigqVfVt6mtBkj3+79le
PcjpUgBGKUy+ryQpqw4Z13cjm7wju7HX81vuLHq9lgFvsG2BlPUyl3wuw4TcC91P
ElBJA580AkKaISFSmK+Jgm4FsR+iL33vTLgw1l5vS1BUfjT3G/MrRu0mrSxqs8I2
c0mASDyDj6ZJUVO6C3fNw4ksws0Abpt8Cf6qFLsA1AzUjFnSdOs98Fw2PZWDxp/y
0Oga3SYWVw50sB1x6oqnbOoUk2h5dwjbwtOms6onjb5XQfsMYTDbryUfQNufvJwF
ei4Mpx9IUlvS1QRGAlYavh5uODgRAD4UC/Rvmq1lePb7v8hXFs05saM6CFtWMe+E
ChytwSjH0eUFV0hHVycNpWIMECL33J9q9gqNRjQOB3H+tB5/WVFfTbGKYANlWSX4
9Tia84eEaKkzhgE9P+wpvW3ULIKh/Nnbl4e18o3awk9Tx6U3W6zA1sGyxgYH4WJs
MrjkWlQHETSv88bP2pr8kgpC4qkKVSmV/JVLxlhTeihopvnXa+sJN18ixfYNOTDC
6WfKCbCDA8f0oabua/Af1jHOeApH63j14dS4zTkoZOicouSeMN/412Usbreq5P6V
e/MqRoQU/ZqDWrL3iuw18Eq4k2ejdZr3OnOuRfiwyCim2D/LgDf2gr9yI7tpt+Je
q8Z2rDQbeRwPv4YNd+cV1ua4szMxCMkGeedXmwTGIM9irL0XffGQ3jhBAxkjDPwe
Pn2WBPGm1N6Fw57hDMcT1SDVJsSpPNx7RuzbfRGdoFJLy8MjgCiYBs1u1Zbak55M
krSckzA9xM3Yu1BU8ERIb16KEVdANqk4uohr+6Xy/b0gftA2K9KayZ5WRh3XGYLI
5I7fJyMNegb/IGrrihHpsXVx8lKE0kL9Wh743gi8OsdM4b6EzSd+AJTbc8rwaGil
Vu/KzMW4auLr/f4ZNfyaNX7mznxARV/2WtMLpLx46V2rH0w8azROVgQ0J3XLCZWi
3LmYoKzgsKyo/Zffdd0hREkpQ4oGIjwDoIt5CsDhSON8v+7WH590Z1T4FSKdDhUO
gkbUN0IXTrS/+ka/1G37YXEOYwcp1OzVVGjqYj4MS2JVfNSguvRwthFhNvBSBNmu
wvt28+hbPIk3oyHHw034xqm93ybawtB3hHuMwa5NYCtLkFXPO2XpqvdnmQ20GFAF
424HxXR/DiGiMPnw9W9Yp1VvyzXUeRQ4fTmyg1hrlvTfyCgLjoKUlyZoeMPgiwzr
K4MMhmKKie23GDvWSzIjQY4VlJFPajlDhcKR+byAQ+bz5ydLXtSdO26h9tCNwI1/
HY8+DGV+vCfZ77PfFJgvnxNVv7oMpXvm9bKvSyDHtbMftwcdwBxyeAQKUd2KaJ5x
dnHdbmQwOJ4hJMolFrsgIUOmJPJ/MMysDPJ/oFafQPS4zty4hmQAfuz8DBQE+qxq
Kvr9o+nuagl99waXot05TsvJllhj58Vv6q83nyueJzWSSOQYJoM1IH6oueJfupvY
O0KWSx3w66BVlWgmZtxMACCBt4gaD8zr91Uqp0KbflRS1/FTEr1Xs6XTIgPn8GMq
i54vfIUt9MGmEVW4JTa9vO1sIAEOerZb/ldvRRoPO2KUsQOefW97zgYGi7jPJ+Du
4WiotJADDr3r368ZQzNU4duwF4e3DUhc5DrQFDo98um8Gc1PhnmEBVxvRgYPKfNv
X7RqDSyZjlceqZzDr8PlT9e0l7VRfqqOk9AUNe3iCVEBGox6XrdXC8Z4De53kENq
VCAL/ZHKPIxvwULJwyskp0PS7UYSOo/qj4QL+kt8w1ABTRpuVNmzzxqy1KE9bR+4
1f4CLzzcB0D1K4LzWfqMEn5KfBaFkwe0hutPmDqKmV7fv+4fjFAncg/i5mfFksuY
kBw0ILM9EFlhRGf/i9oesvPt/ECuISVuictG+vNee2MUGH/U0/+H4RaqpKIuGENM
PXLAoCWVycjfxObMUK5VtCMfBvQ6L84z38sQ/bh9738CSFNqy06UDVbXoIv2bpWR
AA7hcxfoYZSWaueoidnQG/CDTyO5YNkIzzb2wZ0f+AnZJaeYaupxjQp6zZtOnO/g
yIE+VnK0XXf8+dHxe56hUr/KkjvB6btvDpx0ZfZYnsL1ShSH/S+KtzNpd7/07xiQ
/3XRSMLAEx22OVqRbSn1iLglbdgfxn2hBmwUm60UU4tdYu4JjsNtIOhCZAhWjPdQ
+clAv9x2D74lSRRQAtd4ILVJBSQYbQrDZLYqU5eT6x8+08Xnjirr1W9140Tkcf4b
xy7Lxanzi6TH+OqN5cKQKgMlDc3eVatsQ5rCbs5QGJlfCE8MDktS7mUURCKdiVzN
sZbX1ADGSNB7PszGZQPuuUqAdWJVqxXlq/8UdgAEY93RTJ+TDN+pSgXb//ekEn4v
OKzEJ05bSWIKkwV/plnop7mb1FKDoqyVZXI4t+iyhJAsVgd4qc/ZBEiYe5chrc1i
1rZcfeUYoR2Nk/X3Ezgdgk3zzI1lowliB4U80RH/r99U1xnP9BGAWWHji6OgWi1Z
s2xTHM+S/7+437kWzJPQYOv7lRPmrTTqfke1YBr/Tcly/S4ozPH/nH2rXGw83FRZ
x2CvKD6wFl2qBqoUyvgj/NHy1/+8n8xaG8hICRD514DX50fIq3QjWyTh+z+B0M7B
27s9yljorBbmQMm4jwbVRdW4cyZh+b85qP4wTZcyFFc0uCAoaEfH85WtPijlL3QH
oTMh6gglw4/OzpGBSoG9NZjpsbtd0yxwsTJdruQN2wgTXCL17GF5hYpDXucyERvf
P43UfpUDheOhLGwAFNCdYrQU/L4o2LA3zUWqDeXoI5pUIUvTZ0Z++2uUOKxmRd1y
4TRzED7Bcnxn1H0+ySru5uphqxS+tvOUTNkeBAmwNpfGd+9s+u+xpErX4M8LBuKC
QQNZCL0OH2X4Hi94dH5JnmoEAkPNv/KH9I7uJrJtx31MkqgJJCTkM56BqySAXzHG
KncGzT2obkEkaZtEpuK485+jCL2tuXzi5AFeyMeINzNHtPOkI63ESDim2OO7SmcL
tU3+dnieN0jLN93atZXno2hTA+uzaVGrhtp0fMReMhhsaclKXgmDemhgWCZoDwKd
sWIsD9f83VKDISJr7Qo7n2P9RxhP6joPsT0ZyT0mhxJ22wqTfA5MYd238oYVNhhS
wyUFNrYbggNIa/ar2O4/52Myw42Zf8ywBTTxQAUbXFJdXqI4Y4v1J5ds6vFtXs/l
t/D2825G4mFBr9FcWNgNjvmXya4l7VeG75ok8GTdsaJCcNDcBbu8G3xKE+NlTKKr
JgF8HJhJdYTaN86TUupdKuJV0XdbjRZUwz+s5f/V/SzvrGvHf75pY+7F8k7D7OeL
Cj3y8yxLkO0Ct/KfteBWB3x52l7YTefDPYfoVPwQ6wSidfZXoOGzedl8FQHl1HoS
V6M4CUq6tixbrkz+9kajSJk56nfzuWu8XlWNRJ411F1KIH2yXhb2E4r7BedUs35s
OEZU6aTqX9tqZ1s1LlIRMfi+cPdCiedGoxpaK7wvt0ZNT8W9mf0feUsOEE37pC9R
KKgTOZL1OR6YfyhvMlTQBspf/F7YH3kbE6v35mJ1OtdnxWFZ6V6Mav+b5DWh/v/R
azaH6GIQZHnlZTA/SFDVvTUhHS0Xi7+vTuYHCNwcn98lrMyXb6SJU+Ks/Ymk5NZT
feZF3UFcm0Jr7jVPQ4Vk4Ggzm+uUe+hxKDKJOkVxF+OzPlg2Xnp107fDnwHHjTHe
T7SxgyzGCN02ST4HbT8Pn8Hrn478xO6QBleZg5VC+RJAj+gZGdJZ8v1bAP0QWzVK
Oon8ZsH1Y5iSpxbnA6isFSbC5zNP1L/Z3O6b71nvOjbCXflndCbkXh3LPWg/K3KU
qy3TGhApOBuj9gMDI/yOqX7LtmGCd6JLdPFyE6Ev/qSvyaVH13v+QUfIsAv3V4yf
NIynuIrVB/aAvQ7NybQxUwqAQYtGkZrTz/nVyZDD9S5qfJ/wlfMuH8xKAJL+AX2b
R/3k3oTRgdznfiyKVLvpOSqg1G9SGMapWPhS6L/YU1n9wdbQfxLjUuBvriah+oMd
+G3WB2+BBVvjdQMLHWeXTmB1WADj0Chp3RxLCcT9MnaglIgHTHmpNk1CSRpv+rLJ
/E+rzy0U5DSaJ8F9ORla8qB4XcBzJkI7+wlAgz6Q/8XOF+6hzN07eENKM57vpAcc
gtod2UDzG5PgujzbwxbKyZsXgXpmmWSGr3IwIv6fyjyv8s4zan8Jia2GDPSS9rLn
nILlx+FthURaBjO8XI2hjypm7QuPv1TdCLOvZh1yqbYommHE3YXup7kmH766u2K+
XempbOVC0zBGgiO0x9t3kvSsKf5DBzkp617N+AjpKtA8IhaUjLLV2yPlogROVBZN
MBuSQdjWW/PhtdhN6F133emc0T1a6PpL5dAIw5RFflklFWV/IXKqGopv49gNPGGD
nkyMIjf3TUJ2wusLI8NIhFB3/4z9zi0qWdi3vNW3VjZbjEClOuK+dcw6bWUktlkw
XFDcEYd6JxXbAgOdOfWw4Ym6zuvrD8iCfuyVPwsXcOqUQi2Bb+mfPToQreW94YE/
AQDZ50Ef6urAoYl5j6Pr8hdTmiF7ge0X0ttP4GVQ+51BDnxXIrzw25+i9OudKAEG
OjIitfJenjs1HTP8gkNt5sxMk8y/KzQ2Kd7ODwu4BACXXNSVa8QeOYXQQ+ANo07y
nGPJi/QShlICIMxO0fJ3jdWvTtdk3zTldqgQ68Y2hVap3Q7mYFx/qCzcvmxwoirj
CujBDFimtWiZ141sjEG78/9hbI33PHKWg26pwvhN4HHINq3Nq2x95jRAM4RLXs/+
GdRa+8rrJpmNimIk2LXIB5czxuuu/FN4Jn7sKdXOw2VUAu+JEwTwKf+2tO4LKCJ1
5bi3ZGbKa4e5XyfGIZ0IesjR+169spcmkszxznmzGqh7RZDzDY/Be4Uz6/pRH2F3
iV70R4bH6+OjdfING3NuF3NHd5/eok9b6UsfZMxNFtAPB+6a5hqEIdN4X/+ZO6Ao
laxXzyPRS3UfOU0WOKka46X4rC6RLR6Q5lWmvl0KU1h44Q0XJ+dQ6yKSyirT+D2c
PDf9rhGPw8+l01IZpxm4GPbdh951D4NS1MdRuItzW2WS+RzwcE9IF9axO9pwAus8
QCkGHYjGNf4GREWkJg/9+L36SSHgVn+X63ZAGeM+e5Jjv59BKzlQprzIY4xg9IRf
1YCWbJfyHHcCxQ8J5E039KOcRrKB6+n1NgklKTOUoiTHfSmbCI05p4ZFRiEQe2TM
XVAkKD9enk9QTfi/HjeXU6q2SfYXs+VEgmIp8oJS53h4Xk53i0Y0VWjWqKIxAqaF
d74ZcqCjHetRVcXCPYCLV4BFjoUXe/ZA3s1yUuyZxdAJYIwjPEW0yob85sy+EjKU
YmJY9/WmRO4VPvq4GvJaej2abCCCCADGtVtFn2DCM98fktRTdIeLbvYdH3K34Id3
yPzEQ6ftzHNc60DxTzKA9ltVqBY1u6TE/kcEj2oszVLjTNFru9VGhmwcpox0rX+b
bJceIhubHPpdqdL/QAhb4MGF76KJQjL6cI/Q+iL7QjosCexJacEa4OHfSpHfwC/D
ZDPic6Z2uj2PK70EGaQkuQzBhB60kc2KsW+psJPrTvsyUDTnqkfxgBHWYKpsB0+0
Qp60Cye+MN04PhzO4QImnXE0Xwp4rerHhnSkkHsSsCTzi0evd47P+KFI9Wi772gO
7ohl+uqYUxzPfFvHjY5Qp/KgrPHTdn/yl4jNmJULpVZfx28gGn4tsWbX5V93gLBR
aY5zd5G02tOwx3wXZKfUwsGfjdwzSLy1bD/9U4mKrJRWLWvS3TGAMJu1Ys0hWz7i
4h3/b12m3RiJQ47IL6H3RfZm0A6afqJmA0tJ4FvcYQrN+dnheNtKdp0eBFg+jNL4
Ee7RhmC00+5yOzPpVCGsCH+XonjYK8YdXhj4nVIFk8wWylXtIpQqfdY9gQloYu7a
euDe86uV0u0d68pJ2UiE+axeOVcu/RHKHQQVgcH/xPvj8bmNVnAJYtv0pgT1818P
4cgGHwVkf+TexJW1VUVk+Zt5RDumbzIMa3HerrEFHAPauvidsdV4AuQrJXmLa1Zs
08aoecYJYToO00pNE43AYfoQzijfxW6P0pyq/AngxuaqKXZHXJuHo91ZUOwcGUjv
7Dl+g//RLtwPY8DG31cMycW8p2Bvjs7Z406zMgAdOpsGshqafJUCgE4gG1ew8ok/
ck2JTjNOwEJuJgZd9lylmOsCLrwMq9AwrXmNCiEsusTUMurtzcWG2lMFnMd3wiw3
z61aEWnmVLqOwgD0RcIoR/7FjS3xkKZpgyPNAOcEGZf+Zw3Lrm36+Y2CFAA4/f8f
pl6RwjWKpZe6sQ1sxBY3TqyhU3Fa3Doqz1oXxcik42gDalj542oGcTWwT6usDeGu
CalFCXLpmfr2EoaBL1SXSW5D/bDuDdcYn9HAmpnhHzQFeq2/5Mw2BZQU6iOu+BmP
VBrzKXt1/iMqMLrm5iWNy/ovaQhkEGYnr/0444tSzEIngNzvOucfG2QOZXwU44bL
xV78DPvJyMBoOoJng6aaNotY6EmhvVmtMqNa6Cb068mQv1CpNBTB6hKyTFRhIwFD
Ga/cod5cHtvRYDUC9LMcSgjaiLa4JzQf2YrghkbRSCZtdqsgJVyJp1xwWdkxcyg9
paoitYDWcDVR64tz1JmZjnoUEh/a9v7hR0WWiscZpFbYAaOmxvND+yVO+IWgChiZ
Bihvsfwyo+/B1oNF/7/bGJzDmIq4WlY4ubvKQOnwD1YECbfKRBwrF7iZt/5JFUV3
YXfH2uJrtkDj4TE4BZNtoaHLV/IlMlIlROPxRugrBKs9iAomBhpPs8/Pi5WjCg/T
mR8p6QGtzUIoWNyU/GJe5omO/BG2eIUWWWfigkoRX8rZUxGHIAEJ9JFOmMjJw/W+
oUsRHSphGDAf3rToTSXNjnE1p0gNArXlgofbmy7AKGsAxzzMo6BxIRByhBTZgJB9
b8IavHrIO3ar9OXb36zNYAkxw+hO5KAAa8VZKoitvnlM5Bxk1GH5wk+zhN5mexTS
uiS+XOoZPky+m1ZQ4sMTmwcGx74Y3dUcu84u4r3fTFLJmMJghAiej+6iuBAjc5Rn
b2JwE2ywi2cI1k5+arfD8aTs8fJopLUMzbZBp9gBi1GGNMscmKxUHDPf7jkTP/iJ
9WLs7zUvDWRnDsNCZSQMLQCbm6bMMTwhVAQlcHrxfsrZw3UHekyPUYkGlFU+UJzq
LN/U/SZmxMsdqs3hFctukqRWApjlo3w9VgoJnYL1N7OMwSQ1dvLQxq69lascrdsg
EYVUHxnwy1LmljHVJxehSUqwW5krGf3xSvqMsAZek1Ob7JjM7y0Iv/zaK7oCXY8k
jUiJUByPu0AHbzyvE4bzcZXE8svevhDLS9rihqGyYA+S2oxJpjPh7BbLiGGnGG9a
mPn626KBT1pFQjTc8VZgQcb+eYjaotf219kO5JIX0vVoRvouDoLfCPFRTpqKlg6P
oLpe7jM0P7rEX27sCGVXppnSALd6SGfp8qQTmsGZzpuY8CW3AEObOO3kB1QvI9ZQ
rGupki/1K/h1pEBBGj62RNlivoDKRwp/7lVOAc+rg6GMphe3/RV69yQw0wtU6AZ0
WE+DJ7sP/UJpsRE/js3G/nzpqT6ODHoAkIe8HX757V/5BRe8ubKukpk0ZSAqyuuT
FSEhs/KTVkoJ07+c78Foh34WSEeRMGGhXZ6g7gPJvTOLeei46zuWtx15BasugJV9
CQ0zILm0sW3fjR+hTZbzss4BuTikfvk89i8fZ0gKcprzGO9yLDl4SiHUKeoIlbXT
TXDpFGvXoIFNF+1XJjCWnQhvLHQuG407/ykCnG0JO31k21wB4qneHoq0DoEFlgfj
qTTl+ZbRolo2RUXPwoS9U49skxNoQ7BgL8Z20tKZGI/F5aIqOkz9S0aK0uF+lr73
NdvkagWqunsgbVV6YgXPfQaEaD23BqIn5CBWgK17SK3fv1bZqoZEm1WrsbZ21cH6
2rT+Mlqg8bKqvmyARN4SaigKKce0Dj0/TGMIYnV6OGK2PR0Mar90/+0AiaUwkFhd
G5zEUpoaxiqx0CPKO7iLlt7ZZObP8MMXGAKE7KREXb/KZm4OqTxxdh68L5FDZRR0
kHfp+NrE5BTWz3LPBFJTVFnWZpsWcxYKT+ZU5okHh7ymIf/owXshkozKEM7hdxyG
XvZxjnHzrtsd55VLreQJ1sixWK40ShI5TN1r4hdePZakKeERvXxAQOzEGox9s2yj
NsCLJxMGiOftW+UzvOefeI/P7xp95mgCmmXqxWAqaX0BFuouaCPOagO5hhDFDIeT
IjkAG2aBo52mTDjMOIA4FssUG6d7pugzTTs5WUEoHzM8PcLvevCKVHUJjjR2Kbj9
pwQsr+6NVHu4U+WTlOi2Zxa8ilXogGgR9Gx0+z7VyI8Fn7rAGoiisUNeB7jBDp2v
gxHMtbh1HVz/qUo31vRgTtwvXDkR9N5aN84HHxDMAffumRbbBitYnw823kXbJiUX
zkB9/vQa/xzkHARbbpMxb+Fi2KW/snIPHbz+ZthuYugYx5d/1UHBlvCNhAF65L2N
7ZKazqdxN7OBYZM6gFE9XLxYTGYTk0CQXP6YeCp4LnkJa1O/NyLm++CxbjT2BTx3
axDSfViFnpfZMSjW5o2Zu9vdvA5JGyV7aXV0jRahbwSOekdi/AmJ1GOUqtX049Tu
VeDAjIxyFMyiXbJqN+xEtoYK5hcVeRIjVZyVSUrFsXtxtwcU1N5J4hytIPO9yVwt
tk/pvvI6+Wmnl1jYRcYE9GaV+HNJO5IzPDtJobTmsJFXhwuQ/cj2hNMeTqwERbo1
CCGuRozRlt9RYJu61ExckhrPdMTKVYoa2l22Wn1sa/TquVv6vc9jIGt/d+KdLx7s
DBhEI628aFwDPPgitmHJMi8O9eefU/eG+uj5O5QnXkMyE4fJdXnghr/IgXAqMRJq
KqykCbW3E1VhA0zIhlUqurlSigRD2S3W+S6CAJex/DMj0ZQOnJejI/uqvlwrPZXl
fs0hNmMyr1qDILDjJ1C/+i8NxZjn7gkORzdZeOQ5v+d3CeuQuF73CDFuy15fm72V
U2OW3/GknNzMWfgDamhkeCKMpdBLdcsleXAj/uxvD91LFeg8OetjV/FR9/5lXE2A
W10xSH4fkNUfyk8GQWHpSsOSNZYqcwSNcPuo8iXgZQ87pLIDlLhRId1RWOIrf+z1
auoojc4eO87ueB4EZjdHmXrP+BGO6ru5Qy6hA7Z1zbSWa8/kaqkm01f2LEjZvQb2
yNy7O+465c8sFoyPvb6rgYjACb5+KHtzDYwjl6RQip3cXkx2zL1FnGCSxzNlnqOJ
LS+DuGuXw0Aoj4a/sBjNyWObHaIhMDZM4mfrAS7ThQmNFSaRySm/QIMKta0iZgge
0fB8MLBPNzc1b+T9t9x/jM3ATDcvY3ndK9DogFYze2GVZVfUG3qHnahf0JU53bhI
wQDMytjitTW/QlDrTgHKUtD0HbBl5I8zPdx6X+3UUko0RZ9jRV43Ry1SNdmAGck3
EI1FLOqDsYGmOk5kvmz0WwyNNv35pBEWurx49t99pEI0SfBB37JqqISEeri2JIpx
Klft01IZ+teUDvfQtI6j6buM5ZKlaYE6t3bc+0SfWQhlXTfEeRkgXcCwDkwtew/B
P5ukQqbycO3ah61WJeHmqEZCR39iys+Nl6PtdKAkzk3+WzrTDQluDBu1CUJo3m9s
6SNos9nHwbRS9kSLltQ8sjUKPFnVKKStN7MzQDOSSMitf/IdLACB3gESzEK5RAhl
HyT3WoPhKZrzZqiKDLR8hLNYcHjqyVu1/iVn2CkP9Grz7saHJFpWjn56W6RhugT2
aWIU+H08cB0A+Ifan2gUmFfX7PpjFunxaak6i40QuHah+puKbDoc/FQEqmoZEIAP
aAJfO3lJof/ty/KRJTI6+6gEY0wrbG3wwX0qfNq3yiyQ+/5PyXj3dSsIofACOkZT
h9oW0G8hJSlqAGCcL8Q9JyO0gByNqoNyGBfWXEloazigijUjjH040wRUyzLvue+d
GsBobmzdBdAn3hF+Fg3FXy2XfZ/j0eRxhhU7TwHLBF/UyPq36cYoNhu7wBQjYaE4
Tyifj+IF59hMQk45y1T6sout8TJGq1peZPY6pZRskPzgTJ+WbdRhWk/2nA3Tvnd0
xApK0JeAUAYBqTLwIpx1yd3MpPqu7obeB+BWVVTnKcMIFJ+EDJqeB5QzONEksnw6
hDUAQfkT4/vJZ/yho6/jPBbqL44vYWKu8KtZ3ENz6InEbzJexvRIw2xUoX6Zrjz1
lGnife7PuUoE/P6ZXe8/zE53saoxyyR47PhLY18aiXe7gY1C/A63zf5hanTbp18J
DvZVQknDcTBskNbqrHYbVfTzGIu8vllZUCIXMpWxNfA81j4X9k58T9umBXvcuEFL
S2ZD222N1/fWiiEd9UEvc/f6Q+JL/UcrWG8IZnxm1x/9/sSHIiI0pKePLcUbGCIj
kkyJbLW5US9iTDaE3KSpcMNhzwUDqmYy1yOKnEOq632/EOJewXh+Q6RLPC8GazLy
dWHCGBjeXTXrrjyW4yet6YOUc42AosX9pkfyBLac6d+h05uJDqldtHqRVuQVB+pa
rECBlWGGIsQ4kWpanMuzWgvIJX+X4Rl0cL9GNxVpcoO+wpD065VGZPu7pZFiETe2
bBXN5yunPltrJeYr3nD1Hu+EodjAakUJh7KWwWtq/S1A07O10bjlvgRu4U43JYBj
tqwoL0mEinGaf8JXWWOTO9KgE/rlJF6zcgFEBe4KztHqaCs90Z3WdaYmxkrW64OY
141CbW/VlQXxYSy8HrVDbah+x53rjNmd09Unf9+hYNmDFDxM46yZeRv+g2FnYWe4
WrKYDfiCKppopfuJCxeP594KBrx3ao/lPB5glWnozO/FmmoJuFUO8e0Hvh6vbZ5p
H0cZ4f7U87kzvOvxNxkvGCvxVU4SQS096gzRJRHrWaVr2Zl1bStNCxV0BnPy59Ug
eV3sCRNyHqN4qbGPKT9+YLBai+NJsEuPz3i7CVl01CZBpz4j21oLv35+pL0QBzGD
WbRWWOq6gcg/65Q91VVQPBoqhhy6bngawUgLxA/R2L3nQrsU8S1Qf0++PETmAQS+
KliS0+boeLlSRMxx/5B+FCPtUBZOeY8ZDdaFoTIfDt4dAl3NblnBQxNEhIAMc+TE
CRIj6Q1kgDp8m5RvQRjVMtz0oFPQ7VqAQ0rD9qhIHWi69klYqbB+h0DVNeEIgy8d
qHL5VLNWcKXwudu0YbhX7f8t+CnktIrpRt7E6j1bmUf82aMyQBEJ0YoiO1bc2BCz
ARvUBDmz/htByc36Ew/T6pqYj/dystr1fALfyI6Adc2w9/0utW4JfEBDvCBNIB45
Y8pq+10vdpJKR2QF4UXeHfcOpvceH86Rhi06OoUMQmWdQH221IfSTrAcvydm4zCb
uSNBOfTaColVCYltFghuF6bGccR+k1Yc92WRpgt9ugL/mtXPIjuksT6GDKqIzqDS
VIAwfYPdwUHtpbK9sM2PH0uC2oMT7xM52mXmxfPBmgyv2V/ZDCMDiBhfKpZiDAaq
0gMYpT7fkXGhIpSyrCt3kcq/7rT1Z3Rmv9ZL6ENbY9Z6gGJLAWpPea7JTLCB6AfP
+2qrrQqNCNmPvKYA9ONgifxFXYhRIiNUxOX96MDJ0u7SqB/DFGJEf/wSRyWbnoOa
M+M/O4zZm2GstNhV3+bEAyjHnAWVYXJsLot6yNglMSplDqpeAnNLekxhRl0ZHgk5
i4Z87nCdFvx2jwieYIO3m5Q0XNE8k/Fplhm9Vschx+zb/boeYw1WSklFtmRLcFbE
M2MaVYVM2LEWubLga8fL2atU6qQgrcEyRyUsvMgaNChCFa9k8B/Y7CM8MFDr2MuY
Kmzxay2chjCt5HVO1yCbNWTjeo5vEJzXArz8IBzVRJBF5T3a4zjfEUogXbvKEeAm
jkBj65zWKqBLUmF/aLq5PL0cOS2nADKGWFd2mhZ0Fef6Y8X3YhUXsv0Z/zBw8zBZ
h46y3nBdGIwy5R0l6HAlhHrEeT4zBkNH0jiUhwLv4g6vufaQ6JpSu7Hu1uRMtZnK
r35/eq6ccUHJEaUgkiN1VDgpPS9Wx+Awyjw+Vz/ZM+xNxJrzJbHah6KeADma+Oqo
JQlYemXa843HQrsUF+e+DfnhD1BtF/YmK1JlhWTZOlxFNoMTyijYhJWo3N5FLz68
X7zGXsysT15pG8OM6JAb0684Ydr5yckqTs7Di0mq5DZvmDS3zkbq0RdNbyedP4kj
rg60XAkrblAToq2T7vjCsx88O60dkop8jjt+oJCcyL1g3HKowUOgXUvayR2KF7do
dTKH3D35D7/w6YzXtrALCA4Yb0I1crvUvXSVtyNd+XXZj3JMd6ZwTs6+XlJn+Req
uFkjBalJ4VyhUYvS1Chla5OwqPE/gopW9eMpC6ZOjzK6qWjJIxxh/CQuyUIAMjRv
qQNlOIIXpoAzkr/rytEPoP1m3hkfe+3fG2lzOe8oak0g7dSp5K4Hys7/XQu5XnRD
/BxTnIrrcY1CjMnKsfu6w+p/ANDad+niTPMohzkfwq0/JFAhMd1K8u8iJleS7A/j
UP8RXKFAizZI+8WQpeE5i89DugVzkdYCRFQEonQxDr3SIdWpYdyLx8QMp7+AOVxz
jj/FX/fuZq+oDmbWrOYir6deArXhpRVzJYq2HSQ9vkkjDdI+ftHjT578A+0+ln3O
b8lGdkHHa+v/faWvEXKaniRMoIeeThyONV6/ISANdNextENNHaK1CiNxiWgD3BqF
uo5dIgEHIrW15Vsvk5fpFPt59Y6KxCR9QuhrT57ybOr4eHfHIIC//ZBwq2quMKLB
+OLZVPX2yoorKNMGsgS4UEMlgrrPpcrT2G1xjLzlSl/8Dn6LbE7Orb1/cOm7l4Cz
1Dy0FlimSqp6zNX/D18Voql7PTdsgUMqB17LNNq5i7dwc+6W6vDJ4RNvLhZ9WA9C
Aa7+LXzm8Zp5/IFj+my1nJAu2RAwPzmWPlSZRSTyi+3yJ6E6ribBAyVrsb3M7goa
3wieYTnNmIpdTHtm6vebZUuK1+0Q3DIFEyVp9EJfJNuqH/mmj2r4cIqCiFdZqt49
+CeXv/VNgfhKBHGPTFNrvcacW0zLweT/o2/Hqz0jF89st4M5Ko9f+7qYXMlUoRtP
gdp4pA+YAHWRhl1WTlvNcjVUeCrI0Q4X6vWv2diV1S3Oqr4SuAk8uFe9Vn15RbyT
6QcxuhlBu+FJG5Xgbx9CusZFSxYLrzTE00K6BKWIz33waJpCAXRKUOMZX/foa+vf
tNVBiVFxdyRXBAV1TZy84aCJamrrNZkZbw9hzMtrr8Po0UydPvADtVyiQn5W1pz8
A7sIq9CtiPOwzNMoDu5HPuFeXX+pQBtfDzpjIjfWEL6MDJiubLHAIv5xo0E90IIz
9kixdWepbooaCS8FK7LeCloaev4I5Po4Y/NiLQY4lBwmChnjKYI77oZZfTRc4Et1
zVp5Xd1ZnD95Np4f8jAKCNhcLbgcXURk0LAohvtlKhLBJWaXHzKMiYvJIDSeau/B
1GrpHULLsC7PBo8mv7xuLyvpnn43OL0kDHX1SBIPmUVDPc2ykU5yJZMVgbBwosBD
odGHjxiSsKqfsvLBF6Udz+mQHtQf/KoGlGUvyrQ/BtqVFGCgFHGlHJS5NDzc/qgs
IkY9WmOZ7Z4m1fJoAjLLmAGYoA2C3iLFfLjOVAepooKS/DagzJ0tZvXaoMLTveYB
EF6dsRKZtAxiKRys7yKKic2znEy+Rgg9ykTSM8M2DplVkOIJ/b7jIITpcvDWpKFV
PsX8eC2kZOKsooDdUEiEErgkydTqu7Z+6fYkKny2Eo3/r+RChpzWkz5sEWCEUG/i
60ygzLJx9T1l9ow5vb6HK58bhhuSpGXnWZW5MJcnsiiwaIchWBng6vWLIHBpSSRH
vwXkZ3we22fGvJH4kxk0OVPXIjRQcgYlU/cM2yhQpmB1TZ/W5Xlyr0Yl+wwxIS8E
5xKC/T0pCKEtVEAVdMAZSHN1awN67AKcWbXWhVKP1AoQpPa6YJpqCkwe4tPLBeR6
w6lP9KeozbgtRBHterKeyVJKyhaNNDnlm9ISyBnutK3huWFStUEJORHhw5gVUQue
L3hpaUlSUT0uMEpZacKsTVxJicAtfaKJ/CPeYJZ7f7zEs1+RMpIZR5m1LBF9ZUPD
RhoxrZ6dN2SZJ49cFtg6au5RO0PbYXHtAYsrBQb1paosY+p3O0hNbZFsgB3DXKaU
wB+D5GHIqFgn0lx1kCIBk81s8aS/j63p/K6aiE9W2bO4MYu52IbxuxQ27MGmd4GQ
cTMKZLz5yiFHr2toA5rSLEWYuXjR47gMW+7nSkoLRMdIPOwd5aIs2dTOrA+NbQ+V
Pjphwz3AQkCeD9ic9KCZa35ry6S0sJ1lgKLMH7y5p0YXAvPEhzizXRwMrn//cAvK
67ChZfIHCfWQ7iCu2dT9OG2MzVXR60hoom5Y8fE34go6quxwcRmQbuDXzPkUJPXn
ynykNx3r/XlqsrjVpGco6nDodOqvFibB1UwVOwGi9aaPqCT3UGQDjP/fnuHPgf9k
QpkFi572fVQqztwYzdlBTHt44vZmeN1JE1OhDhAgRFx19qQIfCuIrV3wd61hLA9w
N3vZvCTWwGERE8ulukSrQSoUVY82DQmY8Xj7XVa/y0e1BtC6/+BEBtqxeL+qM5Mf
OSJmTREGTTBGg6OARmQkLcasoGlymgjHEXoI85BLr+dT0sBJ6uaz2XrXNLX3/OD4
gXSdam4fwlR8a5O64ncZola8rgAw8CkPare74wVTSVz6DiqtORr5xGh/2YmWxmKs
fOVrZUES07g0KzH6HLCIFMAO9/npEZJ4aBNmsHDfRYP7BLoibWGLioCIV2vCkw6h
fXzSJkiDNNnVp/Nu7JxyL4LwqSamIwspcJ/FvLZu9+l3ev5H7M7PPJcP8M1uAybj
RLXSeHCTJVgteOAxjxVimV6QLWljt0UcJosxTiGuOsTsScIRIzw+wWQHrQML/laM
4zrCqduX9C37yT8S5RbahHGvr5ccw+nuDTwZzMKQ9VF7pxIgYgmbPedzxkOKFEn8
+894AunPJeVAjPSmlxHdbO+QvXUYGvx26wqlIm5QkRzYjDc484EuAcjnQS2YcIMn
cVIZmYldIakLb2h+F+LRwfJ9VoST4cQb8WhgpBPZFL7CgR5FwtDOXNn8gp0cQF05
gr/gPH5d832OV/3A8NXosofZTMUNHR0nRBkbc46qKjEzLu7zV8eh+uuxZNwpGHCs
pzlPNH7gV3zQxAO7p1/c0s7qogzEwzXT7xFsS4ZxgLSrX7JajYz/npMf8WcN4yXU
gYjRclbXw1rTuryfcE8T2bsGx/BTRsGtKKW3NzeuHyn/WEiRf1f98CD9TTZV7J5U
RthAaWbn7i2S6sWR4/OhJdAbGG8g7eqH18y7TmgbfA/130eQ8Z6v8gxNjIxf7HZj
ffJ9U8MX4co9Keq8BkwtJ1xDP/FYo2R58PL97bRCVtbs9ehvimG+uV2RrB1DVCuy
sf0/SdajxREKH7pw9/pKyj894dmzrUK3KrVypKlW/+M2XsRqsydxTCHOI8jiifhM
ewh+saQNgpOoYIzVRAsrcMWiqAqh+dCvNFYKwaN4YxynTGaOr9UfxKncCzbykrB+
34+VUOFjuS8Q3h9o/2Yr7lShXZD4Z2IqbGRUDqUXQOkwHW3afPJFxdHhL/ClHuD8
x/tQfkRUJuE9WHWh8Ht2/Bc70l5ohjpzXYyyB4BERoJ8DnflzLLdwHMEigjnpcOm
HnKYhFnOB2WHUBJrw/hONbhUVU8/Vm0QDdrKg3RvtNtzkUA96mz6t3Jrt62v2Ugm
qLMvY+QQhU83uE5uIFae+INJWi35tYtYacnLd81AN2EbIj85ZZpw/Vs4ZabbCdxK
yd5TuztpWxYXORywfPk11DcOa3PTpm4uNPsq1KQtXFvEyBVsuexNoekPd+IRt0+7
/NZaGm5u4Fc+azip5EDNhohXEpqFkSduVbeuLneSPOOtKi0zDMRyQyQodpYtgx2d
y1IhH7G6n+jkyXqMpg6zotPN3XwdQNQC2UendzqZZ6iuV6twCcckfB3DIfiA2/Mf
XPhSewIod2Zj1CBKahoyrK7cG7YLJ0bfQ81yuJxlMKutOx1Uq3LH1ovY1lGGsb6R
3QkQxZtR1IJm88d2f4YoWzofh2zT1IfYgo8Djx/WWYvINw+ogZ2AJchSxync0Hp/
a38eY2KiAqmLAygvFC/LFw/tfIet+jWeWLeOVEG96ufD5vfypo/rwuraTTOtpTeT
gs2XhuUW2NUBN0M3GSf5fBSEXdsCR1AYB57+b/z26qkjXwBAv71Vp3FiClRSYwQ+
JZ+oyyQWsqgX9j56q+y/4GjmuR8nAzOLkazrgvSqtxkge90S2aB+hyjeUNQxTQ2q
oXnX175eDGtd3zvQQYBzy/AUzNue9izx6aWSsWZECm17stATBhjSkPJJPlGhDUsc
cfeGWbG1IqVzlObECYM7SxJ7+T9TmckY6j9xr8BOcLQEWelfXNOaQnsTjUYeiJgK
F517KRFI6sdzwLfoY3XmimTHn5wGAsWMbpsHyhMfz1mRDrVIo6Wf+136HJ2T9F4V
KQ95ocu6EaxMlG0cdcR3Xcq84J2bW/vv10xATH40JVsKFPi2AvQb9zmVeK3HOL33
v7RXH7UND3NowJRpJoGBqecW7mCtfAg8lFK5ReXZl+g+40AVp18IJZnz+ECJ5+Ts
ZWw4Uk7y7hMnUv5I3Qhc1VW3FFUbVLxkOubt4Fj2XaGm9EnXmvEp/srRLOMAOnq/
HazkeacGHqg+2LHvoYuQJQASwBbvQ7v+Q5QSU0WZfOvstgKgxsGEIQTMCIRTbRyw
mm+grYuIu8/Ozf4Ji4wjVl9iOFPrexp489bQHJ//TIL6xj3Z2NeXcrJaFtVLNJUK
Ss4qlw4XfcHCowFsVf+QX699i6qOF8YQs69iH++hyaKqITQypEZVE0a6sZdfh8S7
1tqrSteX9HtOP0PQYINnUdOHsc3FBr4z2NdseJIJbK9lLLv5RwKBuFXTaSQM43mc
bFQmhEi7KzPpZUU6oH/+EqXMnhprfJBiQYIwN1098Y/UQ/DSv3hJJ2RwzcKlW7FH
G3PMoFXSF3uMDjArtfbQ6cLbIagnTf+qj7VPW5K/3nej8KQ6h51rbgIascFLrboa
QOuuzmWdFUAA4QLWwQsfevpfFatMPP1TMjl+CogQo9T09xGFWG56F/GqKI+vLTx/
iezu107/+97GNZhQL19g5/mVX+md9TPsMrZ2z1AjknkAC7DsTXEXVOWnWa8km6ie
vq0VDbQFxkg5kah5qxJmvpocAtj/PCdY59uxUP9PdAntCGZxQmfbMe+6dfmZQ6gb
yyflmg/48aRYJitW8rzJmI9LcwA6lHArpVusgtzrMXzF8TB36SPmWJXftc7S9z3M
xmfJ+7QjGEZCWRn6tNvL97iWb0ejnZMqolH8Zt9YUqTC23Zl7eyavCAOwSLBRIxg
H4uXFRHRI8T+xRAOQJxH1OzIVKyOfWpSSq4Xn5I2KwPCfZfhp2DefRpKGeSXYFnn
CjzhCDTUIazAUoOMLBmESEJjToR1/dqDuc7Eo6bC6F972Vp1iwBjOd7atxYLDV0q
QJfSbjy87wHsahXmwlhSqt8Q/wiuqH4UBHPDqL5W00d5YS7FgG7FSExs47pP5tNt
B0EdZakg/21N1DLmhvyd3jxrBL3rActbyQ7Jz56npY5zIUhvQyzpS6EY6mAOC7pu
JlrqSoiY0SHA5YYquDe1xoHQNlK5caEbGGQ9yeom4C3nQNfjWHr9WO0zh+PZfhxY
E8vZA6Nypmy3RrEFBztsmIuuQZ8kaM7PAytBLXB9MxLtUDD4VdGtPU+cL59Jqk1d
E5RkKLuCtcjDDYyeKuBgaY0pNsWaq2TJn2yP3qI9E0MmwMD8doHoSJ7ZIMV7xUkx
aPOr9II9mlvY9XtOUafjkj7uuEvnt3qA+G2vePM7u346wCd39eMKX92MQ998/ENQ
19/uZStk89FDJy+i9C5QX3ifLi13FJydJiyd1W2/HQjEOrXST5wPAJPDRDFVgSOX
YNUPc9s1oBq54jHhRePYM6KENZP+InFFr4VQFoWIR/rD4mlr4CMb2rrGHqtENQOL
Wlti35vNfFhpfLABRMh7exKOHJdokC8CzIFuoRnoD75XI4vvBxg+Uae9n4Hi0tlr
bZjFmKQvNpbtlaXTb8jLsXeBQRlTmiF4UsO+Y/LmBHfufDDcLOwbEScMWw4ONK2S
N2c7XBHMo5TmssdmxIFAClOCTuV3XYeAW6m9cZs65nwHa27wLP+XXtLQ8CvPlXLQ
oKZP8JDQUkZvv/XGR/yBqI3PwKH0ggGdVSNJDx4f06OCGrtIX3vInPUOQxLGhema
7TRrFXaeo7N3BVUzZMjAmQQqMzP1ONO8nhSvFgtV83Rknw+jRc449978E1C01Yh5
xkZK3b4jcrXjulNoYs1O7tcJ887k8r2FsSiYcBsuAeFGCfs7DMDZ4wSu8LTXbfna
JyMFNrLP39MK7D8rt7+Upn1g4Y4D59EblhWV3QorILhOqhW5vxNqlah5hDHRkj+W
ecR5RXhJn+uxu+2i2/Yo3c/vDQ/huEx6Bc70kry1rYR+Zyc6Jjj039QZtgRoxQh9
ZyltkGQguC1LPJYwHki2NUrVUwaG087OOYbGR2W8ILbmHqrB0Zs2JjMYWkc0lpvu
J5UpMsSIx5YhpUwYTH4JiYU0F42AcjZ4Kg4Pm+7aS/d59Qn96XBLMHwUgwvQV+wL
wubKiuqdwFSqbRuG1qYc2GgQ5HgFvB5oWo4vBn2BMV6yQuclPMG02FTH/vS8RANs
XDqqZrvzzFsJ3MPbOszUwJVNVBVMpzu+kdQB8v3fBCj74VRzBl91ATSli+Z6tTC/
pR/rK0Pf44w37+dJoSNAVMSaeM/C13zs5YPMLhxN4HtqzazhQaprdl8hQvv3W8hT
rReVNTddmnmWBlwrpKGNXHfDNUJqysyaD1/JQQPkJrUFdEy5BT+L7Ve2TrcRCyOv
fhB9X2AcVsL63pQTlnuIrVAjg8oUqIrNjVdkEzilDrVWn4fprVa4bfuUgycprpYi
BPgt6XpuKp6qV65iJJKQZQbkmSSWk7LfK6D4SFp5Xvs0KZc9ZsVpUVqcnkwNnk8x
QtpmQUL8ELyYZvghyfnI+1KsxC4cC+YWYUVqtJA7oZJYV6UM1tPXD5rZdgcxbIRA
bovsQmdzJ1mOUACyVlI+JeLTfXpw4rb3lQ9NyCelbaA8HhK6OQnLImz+GTy7Y6SZ
J/lfBySi/w7psnUZEzKGmPoRUISRh7VCTKNBN0D3S5Wd8HWTaibUYbuZHBcTTMwW
9N0iLysFfzFHcoIJlNQtPVCFjAxhUPZugr5Lfrp09JDzfN3O1Hq5wnMrjZOT39N0
ZWrvpUciV7Z+vnvmRLsXnnArGIZHi4AXL8L1bInmvRx6XYKq8x64Q0g6+817N5ty
y3vsoA1xmKm+zySZzEEKjFG2HHlGTrtgGC13iPpZWyrL1PzEGIxwBuReULUFf9Z2
1wAxNtvL1jXytwN1fDi1A7slcEr73FQCzmlAx4nazVZkCHrqiOG7U8MH+IDzGm2y
o3GaLBZxvRwZhbXdAYSGMBhY3iQUN+D/thraeha89siZMpNAWIvqc+/ZJduNz3uu
w2GlMZbL6RqOZNUqNMcpzHgX4CkNs6SVPG+gXw2/dv8U66A11FU1aZudVF9azcoT
rRI6QvH7XgIqNYlQON1nO//Bx5f5hVjPkIgE1m5KRb2EMQ08KGmd2u2SUPYXXkGR
7CD6M6y8pOflpxDc4+kEduUxxa0Fok/acRSl4BEZV8s0OXXiFnDtTou0OmGv/fkg
MtyjFyI9T80QJmS0IK70BlLmOR+46kmDuAgLJWCsJw3pMR+YREJcGtQ5Yeh/Sh8F
ZpNSTro8Bzxw19UiO6G6ApSm1HnyiW8B63UWgcWPPIv0LiE7z10mvSYNvKG9Lpac
GfkGczRLPPnkW5bxRB3awuDZmOoBbLhoS0qnbhUJ5zZugqeEypF+INOUh7qORyuR
39O5YiDxVkDVJYa239fimYqcMQjVGQvBNHa504p6BjnZ+au9EEdSgKpKRMw+zlno
im2As7SrzBElFGGpc9aFY4EPpxgjuaRViRLXDIFAwtGsMgKdPEQhJofPhEnn2iZV
0HAIlkDFvOA3I+4qdbVQtMMj4gAB3GrStbC9OOKDetsX1In/y9lYV6Mgi2gqGVKe
YsOiv49T4ySwOmPkeGGaQfeuptBHOGJJYScyYaF5F3XamSAUQm+D5FA47qY7ux/t
05OHEuaYbP0Jq0/kdxHeNX5zMKzJCArf9AjKrMnVXaIKSJt0nN5PnEA51N2pTeKP
YVieEulv9fJGXhZsTPdb3GpVZVAD9gSJQwcf0tvULRBmkGKWxjECddw49Wu2mEzi
UZnESZFROURWggfEpWbCJUcFKDsfmiJERcrlPYN1EhJsSwsFH3VBfIKYHGpZ0uJI
HpKTCxyZLEvNLv5neV/DEmcF5dLTvzMDbcgPkg8W0UjnLuTTHIdyPPxFr1yN0yzc
00ryHGLN/FvXKkD5Of4Vsjx/gEBjueCJegb7ZQSFrnRlmnHPXmhcwgmQ83fHgFPS
nDaBqGTn98H0F1Raz0JXJtYm4+u+9KEwEjeIhr1x3MmeknUD283CjqgJ5ku+G3jh
2FgyDCYPAku1ereB1zKrhtzrsxotK/VuIj6k94K8mDJVcwO2TOAcjwJ/MeDMvcT7
+oXd0ZBqTjrTkr7CPWzUP/HYfhJxmjy66CXJ5xR53QtmKClX+FZSRXXBQniiq+pO
3nfmtwYKZWvovSUmbW+zNyqMlUFA4kmXhPqVvMcJzAzyINMCszBRII/ESEhBk+mc
sejNPYsbzp3iV6eH/KOJy2hKNTQeiLhHnftu6xWQLmQwRGQXtep89Neeisp8buSS
5Bua/5v+QD1QHWDILOCrSPpiM+/9W1lKs6T30bfk+Xqp5AYSIsoidbU6mQMuFW1C
OQySXc4Vps6avNSnJedX8mBcdHUwEvu2DU4StUPsW6HHPsoc7wVzX6TygCNZHgxO
ycLvs4vLuhJ6/TwgTtkfj4J/ewNMpm+xxKhvZe1z4UGRV4Ldzeo+Ae6jQb8MUJAL
mYy4ThJE05Gfoak2fAsWko8QGtRg+kqeFT8t8OFC61YP31XZVeq3B4VZheBoFO+9
agDsnq2YdBnqbiDZaFdYOdb467j2EjcTt0bVpJPPWuZGo/oPvBbhzHjzKQ7pDGV1
K8DelOE/aZns7nKUoN3gqxOQ+lXWeNNs1BhOij1b9p7DoS16e72MAcYRt+YTJYiQ
Msr/esJ+RTwCzDjAUpVhxMiQGNAqT3Xr4YT75UlMQAEwSa52v5gIi00e5xnOiij9
QMJLbvezxvMHbnynU3QcXuFzjECr0wM4ghOlG2lpm4HVQXRx+j/1AJUPZ0wqliuy
OCZgEm8ovyBkBZ+Jsc/YpbSE5PTXHjapJ/0yj3G2RKri9IaK566U5Jtr51OcCAcp
1L+us+AhHVVG45dfFHVIJL/mNebXdP9ti+lFDwzgJIXjOJY1qhgAT8vPv/NSiz15
VuuwOaciEKjdu7beBC5dzkabAeHJAe3cpQMqeFzi5znKBRgxA8Uzkq6QYiNEHT9V
U2eHvoxu2jmzuGy1b+lfB+EjIN56bVLRetJqjs2zIfuogRtPsASaFqJ2vOSQWrvD
QpgWOCc4B/9smCoVIuXOY+2FkJgdPHCbJgqUKThau9riuOpnllY4FEGHv0eeikDl
vZ0umVLECqHI5o6k1Tj9VwZ3Aw/B8/POOqFWKCqmG5UBnj6JImguEvcjLP3kSxyv
tb8yibq8lUjgrlqZnTbRU6jg+i7nmNX03TwHEnnsSujFJLrGLMRptJhOtwLJhuCT
/MjjFwWhLSzrtJca4NIlc+ZStgH7XvVOO4lCJk3FYhZfuq+F3j4ZhHZrVwV22LJ7
LWALrWBDxJXNSfL+p1Qh7KewF9V9XjK6nocsEyePh7FwxJllTXI+NDpqQz7VBhJh
s9I1hz8D33QdsNEYLonVkwXpqbz/7oVrMd0QBG74xuK7pwGwVOJiGLGc6/E/sAQ2
vOvuSs+TwWHwNaaaSj4MnLfT+v7/BPGJMGvxcnrgIxOjzMWV3zeWBfXZlHowBP8W
YJUpcRvlfBp0HEdIPuVP2Q+4YuLnWVaUTpApB4HZxA+Jk5RoHmf06poSHe0dYn2B
8pOhDcTRdv5+KklTBMOYScwIWL22NbeR8VT7P7jHSjjSAZ0yEOYXae0RFgDbzPo6
GPMihwI3OYB83WVYDK4OFr9Cv+DBYh8yrlswtXCFlG0u0lVmEt8wNOUWha8B/skH
3W7806d1Gr/6zOces8d6YY/3jdcjiDZ4T7qdYyCxhEHZH/tzlpoFokyOTVLOrqGw
Fe9fnBXb048SZnlclMHNDcgyn3xSkiVq2heYLcRsib8aUOGJahBxW97la3ZFO8za
Xc/NZWWwpFT66J8OrfIeduJFPvjSI5/Cwy/QV/twhJXPiUTxW6QXvkLYf3rF6sZM
X7fETi9qEAT6WxmXMFPz2Sy7i7FdnlfgZgJkuGNH4MBczKP0jwLycI/ASv0DDnmw
aOowGRjDd4QUgs1A0flXDuroWmOYttpwgZaJ8AlCjmD7W4mHFN45zaXiy0alF8cH
9O2pN9VUbJhRJ//0c9m9WcB4WerAeZGojgCN6qCv/vy92k3sxWjBfna3Eg6rIEMd
soZzku2g2UsLaNH39lNbUm4MW6r1GE4uLwg+unWOpGuEOMIbnSYlYE0UX/EkXPPd
i8esQerfoc7c/fmrNZ9zaR8BnDNWiyvRBOqURA3vrc8KvVNcJhy8R+bPqPt2HoHv
AttCtRXLYZaif31amSH9I2OgteMyRmkcW+algosfcbM42GPWX8+dn5ZZxdct4Q+d
uNhdZumxEpKPH24dbD6dRUPVtvy9ujVgT2rh8Q+maIE2VYBSJ9yCB3nYSWyb8GOH
gy5nQnfiS65P0a4BX/HxAXcF7GvXtGAuFR0li8GQleb3V1DB54wiMIAqpfNZGWeJ
OiirAE7fL8hnN+hB+kRy+BcGRSboQy6ln2JnlbZLltOljRIfQNPPoxCtS1PoHkE0
05RJum1fkYzN/HHfV+skQmlar9CevgOlpgOdjiFObMyTSpOeSnYsmDFpAddMy4uO
9/B2BZjXifQAkdcPjI1WPduQ3aAkGk4L0uVGk8dZGW0+cmYGQfOzp61Z2+W36SIa
kCtzPjLTRBYlr4GY3IvpoTsQDMjxkoNHl30PFILEv1acZLl6vVDi7iKHRU2EYaKH
AuY1nNnO/t74KlTZLCD18LdXy6qcRdgJlT2sZ4/fchUDquSaRzGcBF332EhC6ylY
/Eazzdmc4BV+l6FSiVQazdyU4OqkKG1HYt3feQu30XOxNqhkj63VlF8W4/qTxlQk
SszxI947XOfVQ9hQxcMRinBSYYGAeF4Q5UO/QbBYr9m2TwTWj6hleI9cFJuZ8ZIO
X3nlEEveGts1OInmIpV7kU2W+3GgZVkj3khffWoAiBom0DNLNvn+41RoLcIVLbET
qUkUnYsckNRMnh+CYOpVyInFPaIEPNWJUuruk7WaM13Zn0dIqT5t/hXSjN1apy2H
ADZN3hk0gHq9nxhZJz5aT7Hy4Mk1D8PvDRHIZzrvVl8p1hbJo7mrgx18kmD1vFGk
ypDda82qVs3VGRI1/Z38ZqVnI1hxcawX838rdDxOkw/BI2/IAcIW7Ria4szGrSuV
fbGrDdO9n1rGaZeoaw2yAiafkd16cbPFaqNXAUO2R78VHr+kF00Q8Nnwu4/IEtoz
qmQFiugVvX9vOpVUWe7CWpddw85y45R79uL7ThEAQozk7aD+78fhXg8sS15svnqm
YyNlExh6L9Q9+IQtbK0mhR1I3y2UnOz32uxGl1FMr3YMjyVSexzxUbFZ6qj3Estn
tRnIUqT7Gtj6nMYa1206ihQJH6+PJUmdZSZAJ5PLf4YSeliqJGB08l10xT57hO9a
+APGxCd1cyXoZyF7MwUwHV1VLS8l1GT12jeyeUEpMjG5941v4gX3P+dgDKdDKMDs
3lcHBUIkJspTJFzUIOH/nXibAoDKa0+x8bE2Tq4W8uo3b6aEha580ChsFJY4TKlF
vbzr4Pi3nKnnNCXJZJ00QrguRlFWdniBmto691dNnXsG2cMaTOIXdiA6xslOgL/i
76Mi2o0k0yMGygpc/zrF3CksNpBsN6eBqyoZ+ZJYowwaH0iKlJlbLhh6kBfhuwDi
XBiGQCOoGZmocbpVQfiYW8ujgpPmQEzsyAXyKlLSztjd71Enz21NrsgMUSC2R+n+
J0Nl9lfAc6bEbY2RNJmy/w==
`pragma protect end_protected

// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.1
// ALTERA_TIMESTAMP:Thu Aug 14 16:11:30 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gdy7sAtJbVO6nni5jVkB5fJcmKjTi/FNQpbxnoWnP1gwI07PpcZ1FraX/FB/YMoh
w/3/bm86W7dKq8RN+xAH0I0qK9wfO6JVR3w6d1XeEAZjXpfMzTm8e9wkrYuSegWV
s9qFr8G7HQzGgQkuTqyN4HjaaFx+dKzNLkM0A3/iYAM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9280)
GxPxZbbLm64vAW2eRsOwOUd7VkwnkGfVObOwCOaJeEDOtUPiiSWYNL1E976FCLXH
5qndm1DepQwyWxyNOI6MDtmwBvJAZ3x4x9ZS6f7blFNoi8GY0I2WQ0K/lA8kd25U
3rpHQTd87HturI1iAkayNjvzQSmVygJ4LoeS1gQcUz5zT9r1b6vMFDO8bQj0crO8
sni8gJU/ZYt0bQCR5jTD3+TGdvpeTyCoHlmBt1HtbB+rSkqokiNI0e1q+EU9TwUU
T2QUFRUyEFcHXZGGKkBc/bX5DCamkOod7oaXT86bVHmyFJTgJMHwCf6qOWEU/duX
d19JlZ9KobNFMf+r9Bz6HiWf8+0dN3TOH4ioXYBsh4aDgbfJ8FsfO+h0CgvLQvGI
zaTVP1SKbxfum3gEg3KDOQX0aEPzp0gA1LtKVuFicvnW28F/8Hvhe0PVILOYAoej
Fw1ZYTfZtTGA/jqtpF3X6jTvyj/Dw61xqUAbem16HcrNDWVHgLQWZdQM9MyMqgJX
Dg7iGzQDpKc0fbAg//ulsNmDX2xG9jEt4fiWYlPjItAwmKdgVsHnDPynLQiLGI+v
WPox2VVVFS+B+LZPtUarI8sTfNFWTrZfw8lN+fsK2njl2I18cZVpynsOiphNrlzB
Kj01VhqTZ7ZEOAC7Y7bnmwNc6NGu5di/TBRY6RC2lUhDJ9Q0f1OWJMxT21/vKnMg
JPDTO6fI1KluyutCJvIgI3w7tTp3MeUyOSwSk0s/7GJdTEYupdCC5uLpQiqF6oTo
pg/eilhnbms5rOnhTc5ELUY6+R7DvMjw6xMGQWeCPyjXayQIMkfoTuT62AoPxoZE
8dSB84bgFqBARTytsjirUvZoD17lu75S5muEFEmrDESYX65Fw6+pRDp6G6jGPcvu
j8iLv2B20abVzc0hlW8P+S1uAAW6MhozCbJwbUDYffC4sxpB5G2LSUw2A0AEN5mQ
+fFR/Fe7uzkCgjF7w46kyKp3zD2IrLsJFlfpPtgM17QbYhqYS8QISJCjZ+XX40yt
3OGDwUFZboQlDJt/uGGs4h0fYwQfSq4C7ds2N1tO+EqZ3z0e9gp4zGOJYsVpzhEj
eNy8cgb0oa+YF9MlV0ZEpycNkWkWiFscZGxUTQBLCYeMLzdUitHsT8ci4sHQnCUd
p0rfraNIHgp9tkbWKDVSBv5lZXPBSltQhYBOg3oAl0kOjMn5tD/6/D9urknDNzLI
kW9TtKCpgoH0tSJqpGEj33whi5Ty24vdKl/zGKv6fFtkiS4R1nI2YuJKlAzbPCd6
fly9cUp0Ea2ZvYsOpjqdDi6+EH7Ml4c0aomqv/dW8yK05PQGV6CHmGtfKuSTCf9L
XMTtFWJGtl2xMzVzW3S/VCJYvILqRIN+bsfJunu5K11KPPNiPcVBaUBzZlphxvp8
P0isEbnJc2S0UGbTeGua95/mCJvj5qIe+dAZvV8OJCT8JZimIATTNAihp+6+Gudb
cyPWclF3GlZUPCfrJ/toEt0/Mw3AlBoi1WZrozBSwzUBtDnqdd1/wRYmrZFk5mQb
DaPNRX4wqEBgAv2uIY2aYBSlKx8SqvcxjpbLfpH92eq3fQC/h9AgkfM1rYlmupyM
iRjy4JE82LyPOWt398foyICw9hKQbUOYkPwdfIwcdDv1odyEUZBi9DKFoHcBM5UO
RxQtsUJxycIdOiKqqAxIJD+YxwOMLly797nxcsoe0l1jJbJD+4vlDoETMBpLP3m+
VcDgluUTnpU6IqKiS252aIyFGqNAsqIOVj91pFaJ7qpmP7qxJt8qYlgpymJj1GnM
aowSm+J3lko+1k96ZOG5UrMf8VckDnRwQgNb5jir1VmEqaa6KPXZMIxX59UB5Xai
6aaS3+8Od6ttqLd21Bm0giaE86A364aZLT6+eLUO5nXjirnxGqKAbuEPQV6cjP3p
D6zM71bl9q1RMFGTUTAb9iq/V4XZw9KsQFJe+IwFBVMSJrqj0ZMJCtNlEvsB9zll
osWAmhYgjFBngUpZwv/Vn82S+4SUWeMqtxEcHdgw7Ml2aBIuhZkvdVKKmLbfwS1f
CKy15GDVKVe4qKPGNhEEAeT8R7vdYSAbplHOypCIj/XSu7U7wtHRiDuujZKiSsNq
3EFTyzH4v+6Hv19zhIe6QWW9ZSGTpdqTZv4SqXlrklmmVwI1+Wi32yQ9ywgefXSw
65KVeXelhxlJIsQIko4IWnBkCpk3nWyUWDTAoxlSR6cQZb/Sk/qxr8vLpisFmuT9
n449eq87A1orYBnguBxBQ9jSU7EXwGyU5GyeMXcAB5b1GCx8BKlhPd0fA4MCgnPW
FKqHPd74CTtkTsTQ7ryZBC1PYcKBqNlk0YQauH+THosKrDvCLwGCtYNW4o0vfLuW
D4FGizOC+LX1ewIGmNwuFWxqP/G8sNlG4zaOt7AHOUOiPSAC8H3EDqExdvU+gUN7
hNqG4zNUDwz3xqVJHFvkymwmmq9+MsX/EoXWg/waERMHzbkpL5X6wB6he4nhaFlO
zJCZvrKaVNKNV/m2hKJlCuIf5EPRzMnib9p1B6fpxVO9A8+4hIBr8SiUjPnFKvHH
mG8HR7h1ZwMDqohT7ZXshdtzEijzMIsz9BCjvEEWQg9rL/PBapB0iIBe4UKadKr6
uy3bBSwWHyPu1oJiO1GhbnqDSyRnu3N3GbOlCyXNqZetyFbrvOIm0PEkxmzN48lB
ilkjLPyGQIZOuiIsnwTUHHFgns/RlznrCyvhJT7WOb3Fq/E1xL6/lGxgw2L+cTj0
VBqY9Oh4FhDLfFZ/plltQ1hTBwzcCmzpx8jU/Qf5BnC9lT3huvRjY6L+LeqxOQo0
5DsyrXfJx7CJ03+OUWGNgpovYa6t6msVH7CEyjsJV7GmlY+YaqzT7yGKsSdg+cLP
itLJexIlFqKZCIxW8Q2ho9qFUJ5N9g6aM5rB5un+QffdBTEC8AJf3oIpY14WjPx0
uVuywmZaCRijiC5RvI/hL4TB/We6WSz0eyQpRda4tl4fd0d8ZNhaabqJhdAGlkwl
ZXerxAPFQ3w/EUjWqAiy2kFXmkMoj4oYG3LBf+Nmx/LqE4RrdkfIRqmT7We+hrtD
zxd8PtLsuXXlE4ifXZ6ZsUmrK56cmWg9uuLDlA9+I3WQtJ4MHDQOzQxeXHdu9I6O
8XZ3319NECCuJoRT9r+9PWQRQB5h33vj0F+bdfJ1HA6LB/u74xsEbnsEq8foiVYj
5glFUz64C3cSVf7g3N1mtJ+NMk3onXjxmeVtcV6zDTBbr8hlrRk1KK2MVNnkRhPz
VeifNFbhH4QLA4RFwEZL3sC9IYQAA/8JG9ChTpcRCJj0YAAtTlU0v/Un6hnO11lg
98VuaIUuT36ra1UFCTNYXplFI2bif6FEm3FwTu6lNncRrEqkxOAzD5pnPSwcxCN+
VwJmzqmd1W90Mjv6IMVz5Y3ep/eN73FpRsLEgyPFfyYZbj1EbkHc/l7BTbFHjZwR
xp/BX+5wzPGmq5g5MTGkPflPhoinfdsGOUgkw6kOhRRpFBCgOQWVfVl3Bxy/8LX9
0UvBPG080n+CZdjXMYBBfmHcW5T3UMn95AuB4+jXYMVfyVOO9tjjfLJqmZPoi6GW
CZjEXQ9OvKHSNH5SPxS9Ai2DpJNNo0AtgyTRqGelaI8ZWn9okSPNF47rbpwJ/82I
VjiJv9LYGv85lueRUxNOL57D+nsuRrBhbI2m/y8alL3GhxtTsniNBA66p4WVgmcR
qHLMC9JsYtLV5tk7Aus0afBQ6/pgxybLZ1CVRNNAx9nrMjH+S9r6tf3v1Zu8GWgB
gi8Szl92RMuxO1fov5ynQxNP68ohKygbLvsNU6Q3amhqWcvvU37RMtBfVw5u/WhA
C/pY4kTecm2mSOPELu69XEUrk+J2EmUnh/BrgoCPTNkItLH119YKiyXVi0Ojm8w+
XpRIWyGv06UkF50Fjh3rhO1Em0/AaxcFI3Pqgy9x2fmxNdWY+D9EWS7suzA2M1PF
/fuCDq7jVTdc2IZXR9D07UxFxltLtBhQh3xbx/ZLuXH6je3Pavod8oGnBDGhR+8f
/8csn8bCUFg7dR/8tmEU1/j1XP+wjh0CfN19lAFl7TGBYH1/eYZZBsULOExdyTs7
+6CaIClyDV+RBpqKc6CGKlQSMUB7yVwqSCK78bcLxBh4pjt0HP3mwwPKuTtwgH5Z
ikAkBRd8yISsdWhnGBcfYKMsNQNC/b//NHjp8fNDG8HPNPSAiNtqfrENVAsW6tL8
318oMPevjduJagf9pSU+JZRmOkehgNL5lWvelyTo51SlzSJ8i+R/Gv2QAWX4aFKK
PDCQ429Nqufjos8O1BYPb2n04k5IcFY6AiZLP4hROAlZyWU30vmQ6Q1STc1dT/j8
Idaej2lGmMEIGBRP1MjHXEmzSP3u6eCnGFM38aHRzYeoLdZeZrd0o/7RWYVsTmxc
7vTq5IggRAYIJmbQ0Ch4Z0iXRimCgcMlZ2Bo7hMZfCe4uIAMXcH2xuxjASFhiZRd
1D7mwmQhAwafcj+fr+6zN/UinIyEpc4mt+LDnjsEwAmk/JgaFwcX0BdfbGnQeWeV
jfhNNQfbIXKkF6HOZqWiKyYZvD+BLCXMu9dWNxYS0oV8OX302wois/EkHzgOmWXx
osKntCSyTYJ+MwzGxuoE79fgotrXCveaGfhjxnFy+OAs2xJsgx6lJFG3iMk+YsYF
5m4rhdBfEajSs5uCfVHcjrdOUwOLvfna1mOCnT7S4prAwR+NCuOasIgencHHUCO4
ejmYZZ8fudljudqIcjjdjXC1pCHGA2vCl9rjtv0/ObNZPpknEjfrYYlsjlN5Ws8r
Yk+4iokCci7+NcTnFPjspcEd3i2RBpP/b8uR8OaIuBdfXJ/+T10u0NLT9PAc1wfa
M3jPPvaTfzhFKzaUASTyOHHpWn+NXCyAhgsjUc5ettDg9mVolZVVZc3HWZsz5A8k
I0yOfmRbi8p50p6PFqB7d7klL3efA3tTPArw3ewTbtxSJGThmsgjbB1NyB/HtW6B
vCDWgIGusFx6+K5vZQBnTUC+DcjYOEvxjMmjPU8Mxy8cH65MqUg7Hn/thqhT/mhF
eyXQsXIVlmicQdgr0yyVNyO2ueya0+jF9fkaF8HKkubsHnWbHtYb8pZALdqdbeet
AE7hdlg+c1KJr26APX9HiQlP6PMuq5fOQeW41pAGOxoGhR3TMJpDAJ+kJd9E14Is
ssyhh/uiJPtLP5uvc8UZXZQgijvcivOyjoiZa/VqTPUhwMu4lSMRtoudaOGh2nna
ixTgzK9KuH011zoysIKJZpKhtefqNC3b/f5TveQH9h5fd8Xp1EhsOuSJ+kbsrJI2
VH2YrHkPq6KPnTgO1px8Y2Rf+zOCQIplt+BLC2Snhg0RmdyXwCZ8jKaxkZR66Rgi
HiwmjXFz/05lgzb9YV3ONtOH6l8F15N7kQ+CKrMEMakdylMEpxa/tcggmB3XUVi+
fwdspENQLzM8/LZSvNND8Dd8KM7aLisStOZG4IvB29ndCoXcUEwYDRAsfe4aCj88
nys9hZx7s13Elb8CoGwi6audidBTvx75hxzY0tk6qcviHivGbh1OZ9uPTNxNiGJ4
FpvS8uRi+hGZOvp7hWDazSD+JLOpLDX9Fx1KpS/ZFDpTPTNYPIeNEyLDAlvs9FVa
DN0IMH4CzZvLjaP2Te6TBWSma93fXEE3aLCOly+PZpssOR5+t5jwg+VPZhWnQtMZ
7lHyrMpyt5+/YL3r8ZLEEvG2rAxjBfBHi0Yg1sVZx+ky78uDQyuRlQi9pqMqS4RF
0rL02fEb7PiRV1zqqP4QFy7raaEJmloWtN/qezp+wSVJkEkG0LECpmyYGnktjw45
aqt6TYuTXXQ0g2fWypwKg4LHnuox2ufpIpcm+LWucCA4D98dbDF1G7W/ITU4n9RF
dRJICVcuLY2O+5s0G5um4zV/Zl6tZkg5Um8fZbna4Cuiq2vsmbNbBOh4HsqCIkf3
uQtVHN/QMUHUxFJsRbm93XPVX3hCIjrw0kTDuLgJXGJRsmz2mK9RSGjL7qk3TE+Y
5XEc26Kz86k148cLy3kQEdDJS4ZWcrXkA3fQdf+mcIspc1K0wYztR/7qK4AOwatY
owKj1IeAHGSUVI69RDtXIJdLa/kL5/Pb4OhQV9iYX2VUtXqG7x5eEsPCEv7uv4Bx
YEAlG53Vv55uZZ5vgk0Xa29HxNKLKW15QNzOvcZvvdUppP2IHlJ3c58mgVi5ngxo
YmRdQCi8IJAKCoDU+YludHPX/HqNWDKu9Vk2/DRpxB9WCHfbCLNfxfH2AhIsOV3s
QiL14ujxrlOMfwASfQ1bBFHpM8Jjtzp1loPyRa0SinzjZkMbyGI2VcZWBqfbl3c5
ECXp9qfsAUzXi76t4kZN4UZdiRdBJPrNZToRRFIbAuMs6lZPeLzTqPAVcp93DLcX
+/Lc+8dwduoVNGbdvtvabh255o2uUxqKWQOrpMKo96KaM0IdqXDay/jYTvhs3cXX
IcDnVFotlLsUtQSJYCOnPWfk2+WJc18gruWJcXpnEIRVPBXv0sVP1+xzRpTklhiQ
hYMJANIPzZ5ImICqqJBNi6p+cB1fbaUujYe+tCtTlZZIsWL7Epy7PY79p1FNWXAs
EyI/njr5hOn+G86beBNz2+R6Mlih06DoksO7t2YjOmR7xFP4SX6OSYLrNaKwLzSq
CpZKpvlr9ybCyKZWcyBJZkLywEvZ/9Te7kZKLZfW99//V1Y1RrztabBOcrzJX6Ts
taHARvm7QrtX/08CmvOvulEHwb6nGBIIKHXXT6wRNQ7+eGSorhulsWDGTL1FO8XV
vpu2z07DHmWfcKLu+SGiYn/3SNS5XafxaE+yqzjjQZNEdpsmguj00O2lGZ3mKg7k
f4mIJ9HZ1kKdY/czdo1cyBsfn7K+oBmNwqm3PyUu4xKFiAlOaffZnyg0jmTTp2+v
vljqohsHwgMt090HQKwQUMmt887LoSWF/oiWA3tRndRsB/B3u4AAFvGrp/bO4COt
mnW84Oi4FvlJAUdoC7Gos2BKrtrTu2FaV1eOm4SvAAyebBuVKvPk+uYmpYIuzPRc
JPUfcYysR7pPHc0PnFdhNz+q1AO5Amu+35cYOgiLeixKb8s44RvUPi38VulY9o4e
9M2AEGk3cm6mAJP6IvMz4ZDnnpUy1Sx82BeuNHHEtwPwjk/SPD3MtQ11AEGQaQCs
et3P6brs/bw9ZUi04FT2eAwvJiyZHcFABlGLXM254SOVJGthryMQIBiBJCf0WYFW
Za/Y7Di2K+NrxtkwyBCl3JaJSLHExzpBi0c4vTm5HYzuO9TLeG9j77UZbKIdFH/U
MH5HjxPX7oPf18lP+GadfTodYNwiSSVob0WCpkVGX48TWxHhgeM/PvlNfa2Z1gO3
R+zfS6tCj/ftXW75fHqS8sVL6rNbMj4jkYHfrYNbVSgekFelbL42Pe05IBI7zm6k
BALl8IAf+FBM8Mhc/wXUg/9Pfi8bFhtS08dyr2uOULmVGScVcxSQKoZmmla/mX89
5vArF6zSQU1xx5t3GoGFlOOk8z15m8aEjk6DK72QzyCbV9w9+f+lS/en3WEUJsaY
GSHOwKbDl2bTI/jTGNTGep+YeYgVouiDyuwqOdKmId6E5yS8b/VZ/cq2eB41gi1M
wSqVQ5Qi6+sGo8vWw4sja5pM955KHz6B5fHJo1qyFd0cdIgdpI3uStgB9PNszZ57
xGzd2bU52Pl3K2RVAz+ZiIGsL40t5YMhk/+6zDjUJW5O+SLfKvytCjIs5oWYY2Jy
omIPS7DyaijYTMb/vz0YnZMWWg602vhqcKIvN9sAObmORz8VaC/7Fl++joVjgn+M
g+TBQfVfkK9HBmNsxKr00ySt6PS0qnYjdy8ZE86L9CbDiCpPnRnkgRYKvT9vAzAr
bd97Xiqio1rC+Xg9Zu1H5H2m3/QDOj1rMsaTi7mvOvXOl0eOgLeRKvwt16RD6RYZ
5lzeFuzJqcZXDBNA9HtIpypC4vh1erzvj9ooGqTYLSMGxlLhDl8uVVEGH52JClUd
2WoxMjLXJ6bhqVSuxFXVKXCkcHq2AT2RlrZNW98P4H4HEun138P1DyEUei9weCTr
a7vQKkhC3onf2Dlau5ssSgwMqMOmalvqjtgzD4uV+AVkvDtYeYOzOKOcJUx98zzO
68R67Pz2p372lxMrPWVJaN4WtfKIfwuiDFQ3LfKGuyg/iG5NIJLjuLhHlUqekeSG
15nOeLcHem5IA4suG2IN4uIz51eQ2S1mAuIh+5vFndzKHuaDgDsts1uHeUF/vt2f
IOhWBDiuWttw9EUqpAPnUCq2ZlKuGPtojhfGaBuPHBILpxXr7z/JMnbvayQatGaD
gXhREokMyudfLsjpPsPD3+MmOfN+lvCO7mX12n2TA1OADtnd/uhKuji7bb8Nx0vh
96kkYsctXNr2d6Sq/4Vx727KlhKBpcDkWZQGL0TufsEzkD2/KTunIVKCofSmUvkt
n1AOe8cbOXD7CPvORyqYpAreMUOzrVhDUFqjVBwWzk9KiKYMsxHAm5Ni3byTULn5
MOV7YPKYGCANUCyvcW+pGRQogwoHDUe+2J43RehUg/1I9lNWCnNgmZogVHGVSJrJ
MH0/J/2RtOt4JyrlKB0/efw+kWpq/2UvXpxwjGByWd/xeHpMzxS2jmeYvfvA7hjy
WOw36HXGojDDUkt0bNx4qZPmyMtrXjj3f1I1FPPFaGdoFEU1z7b7cO6ZVlp8w77e
HRWr/o+UfOgRgYN8ylrFG1XIXipk6poo40BMz3cFNWQ27lM3ogC196bk7Lk6zVSC
7XSFAe7z1AYnxB90C1QmyuTq/JsWjYWvD7Omdpx7nmgpCH+eEFauBLMWigu4xCQz
Tl5+rWq1+lARLXq20ADxzBKGCm4FKFNhMYjvfPLHVoPu9fgEbXCWl0Kr46YaEyxT
HsY7VfE0znfR/9wDawbUchn/rGQbEBYJZfJh5SB/Xv2iyOj0DI0e16BcYhaOaUiz
+Ay6PIyAyihUiJXBIOz70kLUNHQdJNNIVDKnB/VL7L6miTsv7EOLM/ctL6iicBbz
QEbqxU4QgW9jrg+vEOufB+BeFISv+mEEE1bpsxw1jfz79l/q0YKJcdWJ+uhyrGhN
ZdkcdTxaAQvxK4Q86GOFxbjdtHSeQcxTi08NKpqaVCNHh0ebzD5dyGxtAXt6F51J
8Mvsy8wPsdBXA3wh4W6SG18MWToWLyZ0ZeoaUvLvJoTGIbSilWPOMg07qjRR53Xc
NqH0Up+3rEa6AUZosXW8CaMIXCx+dpcyY8jucR+FLOVsSvwrlB+NTE/+c58ep+WU
lWVdCMp5Dx7MVlvjxdF4zZACwU6qblaGo7s+UUM/lkbANXnRnqOII6UO2vHyP9ZP
AJQ5wYefKSshzNBDWbppElnxg7Wm+2Fh8RkcXxHi/fOKL3l+2T9R0rV07QNlsoeQ
grYrvnhtHyc77aoXGBNynnx/gOrApzakv3CtCinNUxgrBl9jpl3h+kEc4cPrVTm1
5thB1+SdN9CDld1LTMbDqbJ2jHMTqWqilSSC8PnocQe/C8dNqEGu58JWD9YejV+D
hFhJGSNc+orGCDqqudd7GkVuTFSfKGz3hegqK5JIkcSnQPSB+LGUZxlHPtMCA1vM
CFymlJFjSszdN4dNHr/9Tlat76AMk5NzivIE9yRM6PtE3r9Eho8jWZgYYzZQuCzV
6qpen9sOvwf05keoLlledHu4mq/W58Q9U11YOsZSUE5BzxxCGS5F4zDWHv3BRSju
Sq+yraEqh7UdOowiR9HuurAxDHoOqBEaBFo0xWyllEjYINUBgaHmhs3Jxx/RiwqX
5+G8/FIY35BZp2+zHjDwPJsQv+zUv1nyDF78D8ykwcX88xevDeSOELbTIctWzAbT
d/n/yt2ltVQH6RAkbDG6arIglpWOEdREGfeYQCQaPi4TD5iRm25FTxKFbGuNfy2h
5ZFR4vjIy2B8MaqbEscPS4HVf0+Lht1rKaVnbaXEpLKPoaPrdT0pDjoNIs7LjYDs
OZbYZhDBeu9212kiU/qXShXhd+vLA10WHFbQrHwfpNlvu20kgHrwofvuLoT/aThI
wBxWkMq/wHBQQ3T8VYJofvA3BKobKnOhJVQ7H3Z1ZSapE5C2Gwh7ho7s9uXiONcd
J8/6+7agMb+Uy0X13gxm1r4bIrndH3aOTP+a8Ta+r45OM+dUZwYsjeOtjW4rurhI
teSw5gwdLoq45KW39AqNdo3j9YUagWZe0qh3xClRJkIeWWB4FjOeTryKLqAOTPZH
vhW6EOL3ogzOdCQse9WJV6Y1ghmZv/fQEX9B20FOlMgAtMxlGlrBA0LVk0oE2qgQ
N4GbUNzA62H8QzfBUVkNM+CHuMLp50aUei6Ir2NoeAtq4ihwuyKNNcFynpSLLL6L
2obR83GOeG6/etlk1JU30MyPeFIaEkxEngSPN4uClClFDB89X0RV7ixPif6ovXVR
uUx6YLBWTrDB6gMmPREi3TyepxBCaIfsBQWolaIm9lFX3XXOlqZt0BHzObAvGDew
voxDFEbuP3Ep0pDyDQ0HuqUwAAx+053eEWqCAAtQ2QBbTHm6GHz/nmIJAvtnVmxB
HqIvI/pH2Muuejh6j/j0uwMYhwUxrj0qbUkb4HnLjGYBPuXbWCs/cUuT9QZPEDiB
QdPhikRLcIRPc4KTXUn0iaBaRD6/veR4HEvL11PUDeoRbwqrwo7PmnQin+mxdm/A
o48umFwqj2wo7nsHfWEUeZ0G/GeL8LltOT9Bk3hxq/3UCs9XaBfvuo+phPSh8Tua
tahP6M0Mj55jUxN3aosm9yhC31wGotGSv4ss58rU59MRtRj8N2Wq1XUa47vRNtwy
ToBViM84AzVQOuoqS/Ryxl/vXOgrjntmqdq6oe4YUx2DDMHrC3fZdLfhfS0EJfxq
DK1uXzaOxchQ4iQwXKOV0ATkIzODTh+06hlHtP0aFJS9o90wvkqW2MykpPMnuoN5
zufYB9n0pC3AuRayf/93ixKHyszhbNCosDg3oZsu4e60a0D/PVpQS5lFi3vD7ULV
sI8fUYDHnvbdpASBTK7N+CCD5oHVUg/VIq/xuKWVW1v4JTlgfOLXoDMY2YcBXzMQ
DNlnQngZ2g+n1GuH2lelN8nIgc2DjAjMRn0IPM91WdE+WECkfz2ISFTEvFUCs9ze
JEWEK1c3DOUt7mIgNi0XPaz7nUnyy4ZBo3pOI+/SvUwcFuyV/EdxKiWHxNYR3ACk
OlNum+JX2TGIIL6ftRBs0eBI3HKAfhLURBvO3b3vn/WPZpO2VoRCwbJv8cF5sPlU
sFMRyR0SO+W352ZHBfyEkWUFj3WEM2jdYslIfifZnMafGhwqs3pyrT96VmHkP+xB
O/INwgCic3MfiwhzpAccuUwitbo5HTZls9rtCjwhhcLcW4x9LfO5vvq3FhOYIcTf
bN5OdK4laSKpA+qsMN6aOQ1c24SrZ7VT7QTeFGWnXE4Ogd+L5xPnZJmC3lotfuje
WzQ+hG5WGK5TmE+HA5SJph9iazKa/hQtDg9+I7OW7QKjaG2trU8Bg9Qi1cfVUr1q
cSPX43YqHK6E4AKDBElARnxRz+JoBAHVJdMPxZqGXX4LBk5sxXyOM+AMhQ/Eg9qd
YGuDAb3lu/MJvpdwBkYic6Vs2ZXyjVX5QzvNSRNDxwPTJI8fJSYB89KpBR0ZyMnz
wNuZ6Nm1gPct2zdFoAyxwBKPvGHk/pAFyC+SvSfUYkV1f9j11L5k4JDJuTpmSrRL
sI6m22JBHBg78Z6EZKeb6FS9ShRMHZFftV+qH4uFAsazaQIsP5wt51GcWpFnMewq
B6xTRVIiA6B/iQTord9ptC0fyW3AZHWb6/WLMY2Jil2X3mU5DunyIDnIK2p8K2zb
juGnrPTt8d/yuR5abtVMeLiAVi1VJY2UVXCFtfTnltiwxzTv5cYQz5CUu/EECtuy
6xswxk5Yh7FLlgNs+2UiSdFaz+2ymaZ1Rp5vP/z7lk6hl2+zrTGn8HMvUa0Yk1IZ
vbIYJeD+qmSu3nPotHEz+362Fr2JnONWYyFQzFgRl1jAYBWpDwKnTtLLtr3lSoVy
GNhXmvGk3eBbEgxoW6UzS2BeLRnOoFGceTnfz+xyldE7nld5Kj1kSdX/YOd08/os
BlqxrvIkwJiPDQC3DCI0/vckdTLEjeH4QT8zvLIYV84Az/fMFX3kIkFF95dggRHz
iflFCFC1JiTd3ODHZTlMGfItIsknFbzZkRwuRcga1YUmu1vBrJ4OQg8dZpqToZGq
zG4nliF1XU/y9LPjyOhkp78TmlqplX+bXd4Gfcyo88QejIeG1mPVo4OlgVg8h2Z1
bETTExcHjzfKVJucY0kJGPPKn7j6P7d6oFFCPq111Kuy0JpfLoHzI+WROYrqz4E6
DP+rsp4igoBFpITWGJNNCQ==
`pragma protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���??С�M�4�63�M+�����ӭ��Ni;�Ig�Rs�8aр�s��RŞ@y]�""����s��Q���f�|����a����J0��F}(^��?��T��j<R��X�G��ۖ�Ŗ�t��f��[Y�!�+�F��|q��7��[M��~�@��hD���Ʋ�͡�??5"��b8��Q|*L�^��}y4�.��Y������q�>#z���at�D�bU޻=���}x��94��zH�f�[�̍��_Hߺ�ޯ�̚�©����s�3`Y���W�0Q�ԍ���?�+�FCɺ�7/��:Z���Vm�E$��)���oE�"DA)��aY/V7#��$���oh$��:�,p	ꙷ4��b����]�8,� �Ŕ�O�Tn6��"H��o�;8|�( �Sj0$1����������&.����Q����[�r��^�@lI�`�h��ͺ̀	m�-��N9�NOK)�Fld�������Y��AA�M��f���]�X�726�87c�F9��Y�\v�ͥ�*���ů	��)����u���Ye��@����"�-t*:��ޠQJ����}���\�[��j]�V��3y��~�����w�P���S��^�8R�x]�n|��1E����۵Ԩ���C�ǆT��W�V�;'��m8�mЕ�/U�.6�\�\k��LŽ+��t�<FD�W�� �
�O�`��#�,�c�(��>ʧ�8,�.��T�Q�(}�v[D�H����vK7R��ݜR�AT���ǳ��!aC�l�h�X���l�W���\������:E_�@E�z�'��9�i���l3�T�jD/�{O��o��x(.����)�n&$k��`��34�¸�b<Wq���`'㌌�f!��6��H��ƴ��M�ٚ)�(X�)3�|P��p��&_2���4 �4����5p&OaZ&�~�����N���(�2���B@��J�ʼwl0�yV�
E#��;�#7`�ĝ�TX�ճ�xpO���lTWl�0�����l�%��G������� ���;���x~,�z�J��(kt�'�����uO���o"OFi5.�����}��v��Y�l�7���3��e2�rDz�����Q��~,/%n��c͠K��V�+��	乒b��߸A�~]"���#��Y�-�#�b}ReI�OntYXL���*�_��,綥�E �\왽x�訌Ь�SU��]!j!�p���%!|��П�6#ڜ<Y1+�r�����������H�.�aU����pU���*�� E˹=}i8�Q���r���]7_�cI(>�#g�	���Rٍ����5y!X��O�Sе'�O~MfҐ)�����	*���>�������Fc~�Ow%�=�`��Ni#����D���c%�������UXLP�U/@�a_{U����4�U^��ANنf%n�|g9�`a��͸�"6�cqRz����Q��X��~�ý4T������muθ%�E���,���qz�^�I{n/�/�<T��P	婶y�n*_azZ�
yn��E]}&,`�f3����N?/��Կax� �^>�<0���m�X�+t�3����Lv6�F��}ڛ�@���F<u��#޷�˰ �+��ּ������q%��#N�ق�k�`VW]и{=��N�t�o۾~*��@^^� �+�l��٪�l����(,�eZ�E�)������ (z�h0^��\��a<Z�p����lEbX5��LR��X�h�/�`������p�s�E�(6z�H����"��IqI�Q�~��^qÏ �2V,�����Bx����#�n��5Sf��	;�:��M��5y���z�l��3��3��I�v6ʕ���u�!]M��;�}���S�͑�����hC~��՗���E����:kǡ��Ļ}RDt�j\�#ǳ)�D���BX��;J3P[��Q_����e��'6��9s2�]��<��U�(�JK���~��u7.�
����7������ڟ]5�8�/�9��?&"��J�G�C��r��Ez��s�z��3�Ps���i�\(̸��99�R	�iӞ^��6�)�<��6�bf��ɑ7I����E!Pj�B6d��J��M���'���/���������F�^e� NB֗��#~��REJ������A���i�#�z�:��`{�����D�����ue����F
���t��Fy���s�Z0�B.����C6��(�Uu"5b��C�g��v K<E�x���� ��9@�l���
 �ߐ�4`]?J�Ҧ�X��L�:

ŵ-�#�q ��:K��](0��Vj�C�)��9u���Zv��s�B�zy�NT3�M^cRJ��M���[��ɤɇ�T�I��w��(���D�Vr�~\��đ�N"���=�K�ǹ��b�������z�L� D�x��+8�q���Ԡ�������%	Ц�1p3�a�OTSU�0ཱྀ��#Lv	�5��J`�}�)ti7[�����~8-I����)�6��Iӝ3it۸Fu\p�*�*86Ŧ����Q���k�ג��޴,������2-D=^C�$��$���ZN��Z���O 0��r�M4�ZdI6��� �IS�<�(I�U<m���ʙ����rL�cn�С���ϖ;&ڹ�w˭����;��E�-���H�s�t@v�J6��eoI&{� �m��yӿ̪��T��L`u�I4�S�!���9�%��Y�c�]
�/��� �NO �n��c�pQ�6<2��tpS��`�*�q�&��!:���J��0�O��y�[�	0/V��+�����)pZ	�+ם����������7��{8&�*�3�3�k\�AF���6:"9V� bcԖ	4߿+#jO@�r��t�"����M@Ⱦi	rL�ŉ����&[�Α,O6�R��c���?g5�,�t����;�U��=��Ң;0����Vƣ�)�a&�J�	`'4WI�uv�D|d�X���O&���,��{[U�Z�/��WU|A�b\���+p�Dc
{l�"�#�=S 	�Cέ~�Q@q��U҂_��,��T�S�w�x��9� &�2�xO���$�­J)���v����:��g���͈���{q�x��u����X�\*Z�:?������nnÕޢ���W_�Ja]j�_ol}�{T�=3^"���C��s�PK��S����e��U��3~s��Q�",�U��k��z���>ZI'���ٝ���Ư��h ~9������,A:�K�]:ϪU�x(��C�X���[`���es	�?�r"�]{���s�A��~�9��ʆ	+��B/8�*(��BNc0F�9X�[�J�s��Ü��Ud�@\�v���/�\u�o�����p+މȶ����^�?�P�d.'�a��v�,)'�2%�l�AV��Nٰ����3���Q�9���Y�����S_S�X��O�H`[�'�qsX౜⩧�_	�fZ�u�X
��U%,y�]j�V֘�|c�!���&����ʘ��N�Ǫ�iS*�h�r����V�0K�� �"�a���lu;�M�˟��8���Vpf��m��uE����hr7t망'�g�\M�`��G 2�/�.�zwy�C� :׍=�������ym2�ߌv�WROgx�M�9�|Y���S������ 	����׆�J�n ��6����`��/�b-ý/F�.I_��3�ghR��ؐO-���M�9x�1;�A�l�+:b�Y!���Ҥ��N��
YH��*!���I���gw ��a�@�"q��=�[�2ISY��w��@�=V��_(��kC0���Y8����e��i��_Ž�N���bGy���Ό3S�75������p1�-=�t�;_4��A#xb'�?nLO��>צۣ� 	ǽ�.�7`;o<~K	�������k�w?�y���C]��B�A���F��H�j��z�iU�^<����8�*J�R���]�I���>��^S�h��fe_�˼*Yl��mM $�x%�.�Ȓ�I�J�-sUɕWІ��Q\��'rpu�Ya����;5|�=����6k�����U�W�9^����	H�*9��g��/���Z^0�UCe9��W���=��w2�%|+(��[�zU�M��W褗�v����R��D�|�x�g��御6vw#X���z���?�ƢY@��ܯ��3�ӰH�A˂���,K��oJ�s�	��y�� � -$b�38��g*����Ǡ�Tն>t�Yw�8��?��&���غ�O�{��]�4��s��P���zk!iOF�Sw�B�{\��f����<hٟY����]�e�@F�y���O�]�-K)�i�Ŏb�����r��x����st/c�!�0��q�&�6v�J.�(ڊ�ge�+��������֣�$�6���`/��%�8@28�V�ݧ~�fU�G-?��
AԄ�QX�`U�bt�j�4sP���=�̀!��S�ڤ���#�l�뺉cpT<�A���WQV�]��ᤋ�������@ޗq�8���%#b��r�a+I�Y�¦n�)־������R��A����h�o旝�tٱ?а^��]J�s��I��������9��Y2�)�����ɠ%� ���_f��P���Y�pճ�ҜQ�3�syڗ^R�!;G�Y%�iL)*��{k*t����&2�z��M��چ������+����.ވ[��D�԰/0Ѩ0�4��Y������98�Rw�㚝�!�z���dF��TbC�LPG�r����H��>���i`�S�u����yr���8�i3�PE,�0U6!�ʋ��ȟ4��D�C&��>�^�'��������&��I�]	uA6S-��8�B	�ݰu���y�ZF�P��L���%L	�!�Ɣ-�L��Ey���kl�G��HsR�Ϻ'���Oqi���?9����f��NZ�t�Z���v"��ֽ�h�o�����u�;¤���B��fC4j��ʚ���lB�@���������8�x��l~w�+�׳:X�\�=���Fp�-@lx��#�{����r:̷`�)!6(Fp�e�c��'И��h��ٍR���hl�t՜�>��*VΆ8n{Xn:�S�F�Z���! e�?Ky�$�N #���I������ ���t��0��D0��_���b�T�����~�'G�t��+��6�w��D��T�Y�Y�B�FK�.�ǯ0�>9�����v��]�f;�rC2�}���O,r�&�,]^��E!Y�r�o��@q�4�y�T��{�ֽ�V�^+LGa����bǻT]�.��$m��a4��P8����O�s�w�@7�*����Zi�-��FCw}!�a��$�rp�l�w�L�1���eQ<��$�	�-֤���:h�Q��p3E�	�/�ÿT�����@�����5ޥ���·/8��x�4�ae��������u~v�N'�ʾ�}��w�cʍ�oW4�dPj��)�S���^1/d�p��y�S4-K�F-F����-�G�#���y:�^uј%'�����C�i����]v�W�g`�h��2Wo�Ry�o�������g���0�	1�d`���X������k� Ŝ
�A�� ��[ ���Xa�z�{��s" �]׊�-<o�cUk9�Sd�pj4Zf�beMS���hR	��>��c�pi�
���Bxܡ�N�v���X��Ɇ͖�fY��|���H:e���5���iK\.�I	[3Xc��U������o�34�]+
�X����$���śV�2A,�MDI�vH�j����k���0̰1V����ߙ���Aʴ�T��tO�7ܷ��u�h>����A�W�Pzp�6��b���{��|�~I��}d��t�[b�f*����i9[x�.�8;����`p;�*�g����zc���=��gI�������6y��w���*��/��r��|�;��M�yP�?10)&{�K�gi*�S�X���� <�	j�GƉ�!+34���:ݨHN�⒮�7YZUm���_<$�-�x,��k�"b�t��a�`!�K�#<6h�����Z �s6h{��27�j����g��E�z�5�{�f&΍��������F�
�%&��"Y��O5m-�����$�<{y�Cr���=HA�vα&�\	�|�K�9�vO�Q�M@����}���s3�r&���W�]\,{��j�6}�c�e�rmM��&�-��UoW�����E��Ŗ·�m��ÿI�8[G#�}ȭ󭻺wTG;�􀣅��Vu>P�Q��	:�rE_Wv���)s �}'R�)�,�i��`P�������4ʇ�>�:6��j�x�������)	�(��]�z��Ђ��2Ņ�Zf����eG�R
K�R �+�x��_��Tf�t����_���O�C���3����\i�_����ۼ��w4��b�gtcʯk��зb;%��Xsd��R�!W�dcZ����usɌ����ܙi���wx�J�0FG1Q?�a�#.���9SY<0�'dʋ�9���!U�r4�q���"\�#~OtnXT�I�����.(Ǧq���0N�_ʲ(B���������E��:��f2�ٙ;�m*㙸Yۚ3YYt�ʚ�o�^�[�L]�#���X��ʽJ���s�R8�f�7rQ����)C�l�Иb<FG���8>93U~�]����5��������3S�L���g�aj�>�Ħt���˙��������"A@`1��XS�b4g��[⳼�f���u�ʊ�����IC�PE߅���Z~���s��}�ㇰ�H<.K�o�"(�±
VM���S��sv�1q�
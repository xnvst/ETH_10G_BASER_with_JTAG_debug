// jtag_system.v

// Generated using ACDS version 14.0 205 at 2014.11.09.00:39:26

`timescale 1 ps / 1 ps
module jtag_system (
		input  wire        clk_clk,                       //             clk.clk
		input  wire        reset_reset_n,                 //           reset.reset_n
		output wire        resetrequest_reset,            //    resetrequest.reset
		input  wire        mm_bridge_s0_m0_waitrequest,   // mm_bridge_s0_m0.waitrequest
		input  wire [31:0] mm_bridge_s0_m0_readdata,      //                .readdata
		input  wire        mm_bridge_s0_m0_readdatavalid, //                .readdatavalid
		output wire [3:0]  mm_bridge_s0_m0_burstcount,    //                .burstcount
		output wire [31:0] mm_bridge_s0_m0_writedata,     //                .writedata
		output wire [23:0] mm_bridge_s0_m0_address,       //                .address
		output wire        mm_bridge_s0_m0_write,         //                .write
		output wire        mm_bridge_s0_m0_read,          //                .read
		output wire [3:0]  mm_bridge_s0_m0_byteenable,    //                .byteenable
		output wire        mm_bridge_s0_m0_debugaccess,   //                .debugaccess
		input  wire        mm_bridge_s2_m0_waitrequest,   // mm_bridge_s2_m0.waitrequest
		input  wire [31:0] mm_bridge_s2_m0_readdata,      //                .readdata
		input  wire        mm_bridge_s2_m0_readdatavalid, //                .readdatavalid
		output wire [3:0]  mm_bridge_s2_m0_burstcount,    //                .burstcount
		output wire [31:0] mm_bridge_s2_m0_writedata,     //                .writedata
		output wire [17:0] mm_bridge_s2_m0_address,       //                .address
		output wire        mm_bridge_s2_m0_write,         //                .write
		output wire        mm_bridge_s2_m0_read,          //                .read
		output wire [3:0]  mm_bridge_s2_m0_byteenable,    //                .byteenable
		output wire        mm_bridge_s2_m0_debugaccess,   //                .debugaccess
		input  wire        mm_bridge_s3_m0_waitrequest,   // mm_bridge_s3_m0.waitrequest
		input  wire [31:0] mm_bridge_s3_m0_readdata,      //                .readdata
		input  wire        mm_bridge_s3_m0_readdatavalid, //                .readdatavalid
		output wire [3:0]  mm_bridge_s3_m0_burstcount,    //                .burstcount
		output wire [31:0] mm_bridge_s3_m0_writedata,     //                .writedata
		output wire [23:0] mm_bridge_s3_m0_address,       //                .address
		output wire        mm_bridge_s3_m0_write,         //                .write
		output wire        mm_bridge_s3_m0_read,          //                .read
		output wire [3:0]  mm_bridge_s3_m0_byteenable,    //                .byteenable
		output wire        mm_bridge_s3_m0_debugaccess,   //                .debugaccess
		input  wire        mm_bridge_s1_m0_waitrequest,   // mm_bridge_s1_m0.waitrequest
		input  wire [31:0] mm_bridge_s1_m0_readdata,      //                .readdata
		input  wire        mm_bridge_s1_m0_readdatavalid, //                .readdatavalid
		output wire [3:0]  mm_bridge_s1_m0_burstcount,    //                .burstcount
		output wire [31:0] mm_bridge_s1_m0_writedata,     //                .writedata
		output wire [17:0] mm_bridge_s1_m0_address,       //                .address
		output wire        mm_bridge_s1_m0_write,         //                .write
		output wire        mm_bridge_s1_m0_read,          //                .read
		output wire [3:0]  mm_bridge_s1_m0_byteenable,    //                .byteenable
		output wire        mm_bridge_s1_m0_debugaccess,   //                .debugaccess
		input  wire        mm_bridge_s4_m0_waitrequest,   // mm_bridge_s4_m0.waitrequest
		input  wire [31:0] mm_bridge_s4_m0_readdata,      //                .readdata
		input  wire        mm_bridge_s4_m0_readdatavalid, //                .readdatavalid
		output wire [3:0]  mm_bridge_s4_m0_burstcount,    //                .burstcount
		output wire [31:0] mm_bridge_s4_m0_writedata,     //                .writedata
		output wire [17:0] mm_bridge_s4_m0_address,       //                .address
		output wire        mm_bridge_s4_m0_write,         //                .write
		output wire        mm_bridge_s4_m0_read,          //                .read
		output wire [3:0]  mm_bridge_s4_m0_byteenable,    //                .byteenable
		output wire        mm_bridge_s4_m0_debugaccess,   //                .debugaccess
		input  wire        mm_bridge_s5_m0_waitrequest,   // mm_bridge_s5_m0.waitrequest
		input  wire [31:0] mm_bridge_s5_m0_readdata,      //                .readdata
		input  wire        mm_bridge_s5_m0_readdatavalid, //                .readdatavalid
		output wire [3:0]  mm_bridge_s5_m0_burstcount,    //                .burstcount
		output wire [31:0] mm_bridge_s5_m0_writedata,     //                .writedata
		output wire [17:0] mm_bridge_s5_m0_address,       //                .address
		output wire        mm_bridge_s5_m0_write,         //                .write
		output wire        mm_bridge_s5_m0_read,          //                .read
		output wire [3:0]  mm_bridge_s5_m0_byteenable,    //                .byteenable
		output wire        mm_bridge_s5_m0_debugaccess,   //                .debugaccess
		input  wire        mm_bridge_s6_m0_waitrequest,   // mm_bridge_s6_m0.waitrequest
		input  wire [31:0] mm_bridge_s6_m0_readdata,      //                .readdata
		input  wire        mm_bridge_s6_m0_readdatavalid, //                .readdatavalid
		output wire [3:0]  mm_bridge_s6_m0_burstcount,    //                .burstcount
		output wire [31:0] mm_bridge_s6_m0_writedata,     //                .writedata
		output wire [17:0] mm_bridge_s6_m0_address,       //                .address
		output wire        mm_bridge_s6_m0_write,         //                .write
		output wire        mm_bridge_s6_m0_read,          //                .read
		output wire [3:0]  mm_bridge_s6_m0_byteenable,    //                .byteenable
		output wire        mm_bridge_s6_m0_debugaccess    //                .debugaccess
	);

	wire         jtag_master_master_waitrequest;                      // mm_interconnect_0:jtag_master_master_waitrequest -> jtag_master:master_waitrequest
	wire  [31:0] jtag_master_master_writedata;                        // jtag_master:master_writedata -> mm_interconnect_0:jtag_master_master_writedata
	wire  [31:0] jtag_master_master_address;                          // jtag_master:master_address -> mm_interconnect_0:jtag_master_master_address
	wire         jtag_master_master_write;                            // jtag_master:master_write -> mm_interconnect_0:jtag_master_master_write
	wire         jtag_master_master_read;                             // jtag_master:master_read -> mm_interconnect_0:jtag_master_master_read
	wire  [31:0] jtag_master_master_readdata;                         // mm_interconnect_0:jtag_master_master_readdata -> jtag_master:master_readdata
	wire   [3:0] jtag_master_master_byteenable;                       // jtag_master:master_byteenable -> mm_interconnect_0:jtag_master_master_byteenable
	wire         jtag_master_master_readdatavalid;                    // mm_interconnect_0:jtag_master_master_readdatavalid -> jtag_master:master_readdatavalid
	wire         mm_interconnect_0_mm_bridge_master_s0_waitrequest;   // mm_bridge_master:s0_waitrequest -> mm_interconnect_0:mm_bridge_master_s0_waitrequest
	wire   [3:0] mm_interconnect_0_mm_bridge_master_s0_burstcount;    // mm_interconnect_0:mm_bridge_master_s0_burstcount -> mm_bridge_master:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_bridge_master_s0_writedata;     // mm_interconnect_0:mm_bridge_master_s0_writedata -> mm_bridge_master:s0_writedata
	wire  [31:0] mm_interconnect_0_mm_bridge_master_s0_address;       // mm_interconnect_0:mm_bridge_master_s0_address -> mm_bridge_master:s0_address
	wire         mm_interconnect_0_mm_bridge_master_s0_write;         // mm_interconnect_0:mm_bridge_master_s0_write -> mm_bridge_master:s0_write
	wire         mm_interconnect_0_mm_bridge_master_s0_read;          // mm_interconnect_0:mm_bridge_master_s0_read -> mm_bridge_master:s0_read
	wire  [31:0] mm_interconnect_0_mm_bridge_master_s0_readdata;      // mm_bridge_master:s0_readdata -> mm_interconnect_0:mm_bridge_master_s0_readdata
	wire         mm_interconnect_0_mm_bridge_master_s0_debugaccess;   // mm_interconnect_0:mm_bridge_master_s0_debugaccess -> mm_bridge_master:s0_debugaccess
	wire         mm_interconnect_0_mm_bridge_master_s0_readdatavalid; // mm_bridge_master:s0_readdatavalid -> mm_interconnect_0:mm_bridge_master_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_mm_bridge_master_s0_byteenable;    // mm_interconnect_0:mm_bridge_master_s0_byteenable -> mm_bridge_master:s0_byteenable
	wire   [3:0] mm_bridge_master_m0_burstcount;                      // mm_bridge_master:m0_burstcount -> mm_interconnect_1:mm_bridge_master_m0_burstcount
	wire         mm_bridge_master_m0_waitrequest;                     // mm_interconnect_1:mm_bridge_master_m0_waitrequest -> mm_bridge_master:m0_waitrequest
	wire  [31:0] mm_bridge_master_m0_address;                         // mm_bridge_master:m0_address -> mm_interconnect_1:mm_bridge_master_m0_address
	wire  [31:0] mm_bridge_master_m0_writedata;                       // mm_bridge_master:m0_writedata -> mm_interconnect_1:mm_bridge_master_m0_writedata
	wire         mm_bridge_master_m0_write;                           // mm_bridge_master:m0_write -> mm_interconnect_1:mm_bridge_master_m0_write
	wire         mm_bridge_master_m0_read;                            // mm_bridge_master:m0_read -> mm_interconnect_1:mm_bridge_master_m0_read
	wire  [31:0] mm_bridge_master_m0_readdata;                        // mm_interconnect_1:mm_bridge_master_m0_readdata -> mm_bridge_master:m0_readdata
	wire         mm_bridge_master_m0_debugaccess;                     // mm_bridge_master:m0_debugaccess -> mm_interconnect_1:mm_bridge_master_m0_debugaccess
	wire   [3:0] mm_bridge_master_m0_byteenable;                      // mm_bridge_master:m0_byteenable -> mm_interconnect_1:mm_bridge_master_m0_byteenable
	wire         mm_bridge_master_m0_readdatavalid;                   // mm_interconnect_1:mm_bridge_master_m0_readdatavalid -> mm_bridge_master:m0_readdatavalid
	wire         mm_interconnect_1_mm_bridge_s0_s0_waitrequest;       // mm_bridge_s0:s0_waitrequest -> mm_interconnect_1:mm_bridge_s0_s0_waitrequest
	wire   [3:0] mm_interconnect_1_mm_bridge_s0_s0_burstcount;        // mm_interconnect_1:mm_bridge_s0_s0_burstcount -> mm_bridge_s0:s0_burstcount
	wire  [31:0] mm_interconnect_1_mm_bridge_s0_s0_writedata;         // mm_interconnect_1:mm_bridge_s0_s0_writedata -> mm_bridge_s0:s0_writedata
	wire  [23:0] mm_interconnect_1_mm_bridge_s0_s0_address;           // mm_interconnect_1:mm_bridge_s0_s0_address -> mm_bridge_s0:s0_address
	wire         mm_interconnect_1_mm_bridge_s0_s0_write;             // mm_interconnect_1:mm_bridge_s0_s0_write -> mm_bridge_s0:s0_write
	wire         mm_interconnect_1_mm_bridge_s0_s0_read;              // mm_interconnect_1:mm_bridge_s0_s0_read -> mm_bridge_s0:s0_read
	wire  [31:0] mm_interconnect_1_mm_bridge_s0_s0_readdata;          // mm_bridge_s0:s0_readdata -> mm_interconnect_1:mm_bridge_s0_s0_readdata
	wire         mm_interconnect_1_mm_bridge_s0_s0_debugaccess;       // mm_interconnect_1:mm_bridge_s0_s0_debugaccess -> mm_bridge_s0:s0_debugaccess
	wire         mm_interconnect_1_mm_bridge_s0_s0_readdatavalid;     // mm_bridge_s0:s0_readdatavalid -> mm_interconnect_1:mm_bridge_s0_s0_readdatavalid
	wire   [3:0] mm_interconnect_1_mm_bridge_s0_s0_byteenable;        // mm_interconnect_1:mm_bridge_s0_s0_byteenable -> mm_bridge_s0:s0_byteenable
	wire         mm_interconnect_1_mm_bridge_s1_s0_waitrequest;       // mm_bridge_s1:s0_waitrequest -> mm_interconnect_1:mm_bridge_s1_s0_waitrequest
	wire   [3:0] mm_interconnect_1_mm_bridge_s1_s0_burstcount;        // mm_interconnect_1:mm_bridge_s1_s0_burstcount -> mm_bridge_s1:s0_burstcount
	wire  [31:0] mm_interconnect_1_mm_bridge_s1_s0_writedata;         // mm_interconnect_1:mm_bridge_s1_s0_writedata -> mm_bridge_s1:s0_writedata
	wire  [17:0] mm_interconnect_1_mm_bridge_s1_s0_address;           // mm_interconnect_1:mm_bridge_s1_s0_address -> mm_bridge_s1:s0_address
	wire         mm_interconnect_1_mm_bridge_s1_s0_write;             // mm_interconnect_1:mm_bridge_s1_s0_write -> mm_bridge_s1:s0_write
	wire         mm_interconnect_1_mm_bridge_s1_s0_read;              // mm_interconnect_1:mm_bridge_s1_s0_read -> mm_bridge_s1:s0_read
	wire  [31:0] mm_interconnect_1_mm_bridge_s1_s0_readdata;          // mm_bridge_s1:s0_readdata -> mm_interconnect_1:mm_bridge_s1_s0_readdata
	wire         mm_interconnect_1_mm_bridge_s1_s0_debugaccess;       // mm_interconnect_1:mm_bridge_s1_s0_debugaccess -> mm_bridge_s1:s0_debugaccess
	wire         mm_interconnect_1_mm_bridge_s1_s0_readdatavalid;     // mm_bridge_s1:s0_readdatavalid -> mm_interconnect_1:mm_bridge_s1_s0_readdatavalid
	wire   [3:0] mm_interconnect_1_mm_bridge_s1_s0_byteenable;        // mm_interconnect_1:mm_bridge_s1_s0_byteenable -> mm_bridge_s1:s0_byteenable
	wire         mm_interconnect_1_mm_bridge_s2_s0_waitrequest;       // mm_bridge_s2:s0_waitrequest -> mm_interconnect_1:mm_bridge_s2_s0_waitrequest
	wire   [3:0] mm_interconnect_1_mm_bridge_s2_s0_burstcount;        // mm_interconnect_1:mm_bridge_s2_s0_burstcount -> mm_bridge_s2:s0_burstcount
	wire  [31:0] mm_interconnect_1_mm_bridge_s2_s0_writedata;         // mm_interconnect_1:mm_bridge_s2_s0_writedata -> mm_bridge_s2:s0_writedata
	wire  [17:0] mm_interconnect_1_mm_bridge_s2_s0_address;           // mm_interconnect_1:mm_bridge_s2_s0_address -> mm_bridge_s2:s0_address
	wire         mm_interconnect_1_mm_bridge_s2_s0_write;             // mm_interconnect_1:mm_bridge_s2_s0_write -> mm_bridge_s2:s0_write
	wire         mm_interconnect_1_mm_bridge_s2_s0_read;              // mm_interconnect_1:mm_bridge_s2_s0_read -> mm_bridge_s2:s0_read
	wire  [31:0] mm_interconnect_1_mm_bridge_s2_s0_readdata;          // mm_bridge_s2:s0_readdata -> mm_interconnect_1:mm_bridge_s2_s0_readdata
	wire         mm_interconnect_1_mm_bridge_s2_s0_debugaccess;       // mm_interconnect_1:mm_bridge_s2_s0_debugaccess -> mm_bridge_s2:s0_debugaccess
	wire         mm_interconnect_1_mm_bridge_s2_s0_readdatavalid;     // mm_bridge_s2:s0_readdatavalid -> mm_interconnect_1:mm_bridge_s2_s0_readdatavalid
	wire   [3:0] mm_interconnect_1_mm_bridge_s2_s0_byteenable;        // mm_interconnect_1:mm_bridge_s2_s0_byteenable -> mm_bridge_s2:s0_byteenable
	wire         mm_interconnect_1_mm_bridge_s3_s0_waitrequest;       // mm_bridge_s3:s0_waitrequest -> mm_interconnect_1:mm_bridge_s3_s0_waitrequest
	wire   [3:0] mm_interconnect_1_mm_bridge_s3_s0_burstcount;        // mm_interconnect_1:mm_bridge_s3_s0_burstcount -> mm_bridge_s3:s0_burstcount
	wire  [31:0] mm_interconnect_1_mm_bridge_s3_s0_writedata;         // mm_interconnect_1:mm_bridge_s3_s0_writedata -> mm_bridge_s3:s0_writedata
	wire  [23:0] mm_interconnect_1_mm_bridge_s3_s0_address;           // mm_interconnect_1:mm_bridge_s3_s0_address -> mm_bridge_s3:s0_address
	wire         mm_interconnect_1_mm_bridge_s3_s0_write;             // mm_interconnect_1:mm_bridge_s3_s0_write -> mm_bridge_s3:s0_write
	wire         mm_interconnect_1_mm_bridge_s3_s0_read;              // mm_interconnect_1:mm_bridge_s3_s0_read -> mm_bridge_s3:s0_read
	wire  [31:0] mm_interconnect_1_mm_bridge_s3_s0_readdata;          // mm_bridge_s3:s0_readdata -> mm_interconnect_1:mm_bridge_s3_s0_readdata
	wire         mm_interconnect_1_mm_bridge_s3_s0_debugaccess;       // mm_interconnect_1:mm_bridge_s3_s0_debugaccess -> mm_bridge_s3:s0_debugaccess
	wire         mm_interconnect_1_mm_bridge_s3_s0_readdatavalid;     // mm_bridge_s3:s0_readdatavalid -> mm_interconnect_1:mm_bridge_s3_s0_readdatavalid
	wire   [3:0] mm_interconnect_1_mm_bridge_s3_s0_byteenable;        // mm_interconnect_1:mm_bridge_s3_s0_byteenable -> mm_bridge_s3:s0_byteenable
	wire         mm_interconnect_1_mm_bridge_s4_s0_waitrequest;       // mm_bridge_s4:s0_waitrequest -> mm_interconnect_1:mm_bridge_s4_s0_waitrequest
	wire   [3:0] mm_interconnect_1_mm_bridge_s4_s0_burstcount;        // mm_interconnect_1:mm_bridge_s4_s0_burstcount -> mm_bridge_s4:s0_burstcount
	wire  [31:0] mm_interconnect_1_mm_bridge_s4_s0_writedata;         // mm_interconnect_1:mm_bridge_s4_s0_writedata -> mm_bridge_s4:s0_writedata
	wire  [17:0] mm_interconnect_1_mm_bridge_s4_s0_address;           // mm_interconnect_1:mm_bridge_s4_s0_address -> mm_bridge_s4:s0_address
	wire         mm_interconnect_1_mm_bridge_s4_s0_write;             // mm_interconnect_1:mm_bridge_s4_s0_write -> mm_bridge_s4:s0_write
	wire         mm_interconnect_1_mm_bridge_s4_s0_read;              // mm_interconnect_1:mm_bridge_s4_s0_read -> mm_bridge_s4:s0_read
	wire  [31:0] mm_interconnect_1_mm_bridge_s4_s0_readdata;          // mm_bridge_s4:s0_readdata -> mm_interconnect_1:mm_bridge_s4_s0_readdata
	wire         mm_interconnect_1_mm_bridge_s4_s0_debugaccess;       // mm_interconnect_1:mm_bridge_s4_s0_debugaccess -> mm_bridge_s4:s0_debugaccess
	wire         mm_interconnect_1_mm_bridge_s4_s0_readdatavalid;     // mm_bridge_s4:s0_readdatavalid -> mm_interconnect_1:mm_bridge_s4_s0_readdatavalid
	wire   [3:0] mm_interconnect_1_mm_bridge_s4_s0_byteenable;        // mm_interconnect_1:mm_bridge_s4_s0_byteenable -> mm_bridge_s4:s0_byteenable
	wire         mm_interconnect_1_mm_bridge_s5_s0_waitrequest;       // mm_bridge_s5:s0_waitrequest -> mm_interconnect_1:mm_bridge_s5_s0_waitrequest
	wire   [3:0] mm_interconnect_1_mm_bridge_s5_s0_burstcount;        // mm_interconnect_1:mm_bridge_s5_s0_burstcount -> mm_bridge_s5:s0_burstcount
	wire  [31:0] mm_interconnect_1_mm_bridge_s5_s0_writedata;         // mm_interconnect_1:mm_bridge_s5_s0_writedata -> mm_bridge_s5:s0_writedata
	wire  [17:0] mm_interconnect_1_mm_bridge_s5_s0_address;           // mm_interconnect_1:mm_bridge_s5_s0_address -> mm_bridge_s5:s0_address
	wire         mm_interconnect_1_mm_bridge_s5_s0_write;             // mm_interconnect_1:mm_bridge_s5_s0_write -> mm_bridge_s5:s0_write
	wire         mm_interconnect_1_mm_bridge_s5_s0_read;              // mm_interconnect_1:mm_bridge_s5_s0_read -> mm_bridge_s5:s0_read
	wire  [31:0] mm_interconnect_1_mm_bridge_s5_s0_readdata;          // mm_bridge_s5:s0_readdata -> mm_interconnect_1:mm_bridge_s5_s0_readdata
	wire         mm_interconnect_1_mm_bridge_s5_s0_debugaccess;       // mm_interconnect_1:mm_bridge_s5_s0_debugaccess -> mm_bridge_s5:s0_debugaccess
	wire         mm_interconnect_1_mm_bridge_s5_s0_readdatavalid;     // mm_bridge_s5:s0_readdatavalid -> mm_interconnect_1:mm_bridge_s5_s0_readdatavalid
	wire   [3:0] mm_interconnect_1_mm_bridge_s5_s0_byteenable;        // mm_interconnect_1:mm_bridge_s5_s0_byteenable -> mm_bridge_s5:s0_byteenable
	wire         mm_interconnect_1_mm_bridge_s6_s0_waitrequest;       // mm_bridge_s6:s0_waitrequest -> mm_interconnect_1:mm_bridge_s6_s0_waitrequest
	wire   [3:0] mm_interconnect_1_mm_bridge_s6_s0_burstcount;        // mm_interconnect_1:mm_bridge_s6_s0_burstcount -> mm_bridge_s6:s0_burstcount
	wire  [31:0] mm_interconnect_1_mm_bridge_s6_s0_writedata;         // mm_interconnect_1:mm_bridge_s6_s0_writedata -> mm_bridge_s6:s0_writedata
	wire  [17:0] mm_interconnect_1_mm_bridge_s6_s0_address;           // mm_interconnect_1:mm_bridge_s6_s0_address -> mm_bridge_s6:s0_address
	wire         mm_interconnect_1_mm_bridge_s6_s0_write;             // mm_interconnect_1:mm_bridge_s6_s0_write -> mm_bridge_s6:s0_write
	wire         mm_interconnect_1_mm_bridge_s6_s0_read;              // mm_interconnect_1:mm_bridge_s6_s0_read -> mm_bridge_s6:s0_read
	wire  [31:0] mm_interconnect_1_mm_bridge_s6_s0_readdata;          // mm_bridge_s6:s0_readdata -> mm_interconnect_1:mm_bridge_s6_s0_readdata
	wire         mm_interconnect_1_mm_bridge_s6_s0_debugaccess;       // mm_interconnect_1:mm_bridge_s6_s0_debugaccess -> mm_bridge_s6:s0_debugaccess
	wire         mm_interconnect_1_mm_bridge_s6_s0_readdatavalid;     // mm_bridge_s6:s0_readdatavalid -> mm_interconnect_1:mm_bridge_s6_s0_readdatavalid
	wire   [3:0] mm_interconnect_1_mm_bridge_s6_s0_byteenable;        // mm_interconnect_1:mm_bridge_s6_s0_byteenable -> mm_bridge_s6:s0_byteenable
	wire         rst_controller_reset_out_reset;                      // rst_controller:reset_out -> [mm_bridge_master:reset, mm_bridge_s0:reset, mm_bridge_s1:reset, mm_bridge_s2:reset, mm_bridge_s3:reset, mm_bridge_s4:reset, mm_bridge_s5:reset, mm_bridge_s6:reset, mm_interconnect_0:jtag_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mm_bridge_master_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_bridge_master_reset_reset_bridge_in_reset_reset]

	jtag_system_jtag_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_master (
		.clk_clk              (clk_clk),                          //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                   //    clk_reset.reset
		.master_address       (jtag_master_master_address),       //       master.address
		.master_readdata      (jtag_master_master_readdata),      //             .readdata
		.master_read          (jtag_master_master_read),          //             .read
		.master_write         (jtag_master_master_write),         //             .write
		.master_writedata     (jtag_master_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_master_master_byteenable),    //             .byteenable
		.master_reset_reset   (resetrequest_reset)                // master_reset.reset
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (4),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_master (
		.clk              (clk_clk),                                             //   clk.clk
		.reset            (rst_controller_reset_out_reset),                      // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_master_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_master_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_master_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_master_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_master_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_master_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_master_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_master_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_master_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_master_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_master_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_master_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_master_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_master_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_master_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_master_m0_address),                         //      .address
		.m0_write         (mm_bridge_master_m0_write),                           //      .write
		.m0_read          (mm_bridge_master_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_master_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_master_m0_debugaccess)                      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (24),
		.BURSTCOUNT_WIDTH  (4),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_s0 (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (rst_controller_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_s0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_s0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_s0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_s0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_s0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_s0_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_s0_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_s0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_s0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_s0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_s0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_s0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_s0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_s0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_s0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_s0_m0_address),                         //      .address
		.m0_write         (mm_bridge_s0_m0_write),                           //      .write
		.m0_read          (mm_bridge_s0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_s0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_s0_m0_debugaccess)                      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (18),
		.BURSTCOUNT_WIDTH  (4),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_s1 (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (rst_controller_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_s1_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_s1_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_s1_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_s1_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_s1_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_s1_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_s1_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_s1_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_s1_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_s1_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_s1_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_s1_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_s1_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_s1_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_s1_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_s1_m0_address),                         //      .address
		.m0_write         (mm_bridge_s1_m0_write),                           //      .write
		.m0_read          (mm_bridge_s1_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_s1_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_s1_m0_debugaccess)                      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (18),
		.BURSTCOUNT_WIDTH  (4),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_s2 (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (rst_controller_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_s2_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_s2_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_s2_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_s2_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_s2_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_s2_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_s2_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_s2_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_s2_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_s2_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_s2_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_s2_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_s2_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_s2_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_s2_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_s2_m0_address),                         //      .address
		.m0_write         (mm_bridge_s2_m0_write),                           //      .write
		.m0_read          (mm_bridge_s2_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_s2_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_s2_m0_debugaccess)                      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (24),
		.BURSTCOUNT_WIDTH  (4),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_s3 (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (rst_controller_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_s3_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_s3_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_s3_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_s3_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_s3_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_s3_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_s3_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_s3_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_s3_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_s3_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_s3_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_s3_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_s3_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_s3_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_s3_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_s3_m0_address),                         //      .address
		.m0_write         (mm_bridge_s3_m0_write),                           //      .write
		.m0_read          (mm_bridge_s3_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_s3_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_s3_m0_debugaccess)                      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (18),
		.BURSTCOUNT_WIDTH  (4),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_s4 (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (rst_controller_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_s4_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_s4_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_s4_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_s4_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_s4_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_s4_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_s4_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_s4_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_s4_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_s4_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_s4_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_s4_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_s4_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_s4_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_s4_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_s4_m0_address),                         //      .address
		.m0_write         (mm_bridge_s4_m0_write),                           //      .write
		.m0_read          (mm_bridge_s4_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_s4_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_s4_m0_debugaccess)                      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (18),
		.BURSTCOUNT_WIDTH  (4),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_s5 (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (rst_controller_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_s5_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_s5_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_s5_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_s5_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_s5_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_s5_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_s5_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_s5_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_s5_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_s5_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_s5_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_s5_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_s5_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_s5_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_s5_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_s5_m0_address),                         //      .address
		.m0_write         (mm_bridge_s5_m0_write),                           //      .write
		.m0_read          (mm_bridge_s5_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_s5_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_s5_m0_debugaccess)                      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (18),
		.BURSTCOUNT_WIDTH  (4),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_s6 (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (rst_controller_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_s6_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_s6_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_s6_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_s6_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_s6_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_s6_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_s6_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_s6_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_s6_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_s6_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_s6_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_s6_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_s6_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_s6_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_s6_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_s6_m0_address),                         //      .address
		.m0_write         (mm_bridge_s6_m0_write),                           //      .write
		.m0_read          (mm_bridge_s6_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_s6_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_s6_m0_debugaccess)                      //      .debugaccess
	);

	jtag_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                        (clk_clk),                                             //                                      clk_clk.clk
		.jtag_master_clk_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                      //  jtag_master_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_master_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                      // mm_bridge_master_reset_reset_bridge_in_reset.reset
		.jtag_master_master_address                         (jtag_master_master_address),                          //                           jtag_master_master.address
		.jtag_master_master_waitrequest                     (jtag_master_master_waitrequest),                      //                                             .waitrequest
		.jtag_master_master_byteenable                      (jtag_master_master_byteenable),                       //                                             .byteenable
		.jtag_master_master_read                            (jtag_master_master_read),                             //                                             .read
		.jtag_master_master_readdata                        (jtag_master_master_readdata),                         //                                             .readdata
		.jtag_master_master_readdatavalid                   (jtag_master_master_readdatavalid),                    //                                             .readdatavalid
		.jtag_master_master_write                           (jtag_master_master_write),                            //                                             .write
		.jtag_master_master_writedata                       (jtag_master_master_writedata),                        //                                             .writedata
		.mm_bridge_master_s0_address                        (mm_interconnect_0_mm_bridge_master_s0_address),       //                          mm_bridge_master_s0.address
		.mm_bridge_master_s0_write                          (mm_interconnect_0_mm_bridge_master_s0_write),         //                                             .write
		.mm_bridge_master_s0_read                           (mm_interconnect_0_mm_bridge_master_s0_read),          //                                             .read
		.mm_bridge_master_s0_readdata                       (mm_interconnect_0_mm_bridge_master_s0_readdata),      //                                             .readdata
		.mm_bridge_master_s0_writedata                      (mm_interconnect_0_mm_bridge_master_s0_writedata),     //                                             .writedata
		.mm_bridge_master_s0_burstcount                     (mm_interconnect_0_mm_bridge_master_s0_burstcount),    //                                             .burstcount
		.mm_bridge_master_s0_byteenable                     (mm_interconnect_0_mm_bridge_master_s0_byteenable),    //                                             .byteenable
		.mm_bridge_master_s0_readdatavalid                  (mm_interconnect_0_mm_bridge_master_s0_readdatavalid), //                                             .readdatavalid
		.mm_bridge_master_s0_waitrequest                    (mm_interconnect_0_mm_bridge_master_s0_waitrequest),   //                                             .waitrequest
		.mm_bridge_master_s0_debugaccess                    (mm_interconnect_0_mm_bridge_master_s0_debugaccess)    //                                             .debugaccess
	);

	jtag_system_mm_interconnect_1 mm_interconnect_1 (
		.clk_clk_clk                                        (clk_clk),                                         //                                      clk_clk.clk
		.mm_bridge_master_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                  // mm_bridge_master_reset_reset_bridge_in_reset.reset
		.mm_bridge_master_m0_address                        (mm_bridge_master_m0_address),                     //                          mm_bridge_master_m0.address
		.mm_bridge_master_m0_waitrequest                    (mm_bridge_master_m0_waitrequest),                 //                                             .waitrequest
		.mm_bridge_master_m0_burstcount                     (mm_bridge_master_m0_burstcount),                  //                                             .burstcount
		.mm_bridge_master_m0_byteenable                     (mm_bridge_master_m0_byteenable),                  //                                             .byteenable
		.mm_bridge_master_m0_read                           (mm_bridge_master_m0_read),                        //                                             .read
		.mm_bridge_master_m0_readdata                       (mm_bridge_master_m0_readdata),                    //                                             .readdata
		.mm_bridge_master_m0_readdatavalid                  (mm_bridge_master_m0_readdatavalid),               //                                             .readdatavalid
		.mm_bridge_master_m0_write                          (mm_bridge_master_m0_write),                       //                                             .write
		.mm_bridge_master_m0_writedata                      (mm_bridge_master_m0_writedata),                   //                                             .writedata
		.mm_bridge_master_m0_debugaccess                    (mm_bridge_master_m0_debugaccess),                 //                                             .debugaccess
		.mm_bridge_s0_s0_address                            (mm_interconnect_1_mm_bridge_s0_s0_address),       //                              mm_bridge_s0_s0.address
		.mm_bridge_s0_s0_write                              (mm_interconnect_1_mm_bridge_s0_s0_write),         //                                             .write
		.mm_bridge_s0_s0_read                               (mm_interconnect_1_mm_bridge_s0_s0_read),          //                                             .read
		.mm_bridge_s0_s0_readdata                           (mm_interconnect_1_mm_bridge_s0_s0_readdata),      //                                             .readdata
		.mm_bridge_s0_s0_writedata                          (mm_interconnect_1_mm_bridge_s0_s0_writedata),     //                                             .writedata
		.mm_bridge_s0_s0_burstcount                         (mm_interconnect_1_mm_bridge_s0_s0_burstcount),    //                                             .burstcount
		.mm_bridge_s0_s0_byteenable                         (mm_interconnect_1_mm_bridge_s0_s0_byteenable),    //                                             .byteenable
		.mm_bridge_s0_s0_readdatavalid                      (mm_interconnect_1_mm_bridge_s0_s0_readdatavalid), //                                             .readdatavalid
		.mm_bridge_s0_s0_waitrequest                        (mm_interconnect_1_mm_bridge_s0_s0_waitrequest),   //                                             .waitrequest
		.mm_bridge_s0_s0_debugaccess                        (mm_interconnect_1_mm_bridge_s0_s0_debugaccess),   //                                             .debugaccess
		.mm_bridge_s1_s0_address                            (mm_interconnect_1_mm_bridge_s1_s0_address),       //                              mm_bridge_s1_s0.address
		.mm_bridge_s1_s0_write                              (mm_interconnect_1_mm_bridge_s1_s0_write),         //                                             .write
		.mm_bridge_s1_s0_read                               (mm_interconnect_1_mm_bridge_s1_s0_read),          //                                             .read
		.mm_bridge_s1_s0_readdata                           (mm_interconnect_1_mm_bridge_s1_s0_readdata),      //                                             .readdata
		.mm_bridge_s1_s0_writedata                          (mm_interconnect_1_mm_bridge_s1_s0_writedata),     //                                             .writedata
		.mm_bridge_s1_s0_burstcount                         (mm_interconnect_1_mm_bridge_s1_s0_burstcount),    //                                             .burstcount
		.mm_bridge_s1_s0_byteenable                         (mm_interconnect_1_mm_bridge_s1_s0_byteenable),    //                                             .byteenable
		.mm_bridge_s1_s0_readdatavalid                      (mm_interconnect_1_mm_bridge_s1_s0_readdatavalid), //                                             .readdatavalid
		.mm_bridge_s1_s0_waitrequest                        (mm_interconnect_1_mm_bridge_s1_s0_waitrequest),   //                                             .waitrequest
		.mm_bridge_s1_s0_debugaccess                        (mm_interconnect_1_mm_bridge_s1_s0_debugaccess),   //                                             .debugaccess
		.mm_bridge_s2_s0_address                            (mm_interconnect_1_mm_bridge_s2_s0_address),       //                              mm_bridge_s2_s0.address
		.mm_bridge_s2_s0_write                              (mm_interconnect_1_mm_bridge_s2_s0_write),         //                                             .write
		.mm_bridge_s2_s0_read                               (mm_interconnect_1_mm_bridge_s2_s0_read),          //                                             .read
		.mm_bridge_s2_s0_readdata                           (mm_interconnect_1_mm_bridge_s2_s0_readdata),      //                                             .readdata
		.mm_bridge_s2_s0_writedata                          (mm_interconnect_1_mm_bridge_s2_s0_writedata),     //                                             .writedata
		.mm_bridge_s2_s0_burstcount                         (mm_interconnect_1_mm_bridge_s2_s0_burstcount),    //                                             .burstcount
		.mm_bridge_s2_s0_byteenable                         (mm_interconnect_1_mm_bridge_s2_s0_byteenable),    //                                             .byteenable
		.mm_bridge_s2_s0_readdatavalid                      (mm_interconnect_1_mm_bridge_s2_s0_readdatavalid), //                                             .readdatavalid
		.mm_bridge_s2_s0_waitrequest                        (mm_interconnect_1_mm_bridge_s2_s0_waitrequest),   //                                             .waitrequest
		.mm_bridge_s2_s0_debugaccess                        (mm_interconnect_1_mm_bridge_s2_s0_debugaccess),   //                                             .debugaccess
		.mm_bridge_s3_s0_address                            (mm_interconnect_1_mm_bridge_s3_s0_address),       //                              mm_bridge_s3_s0.address
		.mm_bridge_s3_s0_write                              (mm_interconnect_1_mm_bridge_s3_s0_write),         //                                             .write
		.mm_bridge_s3_s0_read                               (mm_interconnect_1_mm_bridge_s3_s0_read),          //                                             .read
		.mm_bridge_s3_s0_readdata                           (mm_interconnect_1_mm_bridge_s3_s0_readdata),      //                                             .readdata
		.mm_bridge_s3_s0_writedata                          (mm_interconnect_1_mm_bridge_s3_s0_writedata),     //                                             .writedata
		.mm_bridge_s3_s0_burstcount                         (mm_interconnect_1_mm_bridge_s3_s0_burstcount),    //                                             .burstcount
		.mm_bridge_s3_s0_byteenable                         (mm_interconnect_1_mm_bridge_s3_s0_byteenable),    //                                             .byteenable
		.mm_bridge_s3_s0_readdatavalid                      (mm_interconnect_1_mm_bridge_s3_s0_readdatavalid), //                                             .readdatavalid
		.mm_bridge_s3_s0_waitrequest                        (mm_interconnect_1_mm_bridge_s3_s0_waitrequest),   //                                             .waitrequest
		.mm_bridge_s3_s0_debugaccess                        (mm_interconnect_1_mm_bridge_s3_s0_debugaccess),   //                                             .debugaccess
		.mm_bridge_s4_s0_address                            (mm_interconnect_1_mm_bridge_s4_s0_address),       //                              mm_bridge_s4_s0.address
		.mm_bridge_s4_s0_write                              (mm_interconnect_1_mm_bridge_s4_s0_write),         //                                             .write
		.mm_bridge_s4_s0_read                               (mm_interconnect_1_mm_bridge_s4_s0_read),          //                                             .read
		.mm_bridge_s4_s0_readdata                           (mm_interconnect_1_mm_bridge_s4_s0_readdata),      //                                             .readdata
		.mm_bridge_s4_s0_writedata                          (mm_interconnect_1_mm_bridge_s4_s0_writedata),     //                                             .writedata
		.mm_bridge_s4_s0_burstcount                         (mm_interconnect_1_mm_bridge_s4_s0_burstcount),    //                                             .burstcount
		.mm_bridge_s4_s0_byteenable                         (mm_interconnect_1_mm_bridge_s4_s0_byteenable),    //                                             .byteenable
		.mm_bridge_s4_s0_readdatavalid                      (mm_interconnect_1_mm_bridge_s4_s0_readdatavalid), //                                             .readdatavalid
		.mm_bridge_s4_s0_waitrequest                        (mm_interconnect_1_mm_bridge_s4_s0_waitrequest),   //                                             .waitrequest
		.mm_bridge_s4_s0_debugaccess                        (mm_interconnect_1_mm_bridge_s4_s0_debugaccess),   //                                             .debugaccess
		.mm_bridge_s5_s0_address                            (mm_interconnect_1_mm_bridge_s5_s0_address),       //                              mm_bridge_s5_s0.address
		.mm_bridge_s5_s0_write                              (mm_interconnect_1_mm_bridge_s5_s0_write),         //                                             .write
		.mm_bridge_s5_s0_read                               (mm_interconnect_1_mm_bridge_s5_s0_read),          //                                             .read
		.mm_bridge_s5_s0_readdata                           (mm_interconnect_1_mm_bridge_s5_s0_readdata),      //                                             .readdata
		.mm_bridge_s5_s0_writedata                          (mm_interconnect_1_mm_bridge_s5_s0_writedata),     //                                             .writedata
		.mm_bridge_s5_s0_burstcount                         (mm_interconnect_1_mm_bridge_s5_s0_burstcount),    //                                             .burstcount
		.mm_bridge_s5_s0_byteenable                         (mm_interconnect_1_mm_bridge_s5_s0_byteenable),    //                                             .byteenable
		.mm_bridge_s5_s0_readdatavalid                      (mm_interconnect_1_mm_bridge_s5_s0_readdatavalid), //                                             .readdatavalid
		.mm_bridge_s5_s0_waitrequest                        (mm_interconnect_1_mm_bridge_s5_s0_waitrequest),   //                                             .waitrequest
		.mm_bridge_s5_s0_debugaccess                        (mm_interconnect_1_mm_bridge_s5_s0_debugaccess),   //                                             .debugaccess
		.mm_bridge_s6_s0_address                            (mm_interconnect_1_mm_bridge_s6_s0_address),       //                              mm_bridge_s6_s0.address
		.mm_bridge_s6_s0_write                              (mm_interconnect_1_mm_bridge_s6_s0_write),         //                                             .write
		.mm_bridge_s6_s0_read                               (mm_interconnect_1_mm_bridge_s6_s0_read),          //                                             .read
		.mm_bridge_s6_s0_readdata                           (mm_interconnect_1_mm_bridge_s6_s0_readdata),      //                                             .readdata
		.mm_bridge_s6_s0_writedata                          (mm_interconnect_1_mm_bridge_s6_s0_writedata),     //                                             .writedata
		.mm_bridge_s6_s0_burstcount                         (mm_interconnect_1_mm_bridge_s6_s0_burstcount),    //                                             .burstcount
		.mm_bridge_s6_s0_byteenable                         (mm_interconnect_1_mm_bridge_s6_s0_byteenable),    //                                             .byteenable
		.mm_bridge_s6_s0_readdatavalid                      (mm_interconnect_1_mm_bridge_s6_s0_readdatavalid), //                                             .readdatavalid
		.mm_bridge_s6_s0_waitrequest                        (mm_interconnect_1_mm_bridge_s6_s0_waitrequest),   //                                             .waitrequest
		.mm_bridge_s6_s0_debugaccess                        (mm_interconnect_1_mm_bridge_s6_s0_debugaccess)    //                                             .debugaccess
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule

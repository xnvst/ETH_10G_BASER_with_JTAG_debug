// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
o7oOTsPyLa8O8A/AFTzZweteYGjNa/gWjqlNOfVpXbN4IkSO3iyv2p/FtgrfvYlE/sLWi4QaFbeC
aUhT2GRmI4buFpbWTgPdFaretS1+++CeR7XP3MRAhWW8Cx72mBG6dr1cIPnfvoUGHtLhoaeC+OIA
TRECkJPE2jDghrrnrCx8108cHURganiclPuRAZmhGtP1KMw9nn4rqq22q9FAlMyZ+ufYBd0D3asv
EIyZoALAoaIS7YaONkEK+/PE0jpRQ7CHjQXIsMaGj4Lq/AXU+lYo22CE/00EEcHANsyQTpswuuG/
57LCSUJJHboeBsrsgy2TrICRYl+XG2tf0Nfo+w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
QrSEEK1XNCkbsow7Arp4XM1fWcXWclGTS+0QCi1KMVOj/n4BLuR+AiRriAR2yxeiqDPvqt9GN5I9
XTM5JE1VNvFlIhvTqqH54o1HAPTpJj38mutPhYmOC9ex14wHgFA5TlHYOHY+G5W1vauppC+dZUvo
4+UtA27OIsz19zPCuZJpvio5mbBRiwJd+TOtz7SwCgYka3x7dATlc7wGbDai6o3H6GHGwAAoB1sn
NqtKsMLfwsLzSIs1q0nt789PudqgpY1qtwwikGt5fymef+RO9DbWricy7FPaMkp3vlFt+AFm/OfR
l50tePmMdGKe7T1khV1MmlItCTtj1uZIEsbknkJYOOaKWNE2zWHvQy0YpjY816xg11IMW4shTo1l
V/fJJOzudZk30nou1Mstwqu4a5P1mobmIjmzLicuzrYNASSike+X1dt1mXx4udi9Ef3i9eujBBb2
fV2CJqpQ58H9P3mJb9KQHgD8AfWQfu/kltJeaWJSxD1UNSdCWpqtOu8sMzizkuy9Zve0+FJJQN9u
tf/gur2GDPU28kqeW93Wt9zrEpQyeFQYpJ+pvMhruNtGP/tijaEC6LM28o8oVU5uqMHzxYUv+f1k
z8mS3R84kw8WZkRS6MWDuDu5LamkPvNqogNsilw/N0gDbnZ3/TPcLQEu+5sSec6MmTTmFeXO74IO
D8sC/fq0it9K/PJnes+OYDCjP4a12EYj7gUplkL3dz2YJqNuuMvr+iKD0kbcNF2ZEeRauTYUfDNc
uSjG5xpsxHmDfcyjXv0r9TJwzCSVP8alSqdynmyKY7r5DpuHGfkfbI6DfdRBSa9/yll4tIxS3Tme
tp5boqdW0u7Y3OX2+pKBfr1Lm9q3U4z9/17FkxdZZqezKjofRyo65IKfLWii4thBmbIRbc0tJ6gV
UqnI0vu6Q39YDFApF4Fb40wfpX2FExWPYnWY+V5SzSA+NR44Xt86/o8RGX8J/ztWYiTS0CwHIjV4
oQmq0YYSFSLwrrE1agUwCYkbHan9/f/tjFJN2x5gj+80azd9jA/5WnVhSmmHvluWydQAQyUlL460
QMtR5xOI+xzObb88NJlzdkZlRT9zupZEGdwuTTFJoX42nvZK4rHLMXaomczuImJ2shEq7gOW0huU
ZQYY2dDkFxXOn4j989dBhHm19/UEllAZ+Y945gImcPc3ue9RE8IjD080jJh1yO6SYbB6cb7KwhDk
bIlaloeDmCN5lGsP9BEIfN+RrNBB+rOWNtRco5CgeTRn7KtLxIFeHe8vNZ+vHQWTZvdNwpntHUWi
mymY4qdMUAGY0zoktEkE2JttK/VWU1LdfS6CzweZHi94Rpiom5oyYd1mZUk3tmhZ0HM4JD/Bxnfv
lf/ecuOSbRazG+8ZkkR1sqM5PABd86HvH5NPQ9PP4Jtc8K4yR/w6GhKSxwQGfhz71Zk2x8nTe8TI
aOAwxJmbSegkx5kppFX93x3/1NxV9zpoJQCzTvhEOPaCPYlRrKeurWRHupMWNFXXmurKlklHA3hW
Nh8npU0QaKnLEFIYfBQ8EXQYM+nC2x0gshunPEl9870mF9qt2yF5YrjwzRkm1jI0BQGBHUFGk8E7
XaB+dqTKXXGrFHX44iDDENy+dBz4SqanKT5EbQN+MvSq/rCqjdflcG69BnNPnnJtAWe2vW4c4Vhx
FIzZ1QD/3aZm3cEqMxBmoiJS9k5aTskh9SMxeafWWj0roIUyC44RVV4kNpEFDVVjd/mMn0/hZ9sY
yuOgZYKf1zW7Fnnf+KGqJ/DnWxAqIq9ox2LuvEyKJ0nNxMO2zN2B7i9tkH/9iYICWR2JuK3LR6Jg
NiRhOHGLwXzZcMKC54EoujmiChIBPGfVdlq1MbqI+vAJyKXBoYXLmTVI4JACF4n0sPD02zKpkeqW
gP8pIt1niNcYu5oom3x/pubxY2L0zKot2H61uh4hfpav7s1f5p0xD9Eju30iZPaDpnCmls5pN4rt
uKR6+WA79sxbY01lRxq904PdTBKqKCw0N093vL07tWAQTA7PMUOJfQ3/1Pe1eqzhQg4ukTKNmg9A
Dyc24pDEWPx7JRihCo1fSR3xE7YY1Y0hdte0OlPqb87JpTc/5d97jq4XLgw2D+HGZiBK89gL3m4J
wemdFuDDi4UnFhLI97j6szE895dyzIFLkQ5VsEOqznLcsLtQEHBF2YCT/HR6hsYZ9cSa0ru6xaoi
5ohjy6QMJFQGsuxCyN0vIQMx4ITfEv1MIlule57par7+XM7vwg37x8wWom3ZfRRHMDd1dyh2tKcF
s4Vsp7Ymtn9ei1uVZKKMkI4OrbITPcSjBaSqT+P/hltSH9JsJqf7VJU0LJ/F34lutRAoEOoULIrx
ZsauvWPhj/Qyc2AzTlwDBWF7k8MMS6QnzW3Ky0ibiPvxAH/KUZevCAW/hKrNqMbRLiiqHyot6Zlt
YuWwFfLiFTDmIe9KkaTSuzKDxsnPd2LB69R8q2k7vhpyBZsCCb6P2YJM+B2/r12CzsUs/Hu4/k9f
NKDayPE6osIa+/9Nbv1C5F9G1sLjplB+tD+bGKzWKPjFGeCP6hRsadIgtHuSPKGbcJkVlfRTrWI8
jr7XQwBrEGGQd/5SVYFYu1cU/XSKF8ac1BkC94HzgwkTX1v9VAv4Sbs8HXcdgEOuPe3v0avWAhfQ
8Je/RYwLT2y85BQOIihLG9G1zw0r97MljRHiGD3Ro2mbYcpaAFc/Qub8KW7TTLl5rugDiKOZOXS8
GIR6KCRNlncfs9IZBOh/UqAiLR1twgn4BtcNmDpDlg7XE4CgQ3BTO+vVj/JPaIud7XQtmM5WneX1
3BK3KFFK35FMX6qnr/x8Rgf13/p7O7nY6Ew399yFVN4w5NcAn4Y+PD8FTGygdhsKBdvAdnHENLs7
cmjfn9CcXzn8Z0VelSpNtAA1dHaDWt2x/b2hXyLTyRdnwy+T6p5GDyta4O9NDrfdV1Zh8gW0MLXr
2NZaPYlS4bM+qikye1d1dxVSM+exnj7I7SJ21BBiz/HMi87SMEsqD8yxB1eeNi4r7eemRBM41wf1
gSWMqYyHXS/CrbhJmWP6O8QKsmsrCS+BcvXFtZ79oNf/ey7+FeM+n8JA7mmQ0ONPMTr7QS+sRFQp
5wX10M2E9lK4r+ifiTo4UFKmnSRlzMITfhfDN/U6K6iW5WMG3BssK4JEMg/PQOBRb9GqzUJA79Zx
pLlgYd72KrxVFaoBqRXX7UqKk3gYNKyxfd0INRLi0Lyt+BE3WFA2dMXnf+agstVJeseoIr9oLjvF
jWNK7ZuL7rJmyj+2d2vIcRcBgQKk8bqDNtHj+m5pNg7QPyZufTy82/uuq9Lg75uLy9s7FAeXU5PH
9EkvjMo269Y9zNkKUCr3eSnQcz0qUiR3ovZiePYS5v8I8XUwUYzPiQk9eQbcXhjjmD3PwzRQqJOL
vALwh11Pax8MhojcEBFitJoIOmc7OKTUwRg3sDOEUC29xN8TvaIV0g0AcVgxVU/y3Icng5aRYYjI
PuOJ9VhOuedKkK0ch1rLquwpq9OwNJR9fGdSlZFc8iWRbZPjb7b/raMKZs3PDlf5NyzpPM6upGVT
6phkmktSJB8D63MCv1xwy76zjekX78mu9LlMDD+sG9Z3ghU1SO5iETe3vtbWj8of6D6CfqgXGl07
WNNAqfHvVbVvSbcbG88MgufrNyf4acY8m+DcefZk4YCrD7e3kg9S8b0sqUNkECM56nO+N0+b6xpj
wWBnDYR7OG8gNsJjE+14/BEkD9ynIbPfZsyQPGsja6LRFls2b7NVg7JW1hOQkYuR+TxKiGt+utgm
ILr95cCumWoaVs+0xy54NBduceBUcZQP1BbeebpenCNheG/t4V6orfmlCgCe04ZStmF9TndbhL4f
AVbLqW1jS9SallQtATgFEosDyYeY2x0XxziUBXn4DhDnW/8d2KxQoez6jn2D7+5MsxvzbgC6FzCB
ZYUCzLHxOb65OdpYgRr+G7qFRPnqG8xAg2T7WsiB9LA059O3KCrWQTJ1ZHb/9KQEhmRl/R1Pdr5u
c+A/PuCzDpTKC44USwHiMTFotjs5k/yDGnsxrgrAoVBYGx10i9faWtnZpx56sdOIEI8ZnjFI7fBK
TOsdWC4qvuPAbdOlZwQV37kjIJcStPdyIZA2BdL9IFWrJYLcynJqn1EE9FWHxevQC3hblArmgHfc
SHNHCNUO+jjiebcNOjBB72rXVfmQjlDgFPFp/4lQ4y2eq9oQPMPjg1fZiLIyOy9FgyDiJ8XrxOn8
kfnen5dWCk+XUfAtJAw17PUu1DYhLzgeAZ0XOCuUfuEq87C0uJqf3hMVu06psVm4Ek9/pAUoYQF7
aP2qbnJPdprq1UiOmIh59SGfTIk8PDHPO9Devr66/76KT83NOoYx/ElvFAnJNBfbnQaaxonh4DG4
oI3KHDi1D3pbmUAErs5ZpSSDF0CTkDXtdG524B7ctXTqSNocZ4kQYZInhzQdbll8qMwc4QQMyw2O
VrXXxz4lXIObHNxaVbXJzTxO6ZcvgQmAFmIkxrpn8XRDRNW4glMQfMukszc0PonKUibtIgm8Wadv
z6kJmz1DIR3nHvSX/CZDWakuiRI8xThAsZM16MlAVIu+Ein9NzMC1pt05s5o0uWpT3hXlALfOKfc
WLWBtZvc9A6nZ0MleGOuFecm94osrR38sN+SOiwJvs1fl2xSscNbiP/kVNABVBwez8eEMTOy6Tfd
WBSihDaJQY1oUMqH2nkOcIwCEUC0IXGNEmiu9hz+DN93HpH76UPRUEGaabGVdiwNCBQlceG1f4s1
vFqzmHa5idsdAP1lpNwAyBKtfDKaVjNPdQTu8nR7fNrxqbB9P3dayHPka7TnF9LTIxKfYWtX3oPA
0t/Uah3UED5fEePSsY2kbPXzdRNCGRfhLOQOXCBoF/gm8F63pBz7EzQpRTxMEowYgfCsYsCkEv/n
n0q9TFn3RIqvfPiy6e168RYCwh47diLq64YxqUC9lnhmMAuqBo6Mf1WSy8dkEUfR/qmOclouO92K
dzCP1p6F1JZi4Bsxr0bBjel7Y9L8X3PW4J41bLheKBWCbWZxcG+zxVMhrjn+STfeJm/PTw7GYv4v
br5yi20VjlDJzJtZF8oytbc0CmBwYODMxlWqhRCMmyFSQudY3oaNKkXcbt/4v5kJ2oye/Gkf6vck
GpcfgIKjNITe+RxuoptgxwgobFHi1EAr6vZ4hQfV/YRyMtRwx8JGzpjYgVo1+xfVGLWk/WC0+2AI
pPKEMDiMqATrF599sPQitVfGtYtyeNQPNjSLSRtLcfXRIH/31ft7L6VTBCvoG7+coh0z1ZlDWym1
itSH9k5BzJwmeGltbqV4LtVaG5vHXoH0ct6UH3bxhQXFSci1phieYsP/K4UN5TZCWlR0p/P/aGUX
9i6/ThzElzNfR39vtymtDi+lwHuZccguncQZfGsIolu5usIR1cgwlQruPWke8Zx4D3BSOSQkjEMm
xCnRXk15EyY8pvRQvRLvppIJ2dl0KkltJ4aZXk3zEGkMIjw2SZnUeggIPrqKgBfIVe363nH5CyQD
W1NdduQ3b/nfCZH0uEenpqVQn6aJ0lYSfAOangeIOnHS1+Fr2CSV0P/SQhFaA6fjvIkXJkwpMUpi
jNdEvG7scYkUoDLUT8sCihN4q+9IH2iB6ieyyMaj8aTOHV1EgzWrzq6VJ6M59gMD/alP/dU0OHtS
SbrWqlmmYx6ct4bkPz89O9p6jBOhvMel9PCNksVG8mZT7nYHtpM/cOLJAU4+OgDqS+FuetTBZmlT
qqd0i0O+e7zCTVbvlaV5zPOWOLGIBRzNG6qKwe9AALUTQ7E2XWIFjfbbgVe7GSRRRC71Agvkqbnr
cWHQpZMW82/YMiXJ8f2F7wOBCM5FAxPOjQsSBkF1/qzAnTqZysZz9qmH/HA6nVBkgERmDG6+bhZT
gOhZS13l5uxZnwhKrdibVbcXyljuWOBXfa3mQ05VcIS6rkWNYZD+MwZA9iTfgNgMXeW3AdqRzyAm
LnxGtG/DhrH54s9Aqlq6AzfLvCm7FEMt0JYmNQn9PtrrAvUmPQS7SFJUqGMwP++x+Gh09Iu0Dy0L
6k5LXhG1BMdLpb54kxeFj04cXph0bOLEKKfDeks7ZTStT3j+HSyxDil1Hljq05WL1YwnqZoLQrWC
YTPPgTBIZcx1flwWWVDUoxesy7jvEYitlqFOq9oUTORS7y0cBVgWQ8VvDnwnt93SuFQzCNe8ywDj
2a9pFDIf5wGKKMo28+rUWSKE4ffoK5Z5YHajfLHlUDNfXsxNc+ja+np3HHE2yL5cqHg9o3i6/AuJ
CTZllNpJEM/HthQInPKXzbLOnWsrWeR+KAwpT4US8nbXwMlmsCZZg25g4TIZJW3oNsYLzn5LuAUQ
pM6rDaL8q9FmIW1oWF7h6P2bO9NMS5klGWBXAL7n3exQ1xek0x7JMmhQhx7S8ZUPL2BTmykeAqzt
V1JocWSsXjoMoCHcFxkG1RcrrsBgROt+xjkZhln11jLSc3JfPg9Q4ltc3xhpHZ3vk1QFrBTQ05uV
QbQ18vDzjeP0zMDNwYWNZJz/g2mpe1FytqRcJRJMse//BDNM0+4t2osfwLxVtWy0yz4jg8LP90z8
X43YpkMVHHdrkUKBN7p+4g4OVCit+Id6jcGd7kWp3n04ookMgfHaT+3qAlcxHCptd/c3PUvLjngp
8g/WMR5GSf9UYH5M7lly4KvLkYhRA/PbuPVwVw5qIPLTmkJSrISnqWiotRYzW2rtxDMZ6n+Km6dW
kF+5lJDj1M/ycvO1XGXNarj4poWsfMCbVJ0sLV6zGmwB2V1UrY1TPMdyIY+KyJr82zknXbsu/GRH
KmONKfa6jZ983Of+Goq6N14SRfBhjvaSlef5prdHfS8pjp3LrTxSXEE3QEfW1v9JJWQKwC5EJg2y
K9fMRuYO7U9H7EoDTT8V9yPuCE8ai+8+0XphtNelrT9bbUbMnemqytaixEqrxaxlTx9lE4iV1d0z
SUehgQ7FZ9fIPZjXwg0IuO2i3kBXLxLGYyZBl45Lt7JRuzbzpH1k7ui9augDhVFVAR6Fz95S4x+5
6vtMLQU8YaDmil176RQmycsscemq7Dzt8c/WYQFn1TvkgAUMjXHxELAHSLpPBCOSDwNHs0hi526W
15DqpM0mLGSid04CqwV2dLfNvwTpAmKd6jJj/ihcHVXBZOtFK4ULVXw5iqlhVCLfKm2IaK4Ga5cs
Bl1weN3rUCCBuFmm461rZ8l+XlmWP7zHbLJpw1rVFDnG3Uf/v5GIxGwAtO91daQTqWjVKVj/fDzb
6MicbsDmoW/fGBq5lhEABI12MSawI31Yp4gP/ehPNxZ+BdG4kIsOP+TYa/hCzXSpHGboTvP5qRes
PMACRAqywvUeDtweap+or9eIkT2wrrxgp5XPROvLBbRowB68auoTiMhDmkMVEPWDqiuSiWwRdde/
Ae3KDPZmAJoS943zMyuxT2cppg5EKSgc+NeX1BqlBgSoIVcn8icqarhYnuO6nvSI6lYBY+0kvLcF
squWso/uz6Hm3xz4nwr6ASmEzWYpk41lB/Apxa7DR+tUm+25Hj5odw7RCIDqc2k8VbyHF4R4iB9V
JcaoTwHY11YihazcpyXh/a9rI7eSSQNdAdjB7tsC2KoouT8MyWUXRb4LFN/rjNwO5dsGtmNpjNbI
jd63la8ULywNEA92DaHaMQ2ORaSUY884V/anMzqy2Pr95pXT+J8v5fo2m+S9JfTdsHzWNOtcFYJu
Zgp4gVdnNcSVyRswnzY9etY1a1RNl8TEJW9CWO/T67CAuY5Bmm5g7RaQmh9yUcCXlZGCHhb0IAhf
eh1EnBf8AC0JtiUZoxnNQTkIZPz3vgheOZSIJ8R0MgCUOS1D7NtPCXl+ZMhshzqmkuXjTAWWuPlQ
Ha5tp/YHG2SqB3yBN1W1sdllMlG7Fem5JVK9msTZUjNe8J++3427Atj51999I1B/Vq/uVWOY2C32
mGtxr00h0pfaIIetXxAfnfgTf64xaT7eRUc5CZyrCZmf+fkWrakwIKhWFbqbEbXRJyiYmbM7BF8E
KixCaQhudPohWEe0xYjqx3OryExcZ3P1qXtz8zSBbZwwPF64M31rXCJ/HAcxdPveuVMxcetu7oT/
hQ6teajzSKW0vqFUHbus4SANSl1jcKwfT049fdDSfpnhesL9FlY40J09ce4Qs+Ni7LC/uXqNP0c4
j4fEnfeeMTZjzuNT7o71trfCc7ql15URj8vSWbtSDbCiRmyXKlOAPjmtdFBMc6JzNkjxFlQg9Coq
i5NJ2Cija8Xzxpi1biOLPv7DnV5wY6Tx5LP1PbEEkDwpdq1m/39YJvQLT+gFRuQaxNsGda3AQMPm
0QFpCGvrIVF3dZs0Jat1+4aQFNaFfbdzhsXDgVe74KOqPejydo/dpSvGp8C3A5mwbtbIH/XC3OAs
wyE3eXvfs+O/t36ucLO0/P3y1K1d5J+Dtr8ZUV/Tz9j74+Pcis7csGVsASb+jrmhtPXzbkQQ/WMt
TR85oaV87qJYiJmI6k85OBYXVezVzUpHJ55LajG8TiYeN/oFW/oEkfzNqA6fyrZ6LlO3O1zlSeZV
PMsJu+2ZtMltpspialZCuSMm3GP1wj7Ln7hzUMrB73Ky58Mo2MkbYMTzXgykZuH/DpkEkvVpTEY+
r0cxRncGgk8fz1TiHyY3fs3wMv9ToX+ZuDFriiOmPAPQvMu0RkHuaUFbabVUaJsOJsOwSB6ljUnI
/PA0f+4KHGQt9j7KMYTx9nfnEWxooysVp0C1CZfMaBPEsmxrIsdCIxbyioBVlVlS0/OdLuFuKP1R
wl+L6xb5jVOM85y8JiF4LWzTJuyQCvxvGg0aQ/2zduFXAiuBovLj8qm+5wCOSdURxeHIFUGZjqZN
sqg78QObAiA9rKJ/PgDQZneof6XuNvN0bM1MGxMhF/p+fsGbhxJqFobhN2+HGMRdinh5A2rh1Uow
60WnoXzsLvtqDvXt7SVrSfr71Dg8ltulVzqvMPs9kDOj+CPq4Grc/78rp4Rk/8Pnzdlf9A43ZAem
O4a/8V9M1osJqrwyd/uB5L40L9HDt91t8Ydw8aSmCY8gNPZyBWEZYCv58RRAoht/5hARIEqsl1PY
e2n1H5vW4l1YUvXRQEOCKU+PyVySs1DG4JSievTq7fcpLi7PX6CIV8tdKI0hvn8a7QrIPsphV7Se
Rp4kW8GZnc8liwEUvyF/Asi3G4bktDC4nIgk+cDfbuf8UZ1Fbbb7Ynp8vhuv6MLMwMwzLM+kF14m
QZErkUZVQfqjDKMbsCw/0pPrWJpOYqlWSrNQ3Fi0uQNvFxQag1xO/JN+SdI2JXlP0c0+GCcigZUV
orBnZt427k/vd7BuVieFeMbRR1DQC8rcP3mdnvnjhc10/TDWG9aTW+eJr5iVVMnrQqLfXj24wxs/
Qx5UAKtKngytJ7T2A6zUyQXOIgLwg4c/pvckT0UPnyFpEwq0vGNZi3tSyHGKypiU1DK4hZl/+8Zi
0B11Wd1P/CWjhL90PaxJ6xTa0o0vZCyikJRtLtO8BsI1ZCYysEHZYdMMYoUd4lCiI3t7e1g/Ou4T
brCYtw3TBXGjNWEj7EU+LkmJGnz/NA6bBsCjugNzIpIH++tYYG0z0L/J8DLa9o9PmIbMho2rpl8Y
u4dYT7PF7ccbh06kfGLRYdL4HYqvjm4DafEaB1jOmqcZBxXLUD09cLNcYdFh9qwRzExkhhiCmkCI
7qKrZ975eyNOPeAgDkkx+p0fEp2EaIWCyR9PxIjAguOPx0pfE6+Y9OgivNiHkOnuFxIuS5Hzpa+c
VWyicDjuvFDzmblQTv+UIOSxetQKKISq8vGm1seJh8nLnacguXrcThPDCGzhvkGs7/DT85z9Gw6P
D+ZMt/GU/LI/Mi3n4lUwJkrnduEqVw4CnAfF+fOj9EmVZiuqugU7tAtDAsh21GiDnY/6dyjD/gn6
Sv2eKZRo5JHQKkS7gsx4IEIU6346qBYS7Dr2bnDzWLn5gcJYgUyPo33oe48XeXZHd1TZT6wD3AMM
Ko9rMjiNe00iYiGODH61DWpi8JpqusQEIEE7H+RCVRs3TJMctb64fp2Rs0bPP/9RlgqZ9CpGHZfU
ntHJdCfosW5p7XM44YVztBkybOqLVAG9tpXOiiF5sYEhcRu5nfcb4rWOqbdQihk1lgy8bCfKuaDv
Bu3pWg//bqLKwK0//4JAs/7p9FqPYHnPecfDPW7G0zLsyqP9ZL4DwtjoTyvjxqiexAfuZRo/jlfH
udJfRvO2FtafeU6m3OexotBiei4YVg2wU8DOxaSQeCekjb7A+SnWkFJuR5ZSzblaum0OrX4n8d9z
PU8uMmA6w6Ij4sZZxHimlYiOyM9A3Z7iNkVKJ73hbOIWFgd994sGBX66xLD/URX9hP5UmWtdcJn4
a1zSXK77HySzb10NXkEQM0m/WgrfciIAAVafDWPEygmXRZcfYg/QYO4DeE61xS+qI/W6gsmheltO
xdcVFMz6GXNfu3mSStAvxT99ZGJAxCyHUHVjbRV3ZB+TnvKh0w1fjIetbDq9zsVFJQl6cdN4f1lg
jybdHr63XTjt2ErX/zZpNNfn0iD7dQ0FriHME4kARAh1GEfGcGFrJQXiJ/DoxguGhdudMYAcxegW
S1ZTYG7Eq7/vcL/4fwB7RWGA5vuq5bD9hI6lJ10JiLfm4DUTvfxVTIdIDnBWIp7fVf6WAcekSl8J
rPVi8J/9YzAo57Dmb4S2lFtsjHip5ydGjydExNRI6wXITbic2W/qUCSHcJtnMt4rVyHWj/Q17V5I
g/zDR4VlN9NQ/RXMqZhEexo9ou2WJQYYYuLkrpk+hnza6gdl4BHpim23gNFtlH31U2EYbUwtbdnH
6rjKcDfGkn6uH8CveKF/i22hCPgS4mZc/wiZtHiAA4cY4LQ+nzuhMntnZs9uDkGC7v1mj93CF0yJ
/NmTWwqnLoUoSOktHeNFLpqAmaFSdSXG9t5Goi5Kvu5+ocB0yFyuupyaRvoM9fvJliX0YN85JhyE
DxppJzSpjA3IqIVMZcBuq4pQayJb2l+LY2mUomRxoYgT8CeE1hV1Rsd4PTsi1LJ2n3WvR4cl4Y5G
UrAHoz5cjXT8i+ckCKE=
`pragma protect end_protected
